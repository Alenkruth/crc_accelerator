
* cell freepdk45_sram_4kbytes_1rw_32x1024_8
* pin addr0[0]
* pin addr0[1]
* pin addr0[2]
* pin wmask0[0]
* pin wmask0[1]
* pin wmask0[2]
* pin wmask0[3]
* pin din0[0]
* pin din0[1]
* pin din0[2]
* pin dout0[0]
* pin din0[3]
* pin din0[4]
* pin dout0[1]
* pin din0[5]
* pin dout0[2]
* pin din0[6]
* pin din0[7]
* pin dout0[3]
* pin din0[8]
* pin din0[9]
* pin din0[10]
* pin dout0[4]
* pin din0[11]
* pin din0[12]
* pin dout0[5]
* pin din0[13]
* pin dout0[6]
* pin din0[14]
* pin din0[15]
* pin din0[16]
* pin dout0[7]
* pin din0[17]
* pin dout0[8]
* pin din0[18]
* pin din0[19]
* pin dout0[9]
* pin din0[20]
* pin din0[21]
* pin dout0[10]
* pin din0[22]
* pin din0[23]
* pin dout0[11]
* pin din0[24]
* pin din0[25]
* pin dout0[12]
* pin din0[26]
* pin din0[27]
* pin dout0[13]
* pin din0[28]
* pin din0[29]
* pin dout0[14]
* pin din0[30]
* pin din0[31]
* pin dout0[15]
* pin din0[32]
* pin spare_wen0
* pin dout0[16]
* pin dout0[17]
* pin dout0[18]
* pin dout0[19]
* pin dout0[20]
* pin dout0[21]
* pin dout0[22]
* pin dout0[23]
* pin dout0[24]
* pin dout0[25]
* pin dout0[26]
* pin dout0[27]
* pin dout0[28]
* pin csb0
* pin web0
* pin clk0
* pin dout0[29]
* pin dout0[31]
* pin dout0[32]
* pin dout0[30]
* pin addr0[3]
* pin addr0[4]
* pin addr0[5]
* pin addr0[7]
* pin addr0[6]
* pin addr0[8]
* pin addr0[9]
* pin addr0[10]
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 72 73 74 75 76 77 82 84 86 87 88 89 93 94 95 100 101
* net 1 addr0[0]
* net 2 addr0[1]
* net 3 addr0[2]
* net 4 wmask0[0]
* net 5 wmask0[1]
* net 6 wmask0[2]
* net 7 wmask0[3]
* net 8 din0[0]
* net 9 din0[1]
* net 10 din0[2]
* net 11 dout0[0]
* net 12 din0[3]
* net 13 din0[4]
* net 14 dout0[1]
* net 15 din0[5]
* net 16 dout0[2]
* net 17 din0[6]
* net 18 din0[7]
* net 19 dout0[3]
* net 20 din0[8]
* net 21 din0[9]
* net 22 din0[10]
* net 23 dout0[4]
* net 24 din0[11]
* net 25 din0[12]
* net 26 dout0[5]
* net 27 din0[13]
* net 28 dout0[6]
* net 29 din0[14]
* net 30 din0[15]
* net 31 din0[16]
* net 32 dout0[7]
* net 33 din0[17]
* net 34 dout0[8]
* net 35 din0[18]
* net 36 din0[19]
* net 37 dout0[9]
* net 38 din0[20]
* net 39 din0[21]
* net 40 dout0[10]
* net 41 din0[22]
* net 42 din0[23]
* net 43 dout0[11]
* net 44 din0[24]
* net 45 din0[25]
* net 46 dout0[12]
* net 47 din0[26]
* net 48 din0[27]
* net 49 dout0[13]
* net 50 din0[28]
* net 51 din0[29]
* net 52 dout0[14]
* net 53 din0[30]
* net 54 din0[31]
* net 55 dout0[15]
* net 56 din0[32]
* net 57 spare_wen0
* net 58 dout0[16]
* net 59 dout0[17]
* net 60 dout0[18]
* net 61 dout0[19]
* net 62 dout0[20]
* net 63 dout0[21]
* net 64 dout0[22]
* net 65 dout0[23]
* net 66 dout0[24]
* net 67 dout0[25]
* net 68 dout0[26]
* net 69 dout0[27]
* net 70 dout0[28]
* net 72 csb0
* net 73 web0
* net 74 clk0
* net 75 dout0[29]
* net 76 dout0[31]
* net 77 dout0[32]
* net 82 dout0[30]
* net 84 addr0[3]
* net 86 addr0[4]
* net 87 addr0[5]
* net 88 addr0[7]
* net 89 addr0[6]
* net 93 addr0[8]
* net 94 addr0[9]
* net 95 addr0[10]
* net 100 vdd
* net 101 gnd
* cell instance $3 r0 *1 27.29,3.2
X$3 1 142 2 141 3 140 71 100 101
+ freepdk45_sram_4kbytes_1rw_32x1024_8_col_addr_dff
* cell instance $9 r0 *1 35.87,3.2
X$9 4 139 5 137 6 138 7 136 71 100 101
+ freepdk45_sram_4kbytes_1rw_32x1024_8_wmask_dff
* cell instance $18 r0 *1 47.31,3.2
X$18 71 8 135 9 134 10 133 12 132 13 131 15 130 17 129 18 128 20 127 21 126 22
+ 125 24 124 25 123 27 122 29 121 30 120 31 119 33 118 35 117 36 116 38 115 39
+ 114 41 113 42 112 44 111 45 110 47 109 48 108 50 107 51 106 53 105 54 104 56
+ 103 100 101 freepdk45_sram_4kbytes_1rw_32x1024_8_data_dff
* cell instance $26 r0 *1 24.71,11.55
X$26 142 141 140 139 137 138 136 81 135 134 133 132 131 130 129 128 127 126 125
+ 124 123 122 121 120 119 118 117 116 115 114 113 112 111 110 109 108 107 106
+ 105 104 103 102 80 78 11 14 16 19 23 26 28 32 34 37 40 43 46 49 52 55 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 75 82 76 77 79 85 92 91 90 98 97 96 99 83
+ 100 101 freepdk45_sram_4kbytes_1rw_32x1024_8_bank
* cell instance $118 r0 *1 141.69,3.2
X$118 57 102 71 100 101 freepdk45_sram_4kbytes_1rw_32x1024_8_spare_wen_dff
* cell instance $146 r0 *1 3.2525,14.635
X$146 72 71 74 73 78 79 81 83 80 100 101
+ freepdk45_sram_4kbytes_1rw_32x1024_8_control_logic_rw
* cell instance $147 r0 *1 21.57,70.275
X$147 84 85 86 92 87 91 89 90 88 98 93 97 94 96 95 99 71 100 101
+ freepdk45_sram_4kbytes_1rw_32x1024_8_row_addr_dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_spare_wen_dff
* pin din_0
* pin dout_0
* pin clk
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_spare_wen_dff 1 2 3 4 5
* net 1 din_0
* net 2 dout_0
* net 3 clk
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 5 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_spare_wen_dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_wmask_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin clk
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_wmask_dff 1 2 3 4 5 6 7 8 9 10 11
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 din_2
* net 6 dout_2
* net 7 din_3
* net 8 dout_3
* net 9 clk
* net 10 vdd
* net 11 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 9 10 11 dff
* cell instance $2 r0 *1 2.86,0
X$2 4 3 9 10 11 dff
* cell instance $3 r0 *1 5.72,0
X$3 6 5 9 10 11 dff
* cell instance $4 r0 *1 8.58,0
X$4 8 7 9 10 11 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_wmask_dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_control_logic_rw
* pin csb
* pin clk_buf
* pin clk
* pin web
* pin s_en
* pin rbl_bl
* pin w_en
* pin wl_en
* pin p_en_bar
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_control_logic_rw 1 2 4 8 13 14 16
+ 17 18 19 20
* net 1 csb
* net 2 clk_buf
* net 4 clk
* net 8 web
* net 13 s_en
* net 14 rbl_bl
* net 16 w_en
* net 17 wl_en
* net 18 p_en_bar
* net 19 vdd
* net 20 gnd
* cell instance $1 r0 *1 0,0
X$1 1 3 8 10 6 2 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_array
* cell instance $3 r0 *1 6.385,4.94
X$3 9 2 3 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2_0
* cell instance $5 m0 *1 6.385,4.94
X$5 2 7 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
* cell instance $9 r0 *1 6.385,0
X$9 2 4 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_2
* cell instance $17 m0 *1 7.0725,4.94
X$17 5 7 3 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2_0
* cell instance $20 m0 *1 6.385,9.88
X$20 13 12 5 10 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_1
* cell instance $21 m0 *1 6.385,19.76
X$21 17 5 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_3
* cell instance $22 r0 *1 6.385,9.88
X$22 16 6 11 5 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_0
* cell instance $32 m0 *1 6.385,14.82
X$32 9 12 15 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_2
* cell instance $43 r0 *1 6.385,14.82
X$43 12 11 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
* cell instance $45 m0 *1 0,32.11
X$45 12 14 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_delay_chain
* cell instance $52 m0 *1 7.2875,14.82
X$52 18 15 19 20 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_6
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_control_logic_rw

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_col_addr_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin clk
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_col_addr_dff 1 2 3 4 5 6 7 8 9
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 din_2
* net 6 dout_2
* net 7 clk
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 7 8 9 dff
* cell instance $2 r0 *1 2.86,0
X$2 4 3 7 8 9 dff
* cell instance $3 r0 *1 5.72,0
X$3 6 5 7 8 9 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_col_addr_dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_row_addr_dff
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin din_4
* pin dout_4
* pin din_5
* pin dout_5
* pin din_6
* pin dout_6
* pin din_7
* pin dout_7
* pin clk
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_row_addr_dff 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
* net 1 din_0
* net 2 dout_0
* net 3 din_1
* net 4 dout_1
* net 5 din_2
* net 6 dout_2
* net 7 din_3
* net 8 dout_3
* net 9 din_4
* net 10 dout_4
* net 11 din_5
* net 12 dout_5
* net 13 din_6
* net 14 dout_6
* net 15 din_7
* net 16 dout_7
* net 17 clk
* net 18 vdd
* net 19 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 17 18 19 dff
* cell instance $2 m0 *1 0,4.94
X$2 4 3 17 18 19 dff
* cell instance $3 r0 *1 0,4.94
X$3 6 5 17 18 19 dff
* cell instance $4 m0 *1 0,9.88
X$4 8 7 17 18 19 dff
* cell instance $5 r0 *1 0,9.88
X$5 10 9 17 18 19 dff
* cell instance $6 m0 *1 0,14.82
X$6 12 11 17 18 19 dff
* cell instance $7 r0 *1 0,14.82
X$7 14 13 17 18 19 dff
* cell instance $8 m0 *1 0,19.76
X$8 16 15 17 18 19 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_row_addr_dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_data_dff
* pin clk
* pin din_0
* pin dout_0
* pin din_1
* pin dout_1
* pin din_2
* pin dout_2
* pin din_3
* pin dout_3
* pin din_4
* pin dout_4
* pin din_5
* pin dout_5
* pin din_6
* pin dout_6
* pin din_7
* pin dout_7
* pin din_8
* pin dout_8
* pin din_9
* pin dout_9
* pin din_10
* pin dout_10
* pin din_11
* pin dout_11
* pin din_12
* pin dout_12
* pin din_13
* pin dout_13
* pin din_14
* pin dout_14
* pin din_15
* pin dout_15
* pin din_16
* pin dout_16
* pin din_17
* pin dout_17
* pin din_18
* pin dout_18
* pin din_19
* pin dout_19
* pin din_20
* pin dout_20
* pin din_21
* pin dout_21
* pin din_22
* pin dout_22
* pin din_23
* pin dout_23
* pin din_24
* pin dout_24
* pin din_25
* pin dout_25
* pin din_26
* pin dout_26
* pin din_27
* pin dout_27
* pin din_28
* pin dout_28
* pin din_29
* pin dout_29
* pin din_30
* pin dout_30
* pin din_31
* pin dout_31
* pin din_32
* pin dout_32
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_data_dff 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69
* net 1 clk
* net 2 din_0
* net 3 dout_0
* net 4 din_1
* net 5 dout_1
* net 6 din_2
* net 7 dout_2
* net 8 din_3
* net 9 dout_3
* net 10 din_4
* net 11 dout_4
* net 12 din_5
* net 13 dout_5
* net 14 din_6
* net 15 dout_6
* net 16 din_7
* net 17 dout_7
* net 18 din_8
* net 19 dout_8
* net 20 din_9
* net 21 dout_9
* net 22 din_10
* net 23 dout_10
* net 24 din_11
* net 25 dout_11
* net 26 din_12
* net 27 dout_12
* net 28 din_13
* net 29 dout_13
* net 30 din_14
* net 31 dout_14
* net 32 din_15
* net 33 dout_15
* net 34 din_16
* net 35 dout_16
* net 36 din_17
* net 37 dout_17
* net 38 din_18
* net 39 dout_18
* net 40 din_19
* net 41 dout_19
* net 42 din_20
* net 43 dout_20
* net 44 din_21
* net 45 dout_21
* net 46 din_22
* net 47 dout_22
* net 48 din_23
* net 49 dout_23
* net 50 din_24
* net 51 dout_24
* net 52 din_25
* net 53 dout_25
* net 54 din_26
* net 55 dout_26
* net 56 din_27
* net 57 dout_27
* net 58 din_28
* net 59 dout_28
* net 60 din_29
* net 61 dout_29
* net 62 din_30
* net 63 dout_30
* net 64 din_31
* net 65 dout_31
* net 66 din_32
* net 67 dout_32
* net 68 vdd
* net 69 gnd
* cell instance $1 r0 *1 71.5,0
X$1 53 52 1 68 69 dff
* cell instance $2 r0 *1 22.88,0
X$2 19 18 1 68 69 dff
* cell instance $3 r0 *1 20.02,0
X$3 17 16 1 68 69 dff
* cell instance $4 r0 *1 17.16,0
X$4 15 14 1 68 69 dff
* cell instance $5 r0 *1 14.3,0
X$5 13 12 1 68 69 dff
* cell instance $6 r0 *1 11.44,0
X$6 11 10 1 68 69 dff
* cell instance $7 r0 *1 8.58,0
X$7 9 8 1 68 69 dff
* cell instance $8 r0 *1 68.64,0
X$8 51 50 1 68 69 dff
* cell instance $9 r0 *1 2.86,0
X$9 5 4 1 68 69 dff
* cell instance $10 r0 *1 74.36,0
X$10 55 54 1 68 69 dff
* cell instance $11 r0 *1 77.22,0
X$11 57 56 1 68 69 dff
* cell instance $12 r0 *1 80.08,0
X$12 59 58 1 68 69 dff
* cell instance $13 r0 *1 82.94,0
X$13 61 60 1 68 69 dff
* cell instance $14 r0 *1 85.8,0
X$14 63 62 1 68 69 dff
* cell instance $15 r0 *1 88.66,0
X$15 65 64 1 68 69 dff
* cell instance $16 r0 *1 91.52,0
X$16 67 66 1 68 69 dff
* cell instance $17 r0 *1 5.72,0
X$17 7 6 1 68 69 dff
* cell instance $18 r0 *1 45.76,0
X$18 35 34 1 68 69 dff
* cell instance $19 r0 *1 48.62,0
X$19 37 36 1 68 69 dff
* cell instance $20 r0 *1 0,0
X$20 3 2 1 68 69 dff
* cell instance $21 r0 *1 42.9,0
X$21 33 32 1 68 69 dff
* cell instance $22 r0 *1 40.04,0
X$22 31 30 1 68 69 dff
* cell instance $23 r0 *1 37.18,0
X$23 29 28 1 68 69 dff
* cell instance $24 r0 *1 34.32,0
X$24 27 26 1 68 69 dff
* cell instance $25 r0 *1 31.46,0
X$25 25 24 1 68 69 dff
* cell instance $26 r0 *1 28.6,0
X$26 23 22 1 68 69 dff
* cell instance $27 r0 *1 25.74,0
X$27 21 20 1 68 69 dff
* cell instance $28 r0 *1 51.48,0
X$28 39 38 1 68 69 dff
* cell instance $29 r0 *1 54.34,0
X$29 41 40 1 68 69 dff
* cell instance $30 r0 *1 57.2,0
X$30 43 42 1 68 69 dff
* cell instance $31 r0 *1 60.06,0
X$31 45 44 1 68 69 dff
* cell instance $32 r0 *1 62.92,0
X$32 47 46 1 68 69 dff
* cell instance $33 r0 *1 65.78,0
X$33 49 48 1 68 69 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_data_dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_bank
* pin addr0_0
* pin addr0_1
* pin addr0_2
* pin bank_wmask0_0
* pin bank_wmask0_1
* pin bank_wmask0_2
* pin bank_wmask0_3
* pin w_en0
* pin din0_0
* pin din0_1
* pin din0_2
* pin din0_3
* pin din0_4
* pin din0_5
* pin din0_6
* pin din0_7
* pin din0_8
* pin din0_9
* pin din0_10
* pin din0_11
* pin din0_12
* pin din0_13
* pin din0_14
* pin din0_15
* pin din0_16
* pin din0_17
* pin din0_18
* pin din0_19
* pin din0_20
* pin din0_21
* pin din0_22
* pin din0_23
* pin din0_24
* pin din0_25
* pin din0_26
* pin din0_27
* pin din0_28
* pin din0_29
* pin din0_30
* pin din0_31
* pin din0_32
* pin bank_spare_wen0_0
* pin p_en_bar0
* pin s_en0
* pin dout0_0
* pin dout0_1
* pin dout0_2
* pin dout0_3
* pin dout0_4
* pin dout0_5
* pin dout0_6
* pin dout0_7
* pin dout0_8
* pin dout0_9
* pin dout0_10
* pin dout0_11
* pin dout0_12
* pin dout0_13
* pin dout0_14
* pin dout0_15
* pin dout0_16
* pin dout0_17
* pin dout0_18
* pin dout0_19
* pin dout0_20
* pin dout0_21
* pin dout0_22
* pin dout0_23
* pin dout0_24
* pin dout0_25
* pin dout0_26
* pin dout0_27
* pin dout0_28
* pin dout0_29
* pin dout0_30
* pin dout0_31
* pin dout0_32
* pin rbl_bl_0_0
* pin addr0_3
* pin addr0_4
* pin addr0_5
* pin addr0_6
* pin addr0_7
* pin addr0_8
* pin addr0_9
* pin addr0_10
* pin wl_en0
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_bank 1 3 5 7 8 9 10 11 13 14 15 16
+ 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 48 49 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71
+ 72 73 74 75 76 77 78 79 80 81 82 83 84 86 602 603 604 605 606 607 608 609 610
+ 741 742
* net 1 addr0_0
* net 3 addr0_1
* net 5 addr0_2
* net 7 bank_wmask0_0
* net 8 bank_wmask0_1
* net 9 bank_wmask0_2
* net 10 bank_wmask0_3
* net 11 w_en0
* net 13 din0_0
* net 14 din0_1
* net 15 din0_2
* net 16 din0_3
* net 17 din0_4
* net 18 din0_5
* net 19 din0_6
* net 20 din0_7
* net 21 din0_8
* net 22 din0_9
* net 23 din0_10
* net 24 din0_11
* net 25 din0_12
* net 26 din0_13
* net 27 din0_14
* net 28 din0_15
* net 29 din0_16
* net 30 din0_17
* net 31 din0_18
* net 32 din0_19
* net 33 din0_20
* net 34 din0_21
* net 35 din0_22
* net 36 din0_23
* net 37 din0_24
* net 38 din0_25
* net 39 din0_26
* net 40 din0_27
* net 41 din0_28
* net 42 din0_29
* net 43 din0_30
* net 44 din0_31
* net 45 din0_32
* net 46 bank_spare_wen0_0
* net 48 p_en_bar0
* net 49 s_en0
* net 52 dout0_0
* net 53 dout0_1
* net 54 dout0_2
* net 55 dout0_3
* net 56 dout0_4
* net 57 dout0_5
* net 58 dout0_6
* net 59 dout0_7
* net 60 dout0_8
* net 61 dout0_9
* net 62 dout0_10
* net 63 dout0_11
* net 64 dout0_12
* net 65 dout0_13
* net 66 dout0_14
* net 67 dout0_15
* net 68 dout0_16
* net 69 dout0_17
* net 70 dout0_18
* net 71 dout0_19
* net 72 dout0_20
* net 73 dout0_21
* net 74 dout0_22
* net 75 dout0_23
* net 76 dout0_24
* net 77 dout0_25
* net 78 dout0_26
* net 79 dout0_27
* net 80 dout0_28
* net 81 dout0_29
* net 82 dout0_30
* net 83 dout0_31
* net 84 dout0_32
* net 86 rbl_bl_0_0
* net 602 addr0_3
* net 603 addr0_4
* net 604 addr0_5
* net 605 addr0_6
* net 606 addr0_7
* net 607 addr0_8
* net 608 addr0_9
* net 609 addr0_10
* net 610 wl_en0
* net 741 vdd
* net 742 gnd
* cell instance $1 r0 *1 5.415,0.1375
X$1 2 4 6 12 47 51 50 85 1 3 5 741 742
+ freepdk45_sram_4kbytes_1rw_32x1024_8_column_decoder
* cell instance $2 m0 *1 26.49,22.985
X$2 86 87 88 89 90 92 93 94 96 98 99 100 102 103 104 106 108 109 110 111 112
+ 113 114 115 116 117 118 119 120 122 124 125 126 127 128 129 130 131 132 134
+ 135 136 138 139 140 142 143 144 145 146 147 148 149 150 151 152 153 154 155
+ 156 157 158 159 160 161 162 164 165 166 167 168 169 170 171 172 173 174 175
+ 176 177 178 179 180 181 182 183 184 185 186 187 188 190 191 192 194 196 198
+ 200 201 202 203 204 205 206 208 209 210 211 212 213 214 215 216 217 218 219
+ 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
+ 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 276 277 278
+ 279 280 281 282 283 284 286 287 288 289 290 291 292 294 296 297 298 299 300
+ 302 303 304 306 307 308 309 310 312 313 314 315 316 317 318 320 321 322 323
+ 324 325 326 328 329 330 331 332 334 335 336 337 338 339 340 341 342 344 345
+ 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364
+ 365 366 367 368 369 370 371 372 373 374 375 376 378 379 380 381 382 383 384
+ 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403
+ 404 405 406 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 436 437 438 440 441 442 443 444
+ 446 447 448 449 450 451 452 453 454 456 457 458 459 460 461 462 464 465 466
+ 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485
+ 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504
+ 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 524
+ 525 526 527 528 529 530 531 532 534 535 536 537 538 539 540 542 543 544 545
+ 546 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565
+ 566 568 570 571 572 573 574 576 577 578 580 582 584 586 587 588 589 590 592
+ 593 594 595 596 597 598 599 600 601 91 95 97 101 105 107 121 123 133 137 141
+ 163 189 193 195 197 199 207 237 275 285 293 295 301 305 311 319 327 333 48
+ 343 377 407 435 439 445 455 463 523 533 541 547 567 569 575 579 581 583 585
+ 591 85 50 51 47 12 6 4 2 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 49
+ 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 11 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46
+ 7 8 9 10 741 742 freepdk45_sram_4kbytes_1rw_32x1024_8_port_data
* cell instance $20 r0 *1 26.49,22.985
X$20 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107
+ 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126
+ 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145
+ 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259
+ 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278
+ 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297
+ 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316
+ 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335
+ 336 337 338 339 340 341 342 343 674 662 714 611 675 658 657 647 653 642 650
+ 685 649 640 664 630 693 661 663 716 639 698 656 654 619 633 648 687 689 651
+ 676 677 678 699 670 671 665 627 694 669 679 636 710 659 696 680 734 660 708
+ 652 738 666 655 667 718 703 622 727 620 629 616 625 690 736 732 344 345 346
+ 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364 365
+ 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384
+ 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403
+ 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479
+ 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498
+ 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517
+ 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536
+ 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554 555
+ 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573 574
+ 575 576 577 578 579 580 581 582 583 584 585 586 587 588 589 590 591 592 593
+ 594 595 596 597 598 599 600 601 709 707 717 641 706 646 672 711 715 621 618
+ 712 726 729 713 634 691 728 617 673 737 643 735 733 697 692 730 644 623 684
+ 740 739 695 681 722 721 645 731 682 683 686 720 688 719 614 631 612 724 628
+ 723 705 704 613 668 632 638 702 624 725 635 701 700 637 626 615 741 742
+ freepdk45_sram_4kbytes_1rw_32x1024_8_capped_replica_bitcell_array
* cell instance $22 r0 *1 0,25.965
X$22 610 703 710 680 708 696 732 736 714 716 639 636 640 602 603 604 605 606
+ 607 608 609 642 611 627 671 670 678 676 651 648 654 656 619 633 687 689 698
+ 699 694 685 693 690 734 738 718 727 629 630 625 616 620 622 667 666 655 652
+ 660 659 661 662 663 664 649 650 653 647 657 658 675 677 674 679 669 665 668
+ 672 621 673 623 624 628 626 612 613 615 614 617 618 641 643 644 645 634 646
+ 631 632 637 635 638 723 724 725 728 729 717 715 719 720 721 722 740 739 730
+ 733 737 735 731 726 691 692 695 697 681 684 682 683 688 686 707 709 711 706
+ 713 712 701 700 704 702 705 741 742
+ freepdk45_sram_4kbytes_1rw_32x1024_8_port_address
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_bank

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_2
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_2 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_2

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_array
* pin din_0
* pin dout_bar_0
* pin din_1
* pin dout_1
* pin dout_bar_1
* pin clk
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_array 1 3 4 5 6 7 8 9
* net 1 din_0
* net 2 dout_0
* net 3 dout_bar_0
* net 4 din_1
* net 5 dout_1
* net 6 dout_bar_1
* net 7 clk
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 0,0
X$1 3 2 7 1 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_0
* cell instance $2 m0 *1 0,4.94
X$2 6 5 7 4 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pand2_0
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pand2_0 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_1
* cell instance $2 r0 *1 0.75,0
X$2 2 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_1
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pand2_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_6
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_6 5 6 8 9
* net 5 Z
* net 6 A
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 1.375,0
X$1 1 2 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_9
* cell instance $2 r0 *1 0.6875,0
X$2 7 1 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
* cell instance $3 r0 *1 2.0625,0
X$3 2 3 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_17
* cell instance $4 r0 *1 3.3,0
X$4 3 4 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_18
* cell instance $5 r0 *1 6.1875,0
X$5 4 5 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_19
* cell instance $6 r0 *1 0,0
X$6 6 7 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_6

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_delay_chain
* pin out
* pin in
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_delay_chain 1 10 11 12
* net 1 out
* net 10 in
* net 11 vdd
* net 12 gnd
* cell instance $2 r0 *1 0.6875,19.76
X$2 1 37 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $5 r0 *1 1.375,19.76
X$5 1 36 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $8 r0 *1 2.0625,19.76
X$8 1 35 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $11 r0 *1 2.75,19.76
X$11 1 34 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $14 r0 *1 0,19.76
X$14 9 1 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $17 r0 *1 1.375,0
X$17 2 29 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $20 r0 *1 0.6875,0
X$20 2 46 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $23 m0 *1 0,4.94
X$23 2 3 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $25 r0 *1 2.0625,0
X$25 2 45 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $28 r0 *1 2.75,0
X$28 2 47 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $31 r0 *1 0,0
X$31 10 2 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $34 m0 *1 2.0625,4.94
X$34 3 22 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $37 r0 *1 0,4.94
X$37 3 4 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $39 m0 *1 2.75,4.94
X$39 3 23 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $42 m0 *1 0.6875,4.94
X$42 3 16 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $47 m0 *1 1.375,4.94
X$47 3 13 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $50 r0 *1 1.375,4.94
X$50 4 31 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $55 r0 *1 2.75,4.94
X$55 4 33 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $58 r0 *1 2.0625,4.94
X$58 4 32 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $61 m0 *1 0,9.88
X$61 4 5 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $63 r0 *1 0.6875,4.94
X$63 4 30 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $66 m0 *1 2.0625,9.88
X$66 5 15 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $69 r0 *1 0,9.88
X$69 5 6 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $71 m0 *1 0.6875,9.88
X$71 5 27 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $74 m0 *1 2.75,9.88
X$74 5 21 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $79 m0 *1 1.375,9.88
X$79 5 14 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $82 m0 *1 0,14.82
X$82 6 7 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $84 r0 *1 2.0625,9.88
X$84 6 43 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $87 r0 *1 0.6875,9.88
X$87 6 48 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $92 r0 *1 1.375,9.88
X$92 6 44 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $95 r0 *1 2.75,9.88
X$95 6 42 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $100 m0 *1 2.75,14.82
X$100 7 24 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $103 m0 *1 2.0625,14.82
X$103 7 25 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $106 m0 *1 0.6875,14.82
X$106 7 28 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $109 m0 *1 1.375,14.82
X$109 7 26 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $112 r0 *1 0,14.82
X$112 7 8 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $114 r0 *1 1.375,14.82
X$114 8 40 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $117 r0 *1 0.6875,14.82
X$117 8 41 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $120 r0 *1 2.0625,14.82
X$120 8 39 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $123 r0 *1 2.75,14.82
X$123 8 38 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $128 m0 *1 0,19.76
X$128 8 9 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $130 m0 *1 1.375,19.76
X$130 9 19 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $133 m0 *1 0.6875,19.76
X$133 9 20 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $136 m0 *1 2.0625,19.76
X$136 9 18 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* cell instance $139 m0 *1 2.75,19.76
X$139 9 17 11 12 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_delay_chain

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_1
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_1 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0.965,0
X$1 2 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_5
* cell instance $2 r0 *1 0,0
X$2 3 4 5 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_1

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_0
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_0 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0.965,0
X$1 2 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_4
* cell instance $2 r0 *1 0,0
X$2 3 4 5 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pand3_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_3
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_3 2 3 4 5
* net 2 Z
* net 3 A
* net 4 vdd
* net 5 gnd
* cell instance $1 r0 *1 0,0
X$1 3 1 4 5 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_13
* cell instance $2 r0 *1 1.7875,0
X$2 1 2 4 5 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_14
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_3

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_2
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_2 3 4 8 9
* net 3 Z
* net 4 A
* net 8 vdd
* net 9 gnd
* cell instance $1 r0 *1 1.375,0
X$1 1 6 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_9
* cell instance $2 r0 *1 0.6875,0
X$2 5 1 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
* cell instance $3 r0 *1 2.0625,0
X$3 6 2 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_10
* cell instance $4 r0 *1 3.3,0
X$4 2 7 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_11
* cell instance $5 r0 *1 5.9125,0
X$5 7 3 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_12
* cell instance $6 r0 *1 0,0
X$6 4 5 8 9 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_2

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_column_decoder
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin out_4
* pin out_5
* pin out_6
* pin out_7
* pin in_0
* pin in_1
* pin in_2
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_column_decoder 1 2 3 4 5 6 7 8 9
+ 10 11 12 13
* net 1 out_0
* net 2 out_1
* net 3 out_2
* net 4 out_3
* net 5 out_4
* net 6 out_5
* net 7 out_6
* net 8 out_7
* net 9 in_0
* net 10 in_1
* net 11 in_2
* net 12 vdd
* net 13 gnd
* cell instance $1 r0 *1 0,0
X$1 9 10 1 2 11 3 4 6 5 7 8 12 13
+ freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_column_decoder

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_port_address
* pin wl_en
* pin rbl_wl
* pin wl_0
* pin wl_2
* pin wl_1
* pin wl_3
* pin wl_5
* pin wl_4
* pin wl_6
* pin wl_7
* pin wl_8
* pin wl_9
* pin wl_10
* pin addr_0
* pin addr_1
* pin addr_2
* pin addr_3
* pin addr_4
* pin addr_5
* pin addr_6
* pin addr_7
* pin wl_11
* pin wl_12
* pin wl_13
* pin wl_14
* pin wl_15
* pin wl_16
* pin wl_17
* pin wl_18
* pin wl_19
* pin wl_20
* pin wl_21
* pin wl_22
* pin wl_23
* pin wl_24
* pin wl_25
* pin wl_26
* pin wl_27
* pin wl_28
* pin wl_29
* pin wl_30
* pin wl_31
* pin wl_32
* pin wl_33
* pin wl_34
* pin wl_35
* pin wl_36
* pin wl_37
* pin wl_38
* pin wl_39
* pin wl_40
* pin wl_41
* pin wl_42
* pin wl_43
* pin wl_44
* pin wl_45
* pin wl_46
* pin wl_47
* pin wl_48
* pin wl_49
* pin wl_50
* pin wl_51
* pin wl_52
* pin wl_53
* pin wl_54
* pin wl_55
* pin wl_56
* pin wl_57
* pin wl_58
* pin wl_59
* pin wl_60
* pin wl_61
* pin wl_62
* pin wl_63
* pin wl_64
* pin wl_65
* pin wl_67
* pin wl_66
* pin wl_68
* pin wl_69
* pin wl_71
* pin wl_70
* pin wl_72
* pin wl_73
* pin wl_75
* pin wl_74
* pin wl_76
* pin wl_77
* pin wl_78
* pin wl_79
* pin wl_80
* pin wl_81
* pin wl_83
* pin wl_82
* pin wl_84
* pin wl_85
* pin wl_87
* pin wl_86
* pin wl_88
* pin wl_89
* pin wl_90
* pin wl_91
* pin wl_92
* pin wl_93
* pin wl_95
* pin wl_94
* pin wl_96
* pin wl_97
* pin wl_98
* pin wl_99
* pin wl_101
* pin wl_100
* pin wl_102
* pin wl_103
* pin wl_105
* pin wl_104
* pin wl_106
* pin wl_107
* pin wl_108
* pin wl_109
* pin wl_110
* pin wl_111
* pin wl_113
* pin wl_112
* pin wl_114
* pin wl_115
* pin wl_117
* pin wl_116
* pin wl_118
* pin wl_119
* pin wl_121
* pin wl_120
* pin wl_123
* pin wl_122
* pin wl_125
* pin wl_124
* pin wl_127
* pin wl_126
* pin wl_128
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_port_address 1 2 5 8 9 11 14 15 18
+ 19 21 22 25 26 27 28 29 30 31 32 33 34 38 39 41 42 45 47 50 51 53 54 57 59 61
+ 62 64 66 69 70 73 74 77 78 81 82 85 86 89 90 93 94 97 98 101 102 105 106 109
+ 110 113 114 117 118 121 122 125 126 129 130 133 134 137 138 140 142 145 146
+ 149 150 153 154 157 158 161 162 165 166 169 170 173 174 177 178 181 182 185
+ 186 189 190 193 194 197 198 201 202 205 206 209 210 213 214 217 218 221 222
+ 225 226 229 230 233 234 237 238 241 242 245 246 249 250 253 254 257 258 261
+ 262 265 266 268 269 270
* net 1 wl_en
* net 2 rbl_wl
* net 5 wl_0
* net 8 wl_2
* net 9 wl_1
* net 11 wl_3
* net 14 wl_5
* net 15 wl_4
* net 18 wl_6
* net 19 wl_7
* net 21 wl_8
* net 22 wl_9
* net 25 wl_10
* net 26 addr_0
* net 27 addr_1
* net 28 addr_2
* net 29 addr_3
* net 30 addr_4
* net 31 addr_5
* net 32 addr_6
* net 33 addr_7
* net 34 wl_11
* net 38 wl_12
* net 39 wl_13
* net 41 wl_14
* net 42 wl_15
* net 45 wl_16
* net 47 wl_17
* net 50 wl_18
* net 51 wl_19
* net 53 wl_20
* net 54 wl_21
* net 57 wl_22
* net 59 wl_23
* net 61 wl_24
* net 62 wl_25
* net 64 wl_26
* net 66 wl_27
* net 69 wl_28
* net 70 wl_29
* net 73 wl_30
* net 74 wl_31
* net 77 wl_32
* net 78 wl_33
* net 81 wl_34
* net 82 wl_35
* net 85 wl_36
* net 86 wl_37
* net 89 wl_38
* net 90 wl_39
* net 93 wl_40
* net 94 wl_41
* net 97 wl_42
* net 98 wl_43
* net 101 wl_44
* net 102 wl_45
* net 105 wl_46
* net 106 wl_47
* net 109 wl_48
* net 110 wl_49
* net 113 wl_50
* net 114 wl_51
* net 117 wl_52
* net 118 wl_53
* net 121 wl_54
* net 122 wl_55
* net 125 wl_56
* net 126 wl_57
* net 129 wl_58
* net 130 wl_59
* net 133 wl_60
* net 134 wl_61
* net 137 wl_62
* net 138 wl_63
* net 140 wl_64
* net 142 wl_65
* net 145 wl_67
* net 146 wl_66
* net 149 wl_68
* net 150 wl_69
* net 153 wl_71
* net 154 wl_70
* net 157 wl_72
* net 158 wl_73
* net 161 wl_75
* net 162 wl_74
* net 165 wl_76
* net 166 wl_77
* net 169 wl_78
* net 170 wl_79
* net 173 wl_80
* net 174 wl_81
* net 177 wl_83
* net 178 wl_82
* net 181 wl_84
* net 182 wl_85
* net 185 wl_87
* net 186 wl_86
* net 189 wl_88
* net 190 wl_89
* net 193 wl_90
* net 194 wl_91
* net 197 wl_92
* net 198 wl_93
* net 201 wl_95
* net 202 wl_94
* net 205 wl_96
* net 206 wl_97
* net 209 wl_98
* net 210 wl_99
* net 213 wl_101
* net 214 wl_100
* net 217 wl_102
* net 218 wl_103
* net 221 wl_105
* net 222 wl_104
* net 225 wl_106
* net 226 wl_107
* net 229 wl_108
* net 230 wl_109
* net 233 wl_110
* net 234 wl_111
* net 237 wl_113
* net 238 wl_112
* net 241 wl_114
* net 242 wl_115
* net 245 wl_117
* net 246 wl_116
* net 249 wl_118
* net 250 wl_119
* net 253 wl_121
* net 254 wl_120
* net 257 wl_123
* net 258 wl_122
* net 261 wl_125
* net 262 wl_124
* net 265 wl_127
* net 266 wl_126
* net 268 wl_128
* net 269 vdd
* net 270 gnd
* cell instance $1 r0 *1 10.68,0
X$1 4 5 3 9 7 8 6 11 10 15 13 14 12 18 16 19 17 21 20 22 23 25 24 34 36 38 35
+ 39 37 41 40 42 43 45 44 47 46 50 48 51 49 53 52 54 55 57 56 59 58 61 60 62 63
+ 64 65 66 68 69 67 70 72 73 71 74 76 77 75 78 80 81 79 82 84 85 83 86 88 89 87
+ 90 92 93 91 94 96 97 95 98 100 101 99 102 104 105 103 106 108 109 107 110 112
+ 113 111 114 116 117 115 118 120 121 119 122 124 125 123 126 128 129 127 130
+ 132 133 131 134 136 137 135 138 139 140 1 142 141 143 146 145 144 147 149 150
+ 148 151 154 153 152 155 157 158 156 159 162 161 160 163 165 166 164 167 169
+ 170 168 171 173 174 172 175 178 177 176 179 181 182 180 183 186 185 184 187
+ 189 190 188 191 193 194 192 195 197 198 196 199 202 201 200 203 205 206 204
+ 207 209 210 208 211 214 213 212 215 217 218 216 219 222 221 220 223 225 226
+ 224 227 229 230 228 231 233 234 232 235 238 237 236 239 241 242 240 243 246
+ 245 244 247 249 250 248 251 254 253 252 255 258 257 256 259 262 261 260 263
+ 266 265 264 267 268 269 270
+ freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver_array
* cell instance $3 m0 *1 11.24,0
X$3 2 1 269 269 270 freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec_0
* cell instance $4 r0 *1 0,0
X$4 3 4 7 26 27 13 6 10 16 12 29 28 17 23 20 30 31 32 33 24 36 35 37 40 44 43
+ 48 46 49 55 52 60 63 56 58 68 67 65 71 76 72 80 79 75 83 88 84 92 91 87 95 96
+ 100 104 103 99 107 108 112 116 115 111 119 124 120 128 127 123 131 132 136
+ 139 135 141 143 144 147 151 152 148 155 156 159 163 160 164 168 167 171 175
+ 176 172 179 180 183 187 184 188 192 191 195 199 196 200 204 203 207 212 211
+ 208 216 219 215 223 224 220 228 227 231 235 236 232 240 239 243 244 248 247
+ 252 255 251 259 260 256 264 263 267 269 270
+ freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_decoder
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_port_address

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_port_data
* pin rbl_bl
* pin rbl_br
* pin bl_0
* pin br_0
* pin bl_1
* pin bl_2
* pin br_2
* pin bl_3
* pin bl_4
* pin bl_5
* pin br_5
* pin bl_6
* pin bl_7
* pin br_7
* pin bl_8
* pin bl_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin bl_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin bl_23
* pin br_23
* pin bl_24
* pin bl_25
* pin br_25
* pin bl_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin bl_51
* pin br_51
* pin bl_52
* pin bl_53
* pin bl_54
* pin bl_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin bl_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin bl_107
* pin br_107
* pin bl_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin bl_128
* pin br_128
* pin bl_129
* pin br_129
* pin bl_130
* pin br_130
* pin bl_131
* pin br_131
* pin bl_132
* pin br_132
* pin bl_133
* pin br_133
* pin bl_134
* pin br_134
* pin bl_135
* pin br_135
* pin bl_136
* pin br_136
* pin bl_137
* pin br_137
* pin bl_138
* pin br_138
* pin bl_139
* pin br_139
* pin bl_140
* pin br_140
* pin bl_141
* pin br_141
* pin bl_142
* pin br_142
* pin bl_143
* pin br_143
* pin bl_144
* pin bl_145
* pin br_145
* pin bl_146
* pin br_146
* pin bl_147
* pin br_147
* pin bl_148
* pin br_148
* pin bl_149
* pin br_149
* pin bl_150
* pin br_150
* pin bl_151
* pin br_151
* pin bl_152
* pin br_152
* pin bl_153
* pin br_153
* pin bl_154
* pin br_154
* pin bl_155
* pin br_155
* pin bl_156
* pin br_156
* pin bl_157
* pin br_157
* pin bl_158
* pin br_158
* pin bl_159
* pin bl_160
* pin br_160
* pin bl_161
* pin br_161
* pin bl_162
* pin br_162
* pin bl_163
* pin br_163
* pin bl_164
* pin br_164
* pin bl_165
* pin br_165
* pin bl_166
* pin br_166
* pin bl_167
* pin br_167
* pin bl_168
* pin br_168
* pin bl_169
* pin br_169
* pin bl_170
* pin br_170
* pin bl_171
* pin br_171
* pin bl_172
* pin br_172
* pin bl_173
* pin bl_174
* pin br_174
* pin bl_175
* pin bl_176
* pin br_176
* pin bl_177
* pin br_177
* pin bl_178
* pin bl_179
* pin br_179
* pin bl_180
* pin br_180
* pin bl_181
* pin br_181
* pin bl_182
* pin br_182
* pin bl_183
* pin bl_184
* pin br_184
* pin bl_185
* pin br_185
* pin bl_186
* pin br_186
* pin bl_187
* pin bl_188
* pin br_188
* pin bl_189
* pin br_189
* pin bl_190
* pin br_190
* pin bl_191
* pin br_191
* pin bl_192
* pin br_192
* pin bl_193
* pin br_193
* pin bl_194
* pin br_194
* pin bl_195
* pin br_195
* pin bl_196
* pin br_196
* pin bl_197
* pin br_197
* pin bl_198
* pin br_198
* pin bl_199
* pin br_199
* pin bl_200
* pin br_200
* pin bl_201
* pin br_201
* pin bl_202
* pin br_202
* pin bl_203
* pin br_203
* pin bl_204
* pin br_204
* pin bl_205
* pin br_205
* pin bl_206
* pin br_206
* pin bl_207
* pin br_207
* pin bl_208
* pin br_208
* pin bl_209
* pin br_209
* pin bl_210
* pin br_210
* pin bl_211
* pin br_211
* pin bl_212
* pin br_212
* pin bl_213
* pin br_213
* pin bl_214
* pin br_214
* pin bl_215
* pin br_215
* pin bl_216
* pin br_216
* pin bl_217
* pin bl_218
* pin br_218
* pin bl_219
* pin br_219
* pin bl_220
* pin br_220
* pin bl_221
* pin br_221
* pin bl_222
* pin bl_223
* pin br_223
* pin bl_224
* pin br_224
* pin bl_225
* pin br_225
* pin bl_226
* pin bl_227
* pin br_227
* pin bl_228
* pin br_228
* pin bl_229
* pin bl_230
* pin br_230
* pin bl_231
* pin br_231
* pin bl_232
* pin br_232
* pin bl_233
* pin br_233
* pin bl_234
* pin br_234
* pin bl_235
* pin br_235
* pin bl_236
* pin br_236
* pin bl_237
* pin br_237
* pin bl_238
* pin br_238
* pin bl_239
* pin bl_240
* pin bl_241
* pin br_241
* pin bl_242
* pin br_242
* pin bl_243
* pin bl_244
* pin br_244
* pin bl_245
* pin bl_246
* pin bl_247
* pin bl_248
* pin bl_249
* pin br_249
* pin bl_250
* pin br_250
* pin bl_251
* pin bl_252
* pin br_252
* pin bl_253
* pin br_253
* pin bl_254
* pin br_254
* pin bl_255
* pin br_255
* pin sparebl_0
* pin sparebr_0
* pin br_1
* pin br_3
* pin br_4
* pin br_6
* pin br_8
* pin br_9
* pin br_16
* pin br_17
* pin br_22
* pin br_24
* pin br_26
* pin br_37
* pin br_50
* pin br_52
* pin br_53
* pin br_54
* pin br_55
* pin br_59
* pin br_74
* pin br_93
* pin br_98
* pin br_102
* pin br_103
* pin br_106
* pin br_108
* pin br_111
* pin br_115
* pin br_119
* pin br_122
* pin p_en_bar
* pin br_127
* pin br_144
* pin br_159
* pin br_173
* pin br_175
* pin br_178
* pin br_183
* pin br_187
* pin br_217
* pin br_222
* pin br_226
* pin br_229
* pin br_239
* pin br_240
* pin br_243
* pin br_245
* pin br_246
* pin br_247
* pin br_248
* pin br_251
* pin sel_7
* pin sel_6
* pin sel_5
* pin sel_4
* pin sel_3
* pin sel_2
* pin sel_1
* pin sel_0
* pin dout_0
* pin dout_1
* pin dout_2
* pin dout_3
* pin dout_4
* pin dout_5
* pin dout_6
* pin dout_7
* pin dout_8
* pin dout_9
* pin dout_10
* pin dout_11
* pin dout_12
* pin dout_13
* pin dout_14
* pin dout_15
* pin s_en
* pin dout_16
* pin dout_17
* pin dout_18
* pin dout_19
* pin dout_20
* pin dout_21
* pin dout_22
* pin dout_23
* pin dout_24
* pin dout_25
* pin dout_26
* pin dout_27
* pin dout_28
* pin dout_29
* pin dout_30
* pin dout_31
* pin dout_32
* pin din_0
* pin din_1
* pin din_2
* pin din_3
* pin din_4
* pin din_5
* pin din_6
* pin din_7
* pin din_8
* pin din_9
* pin din_10
* pin din_11
* pin din_12
* pin din_13
* pin din_14
* pin din_15
* pin w_en
* pin din_16
* pin din_17
* pin din_18
* pin din_19
* pin din_20
* pin din_21
* pin din_22
* pin din_23
* pin din_24
* pin din_25
* pin din_26
* pin din_27
* pin din_28
* pin din_29
* pin din_30
* pin din_31
* pin din_32
* pin bank_spare_wen0
* pin bank_wmask_0
* pin bank_wmask_1
* pin bank_wmask_2
* pin bank_wmask_3
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_port_data 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37
+ 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89
+ 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110 111
+ 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129 130
+ 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148 149
+ 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167 168
+ 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186 187
+ 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205 206
+ 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224 225
+ 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263
+ 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282
+ 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339
+ 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358
+ 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377
+ 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396
+ 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415
+ 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434
+ 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453
+ 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472
+ 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491
+ 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 590 591 592 593
+ 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610 611 612
+ 613 614 615 616 617 618 619 620 621 622 623 624 626 627 628 629 630 631 632
+ 633 635 636 637 638 639 640 641 642 643 645 646 647 648 649 650 651 652 654
+ 655 656 657 658 659 660 661 662 663 664 665 666 667 668
* net 1 rbl_bl
* net 2 rbl_br
* net 3 bl_0
* net 4 br_0
* net 5 bl_1
* net 6 bl_2
* net 7 br_2
* net 8 bl_3
* net 9 bl_4
* net 10 bl_5
* net 11 br_5
* net 12 bl_6
* net 13 bl_7
* net 14 br_7
* net 15 bl_8
* net 16 bl_9
* net 17 bl_10
* net 18 br_10
* net 19 bl_11
* net 20 br_11
* net 21 bl_12
* net 22 br_12
* net 23 bl_13
* net 24 br_13
* net 25 bl_14
* net 26 br_14
* net 27 bl_15
* net 28 br_15
* net 29 bl_16
* net 30 bl_17
* net 31 bl_18
* net 32 br_18
* net 33 bl_19
* net 34 br_19
* net 35 bl_20
* net 36 br_20
* net 37 bl_21
* net 38 br_21
* net 39 bl_22
* net 40 bl_23
* net 41 br_23
* net 42 bl_24
* net 43 bl_25
* net 44 br_25
* net 45 bl_26
* net 46 bl_27
* net 47 br_27
* net 48 bl_28
* net 49 br_28
* net 50 bl_29
* net 51 br_29
* net 52 bl_30
* net 53 br_30
* net 54 bl_31
* net 55 br_31
* net 56 bl_32
* net 57 br_32
* net 58 bl_33
* net 59 br_33
* net 60 bl_34
* net 61 br_34
* net 62 bl_35
* net 63 br_35
* net 64 bl_36
* net 65 br_36
* net 66 bl_37
* net 67 bl_38
* net 68 br_38
* net 69 bl_39
* net 70 br_39
* net 71 bl_40
* net 72 br_40
* net 73 bl_41
* net 74 br_41
* net 75 bl_42
* net 76 br_42
* net 77 bl_43
* net 78 br_43
* net 79 bl_44
* net 80 br_44
* net 81 bl_45
* net 82 br_45
* net 83 bl_46
* net 84 br_46
* net 85 bl_47
* net 86 br_47
* net 87 bl_48
* net 88 br_48
* net 89 bl_49
* net 90 br_49
* net 91 bl_50
* net 92 bl_51
* net 93 br_51
* net 94 bl_52
* net 95 bl_53
* net 96 bl_54
* net 97 bl_55
* net 98 bl_56
* net 99 br_56
* net 100 bl_57
* net 101 br_57
* net 102 bl_58
* net 103 br_58
* net 104 bl_59
* net 105 bl_60
* net 106 br_60
* net 107 bl_61
* net 108 br_61
* net 109 bl_62
* net 110 br_62
* net 111 bl_63
* net 112 br_63
* net 113 bl_64
* net 114 br_64
* net 115 bl_65
* net 116 br_65
* net 117 bl_66
* net 118 br_66
* net 119 bl_67
* net 120 br_67
* net 121 bl_68
* net 122 br_68
* net 123 bl_69
* net 124 br_69
* net 125 bl_70
* net 126 br_70
* net 127 bl_71
* net 128 br_71
* net 129 bl_72
* net 130 br_72
* net 131 bl_73
* net 132 br_73
* net 133 bl_74
* net 134 bl_75
* net 135 br_75
* net 136 bl_76
* net 137 br_76
* net 138 bl_77
* net 139 br_77
* net 140 bl_78
* net 141 br_78
* net 142 bl_79
* net 143 br_79
* net 144 bl_80
* net 145 br_80
* net 146 bl_81
* net 147 br_81
* net 148 bl_82
* net 149 br_82
* net 150 bl_83
* net 151 br_83
* net 152 bl_84
* net 153 br_84
* net 154 bl_85
* net 155 br_85
* net 156 bl_86
* net 157 br_86
* net 158 bl_87
* net 159 br_87
* net 160 bl_88
* net 161 br_88
* net 162 bl_89
* net 163 br_89
* net 164 bl_90
* net 165 br_90
* net 166 bl_91
* net 167 br_91
* net 168 bl_92
* net 169 br_92
* net 170 bl_93
* net 171 bl_94
* net 172 br_94
* net 173 bl_95
* net 174 br_95
* net 175 bl_96
* net 176 br_96
* net 177 bl_97
* net 178 br_97
* net 179 bl_98
* net 180 bl_99
* net 181 br_99
* net 182 bl_100
* net 183 br_100
* net 184 bl_101
* net 185 br_101
* net 186 bl_102
* net 187 bl_103
* net 188 bl_104
* net 189 br_104
* net 190 bl_105
* net 191 br_105
* net 192 bl_106
* net 193 bl_107
* net 194 br_107
* net 195 bl_108
* net 196 bl_109
* net 197 br_109
* net 198 bl_110
* net 199 br_110
* net 200 bl_111
* net 201 bl_112
* net 202 br_112
* net 203 bl_113
* net 204 br_113
* net 205 bl_114
* net 206 br_114
* net 207 bl_115
* net 208 bl_116
* net 209 br_116
* net 210 bl_117
* net 211 br_117
* net 212 bl_118
* net 213 br_118
* net 214 bl_119
* net 215 bl_120
* net 216 br_120
* net 217 bl_121
* net 218 br_121
* net 219 bl_122
* net 220 bl_123
* net 221 br_123
* net 222 bl_124
* net 223 br_124
* net 224 bl_125
* net 225 br_125
* net 226 bl_126
* net 227 br_126
* net 228 bl_127
* net 229 bl_128
* net 230 br_128
* net 231 bl_129
* net 232 br_129
* net 233 bl_130
* net 234 br_130
* net 235 bl_131
* net 236 br_131
* net 237 bl_132
* net 238 br_132
* net 239 bl_133
* net 240 br_133
* net 241 bl_134
* net 242 br_134
* net 243 bl_135
* net 244 br_135
* net 245 bl_136
* net 246 br_136
* net 247 bl_137
* net 248 br_137
* net 249 bl_138
* net 250 br_138
* net 251 bl_139
* net 252 br_139
* net 253 bl_140
* net 254 br_140
* net 255 bl_141
* net 256 br_141
* net 257 bl_142
* net 258 br_142
* net 259 bl_143
* net 260 br_143
* net 261 bl_144
* net 262 bl_145
* net 263 br_145
* net 264 bl_146
* net 265 br_146
* net 266 bl_147
* net 267 br_147
* net 268 bl_148
* net 269 br_148
* net 270 bl_149
* net 271 br_149
* net 272 bl_150
* net 273 br_150
* net 274 bl_151
* net 275 br_151
* net 276 bl_152
* net 277 br_152
* net 278 bl_153
* net 279 br_153
* net 280 bl_154
* net 281 br_154
* net 282 bl_155
* net 283 br_155
* net 284 bl_156
* net 285 br_156
* net 286 bl_157
* net 287 br_157
* net 288 bl_158
* net 289 br_158
* net 290 bl_159
* net 291 bl_160
* net 292 br_160
* net 293 bl_161
* net 294 br_161
* net 295 bl_162
* net 296 br_162
* net 297 bl_163
* net 298 br_163
* net 299 bl_164
* net 300 br_164
* net 301 bl_165
* net 302 br_165
* net 303 bl_166
* net 304 br_166
* net 305 bl_167
* net 306 br_167
* net 307 bl_168
* net 308 br_168
* net 309 bl_169
* net 310 br_169
* net 311 bl_170
* net 312 br_170
* net 313 bl_171
* net 314 br_171
* net 315 bl_172
* net 316 br_172
* net 317 bl_173
* net 318 bl_174
* net 319 br_174
* net 320 bl_175
* net 321 bl_176
* net 322 br_176
* net 323 bl_177
* net 324 br_177
* net 325 bl_178
* net 326 bl_179
* net 327 br_179
* net 328 bl_180
* net 329 br_180
* net 330 bl_181
* net 331 br_181
* net 332 bl_182
* net 333 br_182
* net 334 bl_183
* net 335 bl_184
* net 336 br_184
* net 337 bl_185
* net 338 br_185
* net 339 bl_186
* net 340 br_186
* net 341 bl_187
* net 342 bl_188
* net 343 br_188
* net 344 bl_189
* net 345 br_189
* net 346 bl_190
* net 347 br_190
* net 348 bl_191
* net 349 br_191
* net 350 bl_192
* net 351 br_192
* net 352 bl_193
* net 353 br_193
* net 354 bl_194
* net 355 br_194
* net 356 bl_195
* net 357 br_195
* net 358 bl_196
* net 359 br_196
* net 360 bl_197
* net 361 br_197
* net 362 bl_198
* net 363 br_198
* net 364 bl_199
* net 365 br_199
* net 366 bl_200
* net 367 br_200
* net 368 bl_201
* net 369 br_201
* net 370 bl_202
* net 371 br_202
* net 372 bl_203
* net 373 br_203
* net 374 bl_204
* net 375 br_204
* net 376 bl_205
* net 377 br_205
* net 378 bl_206
* net 379 br_206
* net 380 bl_207
* net 381 br_207
* net 382 bl_208
* net 383 br_208
* net 384 bl_209
* net 385 br_209
* net 386 bl_210
* net 387 br_210
* net 388 bl_211
* net 389 br_211
* net 390 bl_212
* net 391 br_212
* net 392 bl_213
* net 393 br_213
* net 394 bl_214
* net 395 br_214
* net 396 bl_215
* net 397 br_215
* net 398 bl_216
* net 399 br_216
* net 400 bl_217
* net 401 bl_218
* net 402 br_218
* net 403 bl_219
* net 404 br_219
* net 405 bl_220
* net 406 br_220
* net 407 bl_221
* net 408 br_221
* net 409 bl_222
* net 410 bl_223
* net 411 br_223
* net 412 bl_224
* net 413 br_224
* net 414 bl_225
* net 415 br_225
* net 416 bl_226
* net 417 bl_227
* net 418 br_227
* net 419 bl_228
* net 420 br_228
* net 421 bl_229
* net 422 bl_230
* net 423 br_230
* net 424 bl_231
* net 425 br_231
* net 426 bl_232
* net 427 br_232
* net 428 bl_233
* net 429 br_233
* net 430 bl_234
* net 431 br_234
* net 432 bl_235
* net 433 br_235
* net 434 bl_236
* net 435 br_236
* net 436 bl_237
* net 437 br_237
* net 438 bl_238
* net 439 br_238
* net 440 bl_239
* net 441 bl_240
* net 442 bl_241
* net 443 br_241
* net 444 bl_242
* net 445 br_242
* net 446 bl_243
* net 447 bl_244
* net 448 br_244
* net 449 bl_245
* net 450 bl_246
* net 451 bl_247
* net 452 bl_248
* net 453 bl_249
* net 454 br_249
* net 455 bl_250
* net 456 br_250
* net 457 bl_251
* net 458 bl_252
* net 459 br_252
* net 460 bl_253
* net 461 br_253
* net 462 bl_254
* net 463 br_254
* net 464 bl_255
* net 465 br_255
* net 466 sparebl_0
* net 467 sparebr_0
* net 468 br_1
* net 469 br_3
* net 470 br_4
* net 471 br_6
* net 472 br_8
* net 473 br_9
* net 474 br_16
* net 475 br_17
* net 476 br_22
* net 477 br_24
* net 478 br_26
* net 479 br_37
* net 480 br_50
* net 481 br_52
* net 482 br_53
* net 483 br_54
* net 484 br_55
* net 485 br_59
* net 486 br_74
* net 487 br_93
* net 488 br_98
* net 489 br_102
* net 490 br_103
* net 491 br_106
* net 492 br_108
* net 493 br_111
* net 494 br_115
* net 495 br_119
* net 496 br_122
* net 497 p_en_bar
* net 498 br_127
* net 499 br_144
* net 500 br_159
* net 501 br_173
* net 502 br_175
* net 503 br_178
* net 504 br_183
* net 505 br_187
* net 506 br_217
* net 507 br_222
* net 508 br_226
* net 509 br_229
* net 510 br_239
* net 511 br_240
* net 512 br_243
* net 513 br_245
* net 514 br_246
* net 515 br_247
* net 516 br_248
* net 517 br_251
* net 518 sel_7
* net 519 sel_6
* net 520 sel_5
* net 521 sel_4
* net 522 sel_3
* net 523 sel_2
* net 524 sel_1
* net 525 sel_0
* net 590 dout_0
* net 591 dout_1
* net 592 dout_2
* net 593 dout_3
* net 594 dout_4
* net 595 dout_5
* net 596 dout_6
* net 597 dout_7
* net 598 dout_8
* net 599 dout_9
* net 600 dout_10
* net 601 dout_11
* net 602 dout_12
* net 603 dout_13
* net 604 dout_14
* net 605 dout_15
* net 606 s_en
* net 607 dout_16
* net 608 dout_17
* net 609 dout_18
* net 610 dout_19
* net 611 dout_20
* net 612 dout_21
* net 613 dout_22
* net 614 dout_23
* net 615 dout_24
* net 616 dout_25
* net 617 dout_26
* net 618 dout_27
* net 619 dout_28
* net 620 dout_29
* net 621 dout_30
* net 622 dout_31
* net 623 dout_32
* net 624 din_0
* net 625 wdriver_sel_0
* net 626 din_1
* net 627 din_2
* net 628 din_3
* net 629 din_4
* net 630 din_5
* net 631 din_6
* net 632 din_7
* net 633 din_8
* net 634 wdriver_sel_1
* net 635 din_9
* net 636 din_10
* net 637 din_11
* net 638 din_12
* net 639 din_13
* net 640 din_14
* net 641 din_15
* net 642 w_en
* net 643 din_16
* net 644 wdriver_sel_2
* net 645 din_17
* net 646 din_18
* net 647 din_19
* net 648 din_20
* net 649 din_21
* net 650 din_22
* net 651 din_23
* net 652 din_24
* net 653 wdriver_sel_3
* net 654 din_25
* net 655 din_26
* net 656 din_27
* net 657 din_28
* net 658 din_29
* net 659 din_30
* net 660 din_31
* net 661 din_32
* net 662 bank_spare_wen0
* net 663 bank_wmask_0
* net 664 bank_wmask_1
* net 665 bank_wmask_2
* net 666 bank_wmask_3
* net 667 vdd
* net 668 gnd
* cell instance $1 m0 *1 0,1.845
X$1 497 1 2 3 4 5 468 6 7 8 469 9 470 10 11 12 471 13 14 15 472 16 473 17 18 19
+ 20 21 22 23 24 25 26 27 28 29 474 30 475 31 32 33 34 35 36 37 38 39 476 40 41
+ 42 477 43 44 45 478 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 479 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 480 92 93 94 481 95 482 96 483 97 484 98 99 100 101 102 103 104 485
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 486 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 487 171 172 173 174 175 176 177 178
+ 179 488 180 181 182 183 184 185 186 489 187 490 188 189 190 191 192 491 193
+ 194 195 492 196 197 198 199 200 493 201 202 203 204 205 206 207 494 208 209
+ 210 211 212 213 214 495 215 216 217 218 219 496 220 221 222 223 224 225 226
+ 227 228 498 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 499 262
+ 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 500 291 292 293 294 295 296 297 298 299
+ 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 501
+ 318 319 320 502 321 322 323 324 325 503 326 327 328 329 330 331 332 333 334
+ 504 335 336 337 338 339 340 341 505 342 343 344 345 346 347 348 349 350 351
+ 352 353 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370
+ 371 372 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389
+ 390 391 392 393 394 395 396 397 398 399 400 506 401 402 403 404 405 406 407
+ 408 409 507 410 411 412 413 414 415 416 508 417 418 419 420 421 509 422 423
+ 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 510 441
+ 511 442 443 444 445 446 512 447 448 449 513 450 514 451 515 452 516 453 454
+ 455 456 457 517 458 459 460 461 462 463 464 465 466 467 667
+ freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_array
* cell instance $2 m0 *1 0,5.58
X$2 557 556 555 554 553 552 551 550 549 548 547 546 545 544 526 543 542 541 540
+ 539 538 537 536 535 534 533 532 531 530 529 528 527 525 524 523 522 589 588
+ 587 558 586 585 584 559 583 582 581 560 580 579 578 577 561 576 575 574 562
+ 573 572 571 563 570 569 568 564 567 566 565 521 520 519 518 3 4 5 468 6 7 8
+ 469 9 470 10 11 12 471 13 14 15 472 16 473 17 18 19 20 21 22 23 24 25 26 27
+ 28 29 474 30 475 31 32 33 34 35 36 37 38 39 476 40 41 42 477 43 44 45 478 46
+ 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 479 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 480 92 93 94
+ 481 95 482 96 483 97 484 98 99 100 101 102 103 104 485 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 486 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 487 171 172 173 174 175 176 177 178 179 488 180 181 182
+ 183 184 185 186 489 187 490 188 189 190 191 192 491 193 194 195 492 196 197
+ 198 199 200 493 201 202 203 204 205 206 207 494 208 209 210 211 212 213 214
+ 495 215 216 217 218 219 496 220 221 222 223 224 225 226 227 228 498 229 230
+ 231 232 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249
+ 250 251 252 253 254 255 256 257 258 259 260 261 499 262 263 264 265 266 267
+ 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286
+ 287 288 289 290 500 291 292 293 294 295 296 297 298 299 300 301 302 303 304
+ 305 306 307 308 309 310 311 312 313 314 315 316 317 501 318 319 320 502 321
+ 322 323 324 325 503 326 327 328 329 330 331 332 333 334 504 335 336 337 338
+ 339 340 341 505 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356
+ 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375
+ 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394
+ 395 396 397 398 399 400 506 401 402 403 404 405 406 407 408 409 507 410 411
+ 412 413 414 415 416 508 417 418 419 420 421 509 422 423 424 425 426 427 428
+ 429 430 431 432 433 434 435 436 437 438 439 440 510 441 511 442 443 444 445
+ 446 512 447 448 449 513 450 514 451 515 452 516 453 454 455 456 457 517 458
+ 459 460 461 462 463 464 465 668
+ freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux_array
* cell instance $3 m0 *1 0,10.97
X$3 590 558 526 591 559 527 592 560 528 593 561 529 594 562 530 595 563 531 596
+ 564 532 597 565 533 598 566 534 599 567 535 600 568 536 601 569 537 602 570
+ 538 603 571 539 604 572 540 605 573 541 607 574 542 608 575 543 609 576 544
+ 610 577 545 611 578 546 612 579 547 613 580 548 614 581 549 615 582 550 616
+ 583 551 617 584 552 618 585 553 619 586 554 620 587 555 621 588 556 622 589
+ 557 623 466 467 606 667 668
+ freepdk45_sram_4kbytes_1rw_32x1024_8_sense_amp_array
* cell instance $4 m0 *1 0,15.65
X$4 624 626 627 628 629 630 631 632 633 635 636 637 638 639 640 641 643 645 646
+ 647 648 649 650 651 652 654 655 656 657 658 659 660 661 526 527 528 529 625
+ 530 531 532 533 534 535 536 537 634 538 539 540 541 542 543 544 545 644 546
+ 547 548 549 550 551 552 553 653 554 555 556 557 467 662 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 466 667 668
+ freepdk45_sram_4kbytes_1rw_32x1024_8_write_driver_array
* cell instance $5 m0 *1 0,17.975
X$5 625 634 644 653 663 664 665 666 642 667 668
+ freepdk45_sram_4kbytes_1rw_32x1024_8_write_mask_and_array
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_port_data

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_capped_replica_bitcell_array
* pin rbl_bl_0_0
* pin rbl_br_0_0
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin bl_0_2
* pin br_0_2
* pin bl_0_3
* pin br_0_3
* pin bl_0_4
* pin br_0_4
* pin bl_0_5
* pin br_0_5
* pin bl_0_6
* pin br_0_6
* pin bl_0_7
* pin br_0_7
* pin bl_0_8
* pin br_0_8
* pin bl_0_9
* pin br_0_9
* pin bl_0_10
* pin br_0_10
* pin bl_0_11
* pin br_0_11
* pin bl_0_12
* pin br_0_12
* pin bl_0_13
* pin br_0_13
* pin bl_0_14
* pin br_0_14
* pin bl_0_15
* pin br_0_15
* pin bl_0_16
* pin br_0_16
* pin bl_0_17
* pin br_0_17
* pin bl_0_18
* pin br_0_18
* pin bl_0_19
* pin br_0_19
* pin bl_0_20
* pin br_0_20
* pin bl_0_21
* pin br_0_21
* pin bl_0_22
* pin br_0_22
* pin bl_0_23
* pin br_0_23
* pin bl_0_24
* pin br_0_24
* pin bl_0_25
* pin br_0_25
* pin bl_0_26
* pin br_0_26
* pin bl_0_27
* pin br_0_27
* pin bl_0_28
* pin br_0_28
* pin bl_0_29
* pin br_0_29
* pin bl_0_30
* pin br_0_30
* pin bl_0_31
* pin br_0_31
* pin bl_0_32
* pin br_0_32
* pin bl_0_33
* pin br_0_33
* pin bl_0_34
* pin br_0_34
* pin bl_0_35
* pin br_0_35
* pin bl_0_36
* pin br_0_36
* pin bl_0_37
* pin br_0_37
* pin bl_0_38
* pin br_0_38
* pin bl_0_39
* pin br_0_39
* pin bl_0_40
* pin br_0_40
* pin bl_0_41
* pin br_0_41
* pin bl_0_42
* pin br_0_42
* pin bl_0_43
* pin br_0_43
* pin bl_0_44
* pin br_0_44
* pin bl_0_45
* pin br_0_45
* pin bl_0_46
* pin br_0_46
* pin bl_0_47
* pin br_0_47
* pin bl_0_48
* pin br_0_48
* pin bl_0_49
* pin br_0_49
* pin bl_0_50
* pin br_0_50
* pin bl_0_51
* pin br_0_51
* pin bl_0_52
* pin br_0_52
* pin bl_0_53
* pin br_0_53
* pin bl_0_54
* pin br_0_54
* pin bl_0_55
* pin br_0_55
* pin bl_0_56
* pin br_0_56
* pin bl_0_57
* pin br_0_57
* pin bl_0_58
* pin br_0_58
* pin bl_0_59
* pin br_0_59
* pin bl_0_60
* pin br_0_60
* pin bl_0_61
* pin br_0_61
* pin bl_0_62
* pin br_0_62
* pin bl_0_63
* pin br_0_63
* pin bl_0_64
* pin br_0_64
* pin bl_0_65
* pin br_0_65
* pin bl_0_66
* pin br_0_66
* pin bl_0_67
* pin br_0_67
* pin bl_0_68
* pin br_0_68
* pin bl_0_69
* pin br_0_69
* pin bl_0_70
* pin br_0_70
* pin bl_0_71
* pin br_0_71
* pin bl_0_72
* pin br_0_72
* pin bl_0_73
* pin br_0_73
* pin bl_0_74
* pin br_0_74
* pin bl_0_75
* pin br_0_75
* pin bl_0_76
* pin br_0_76
* pin bl_0_77
* pin br_0_77
* pin bl_0_78
* pin br_0_78
* pin bl_0_79
* pin br_0_79
* pin bl_0_80
* pin br_0_80
* pin bl_0_81
* pin br_0_81
* pin bl_0_82
* pin br_0_82
* pin bl_0_83
* pin br_0_83
* pin bl_0_84
* pin br_0_84
* pin bl_0_85
* pin br_0_85
* pin bl_0_86
* pin br_0_86
* pin bl_0_87
* pin br_0_87
* pin bl_0_88
* pin br_0_88
* pin bl_0_89
* pin br_0_89
* pin bl_0_90
* pin br_0_90
* pin bl_0_91
* pin br_0_91
* pin bl_0_92
* pin br_0_92
* pin bl_0_93
* pin br_0_93
* pin bl_0_94
* pin br_0_94
* pin bl_0_95
* pin br_0_95
* pin bl_0_96
* pin br_0_96
* pin bl_0_97
* pin br_0_97
* pin bl_0_98
* pin br_0_98
* pin bl_0_99
* pin br_0_99
* pin bl_0_100
* pin br_0_100
* pin bl_0_101
* pin br_0_101
* pin bl_0_102
* pin br_0_102
* pin bl_0_103
* pin br_0_103
* pin bl_0_104
* pin br_0_104
* pin bl_0_105
* pin br_0_105
* pin bl_0_106
* pin br_0_106
* pin bl_0_107
* pin br_0_107
* pin bl_0_108
* pin br_0_108
* pin bl_0_109
* pin br_0_109
* pin bl_0_110
* pin br_0_110
* pin bl_0_111
* pin br_0_111
* pin bl_0_112
* pin br_0_112
* pin bl_0_113
* pin br_0_113
* pin bl_0_114
* pin br_0_114
* pin bl_0_115
* pin br_0_115
* pin bl_0_116
* pin br_0_116
* pin bl_0_117
* pin br_0_117
* pin bl_0_118
* pin br_0_118
* pin bl_0_119
* pin br_0_119
* pin bl_0_120
* pin br_0_120
* pin bl_0_121
* pin br_0_121
* pin bl_0_122
* pin br_0_122
* pin bl_0_123
* pin br_0_123
* pin bl_0_124
* pin br_0_124
* pin bl_0_125
* pin br_0_125
* pin bl_0_126
* pin br_0_126
* pin bl_0_127
* pin br_0_127
* pin wl_0_60
* pin wl_0_49
* pin wl_0_6
* pin wl_0_12
* pin wl_0_58
* pin wl_0_57
* pin wl_0_56
* pin wl_0_55
* pin wl_0_54
* pin wl_0_11
* pin wl_0_53
* pin wl_0_29
* pin wl_0_52
* pin wl_0_10
* pin wl_0_51
* pin wl_0_37
* pin wl_0_30
* pin wl_0_48
* pin wl_0_50
* pin wl_0_7
* pin wl_0_8
* pin wl_0_26
* pin wl_0_21
* pin wl_0_20
* pin wl_0_22
* pin wl_0_23
* pin wl_0_19
* pin wl_0_24
* pin wl_0_25
* pin wl_0_18
* pin wl_0_17
* pin wl_0_59
* pin wl_0_16
* pin wl_0_27
* pin wl_0_15
* pin wl_0_14
* pin wl_0_63
* pin wl_0_13
* pin wl_0_28
* pin wl_0_62
* pin wl_0_61
* pin wl_0_9
* pin wl_0_0
* pin wl_0_47
* pin wl_0_3
* pin wl_0_2
* pin wl_0_32
* pin wl_0_46
* pin wl_0_1
* pin wl_0_45
* pin wl_0_33
* pin wl_0_43
* pin wl_0_44
* pin wl_0_42
* pin wl_0_34
* pin rbl_wl_0_0
* pin wl_0_41
* pin wl_0_35
* pin wl_0_40
* pin wl_0_36
* pin wl_0_39
* pin wl_0_38
* pin wl_0_31
* pin wl_0_4
* pin wl_0_5
* pin bl_0_128
* pin br_0_128
* pin bl_0_129
* pin br_0_129
* pin bl_0_130
* pin br_0_130
* pin bl_0_131
* pin br_0_131
* pin bl_0_132
* pin br_0_132
* pin bl_0_133
* pin br_0_133
* pin bl_0_134
* pin br_0_134
* pin bl_0_135
* pin br_0_135
* pin bl_0_136
* pin br_0_136
* pin bl_0_137
* pin br_0_137
* pin bl_0_138
* pin br_0_138
* pin bl_0_139
* pin br_0_139
* pin bl_0_140
* pin br_0_140
* pin bl_0_141
* pin br_0_141
* pin bl_0_142
* pin br_0_142
* pin bl_0_143
* pin br_0_143
* pin bl_0_144
* pin br_0_144
* pin bl_0_145
* pin br_0_145
* pin bl_0_146
* pin br_0_146
* pin bl_0_147
* pin br_0_147
* pin bl_0_148
* pin br_0_148
* pin bl_0_149
* pin br_0_149
* pin bl_0_150
* pin br_0_150
* pin bl_0_151
* pin br_0_151
* pin bl_0_152
* pin br_0_152
* pin bl_0_153
* pin br_0_153
* pin bl_0_154
* pin br_0_154
* pin bl_0_155
* pin br_0_155
* pin bl_0_156
* pin br_0_156
* pin bl_0_157
* pin br_0_157
* pin bl_0_158
* pin br_0_158
* pin bl_0_159
* pin br_0_159
* pin bl_0_160
* pin br_0_160
* pin bl_0_161
* pin br_0_161
* pin bl_0_162
* pin br_0_162
* pin bl_0_163
* pin br_0_163
* pin bl_0_164
* pin br_0_164
* pin bl_0_165
* pin br_0_165
* pin bl_0_166
* pin br_0_166
* pin bl_0_167
* pin br_0_167
* pin bl_0_168
* pin br_0_168
* pin bl_0_169
* pin br_0_169
* pin bl_0_170
* pin br_0_170
* pin bl_0_171
* pin br_0_171
* pin bl_0_172
* pin br_0_172
* pin bl_0_173
* pin br_0_173
* pin bl_0_174
* pin br_0_174
* pin bl_0_175
* pin br_0_175
* pin bl_0_176
* pin br_0_176
* pin bl_0_177
* pin br_0_177
* pin bl_0_178
* pin br_0_178
* pin bl_0_179
* pin br_0_179
* pin bl_0_180
* pin br_0_180
* pin bl_0_181
* pin br_0_181
* pin bl_0_182
* pin br_0_182
* pin bl_0_183
* pin br_0_183
* pin bl_0_184
* pin br_0_184
* pin bl_0_185
* pin br_0_185
* pin bl_0_186
* pin br_0_186
* pin bl_0_187
* pin br_0_187
* pin bl_0_188
* pin br_0_188
* pin bl_0_189
* pin br_0_189
* pin bl_0_190
* pin br_0_190
* pin bl_0_191
* pin br_0_191
* pin bl_0_192
* pin br_0_192
* pin bl_0_193
* pin br_0_193
* pin bl_0_194
* pin br_0_194
* pin bl_0_195
* pin br_0_195
* pin bl_0_196
* pin br_0_196
* pin bl_0_197
* pin br_0_197
* pin bl_0_198
* pin br_0_198
* pin bl_0_199
* pin br_0_199
* pin bl_0_200
* pin br_0_200
* pin bl_0_201
* pin br_0_201
* pin bl_0_202
* pin br_0_202
* pin bl_0_203
* pin br_0_203
* pin bl_0_204
* pin br_0_204
* pin bl_0_205
* pin br_0_205
* pin bl_0_206
* pin br_0_206
* pin bl_0_207
* pin br_0_207
* pin bl_0_208
* pin br_0_208
* pin bl_0_209
* pin br_0_209
* pin bl_0_210
* pin br_0_210
* pin bl_0_211
* pin br_0_211
* pin bl_0_212
* pin br_0_212
* pin bl_0_213
* pin br_0_213
* pin bl_0_214
* pin br_0_214
* pin bl_0_215
* pin br_0_215
* pin bl_0_216
* pin br_0_216
* pin bl_0_217
* pin br_0_217
* pin bl_0_218
* pin br_0_218
* pin bl_0_219
* pin br_0_219
* pin bl_0_220
* pin br_0_220
* pin bl_0_221
* pin br_0_221
* pin bl_0_222
* pin br_0_222
* pin bl_0_223
* pin br_0_223
* pin bl_0_224
* pin br_0_224
* pin bl_0_225
* pin br_0_225
* pin bl_0_226
* pin br_0_226
* pin bl_0_227
* pin br_0_227
* pin bl_0_228
* pin br_0_228
* pin bl_0_229
* pin br_0_229
* pin bl_0_230
* pin br_0_230
* pin bl_0_231
* pin br_0_231
* pin bl_0_232
* pin br_0_232
* pin bl_0_233
* pin br_0_233
* pin bl_0_234
* pin br_0_234
* pin bl_0_235
* pin br_0_235
* pin bl_0_236
* pin br_0_236
* pin bl_0_237
* pin br_0_237
* pin bl_0_238
* pin br_0_238
* pin bl_0_239
* pin br_0_239
* pin bl_0_240
* pin br_0_240
* pin bl_0_241
* pin br_0_241
* pin bl_0_242
* pin br_0_242
* pin bl_0_243
* pin br_0_243
* pin bl_0_244
* pin br_0_244
* pin bl_0_245
* pin br_0_245
* pin bl_0_246
* pin br_0_246
* pin bl_0_247
* pin br_0_247
* pin bl_0_248
* pin br_0_248
* pin bl_0_249
* pin br_0_249
* pin bl_0_250
* pin br_0_250
* pin bl_0_251
* pin br_0_251
* pin bl_0_252
* pin br_0_252
* pin bl_0_253
* pin br_0_253
* pin bl_0_254
* pin br_0_254
* pin bl_0_255
* pin br_0_255
* pin bl_0_256
* pin br_0_256
* pin wl_0_119
* pin wl_0_118
* pin wl_0_95
* pin wl_0_78
* pin wl_0_120
* pin wl_0_82
* pin wl_0_65
* pin wl_0_121
* pin wl_0_94
* pin wl_0_67
* pin wl_0_77
* pin wl_0_122
* pin wl_0_107
* pin wl_0_93
* pin wl_0_123
* pin wl_0_83
* pin wl_0_108
* pin wl_0_92
* pin wl_0_76
* pin wl_0_66
* pin wl_0_105
* pin wl_0_79
* pin wl_0_104
* pin wl_0_103
* pin wl_0_111
* pin wl_0_109
* pin wl_0_102
* pin wl_0_80
* pin wl_0_68
* pin wl_0_112
* pin wl_0_101
* pin wl_0_100
* pin wl_0_110
* pin wl_0_113
* pin wl_0_99
* pin wl_0_98
* pin wl_0_81
* pin wl_0_106
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_97
* pin wl_0_117
* pin wl_0_96
* pin wl_0_74
* pin wl_0_84
* pin wl_0_72
* pin wl_0_90
* pin wl_0_71
* pin wl_0_89
* pin wl_0_128
* pin wl_0_127
* pin wl_0_73
* pin wl_0_64
* pin wl_0_85
* pin wl_0_88
* pin wl_0_126
* pin wl_0_69
* pin wl_0_91
* pin wl_0_86
* pin wl_0_125
* pin wl_0_124
* pin wl_0_87
* pin wl_0_70
* pin wl_0_75
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_capped_replica_bitcell_array 1 2 3
+ 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31
+ 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57
+ 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
+ 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125
+ 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
+ 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258
+ 259 260 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277
+ 278 279 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296
+ 297 298 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315
+ 316 317 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334
+ 335 336 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353
+ 354 355 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372
+ 373 374 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391
+ 392 393 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410
+ 411 412 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429
+ 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448
+ 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467
+ 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486
+ 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505
+ 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524
+ 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543
+ 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581
+ 582 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600
+ 601 602 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619
+ 620 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 639 640 641 642 643 644 645 646 647 648
* net 1 rbl_bl_0_0
* net 2 rbl_br_0_0
* net 3 bl_0_0
* net 4 br_0_0
* net 5 bl_0_1
* net 6 br_0_1
* net 7 bl_0_2
* net 8 br_0_2
* net 9 bl_0_3
* net 10 br_0_3
* net 11 bl_0_4
* net 12 br_0_4
* net 13 bl_0_5
* net 14 br_0_5
* net 15 bl_0_6
* net 16 br_0_6
* net 17 bl_0_7
* net 18 br_0_7
* net 19 bl_0_8
* net 20 br_0_8
* net 21 bl_0_9
* net 22 br_0_9
* net 23 bl_0_10
* net 24 br_0_10
* net 25 bl_0_11
* net 26 br_0_11
* net 27 bl_0_12
* net 28 br_0_12
* net 29 bl_0_13
* net 30 br_0_13
* net 31 bl_0_14
* net 32 br_0_14
* net 33 bl_0_15
* net 34 br_0_15
* net 35 bl_0_16
* net 36 br_0_16
* net 37 bl_0_17
* net 38 br_0_17
* net 39 bl_0_18
* net 40 br_0_18
* net 41 bl_0_19
* net 42 br_0_19
* net 43 bl_0_20
* net 44 br_0_20
* net 45 bl_0_21
* net 46 br_0_21
* net 47 bl_0_22
* net 48 br_0_22
* net 49 bl_0_23
* net 50 br_0_23
* net 51 bl_0_24
* net 52 br_0_24
* net 53 bl_0_25
* net 54 br_0_25
* net 55 bl_0_26
* net 56 br_0_26
* net 57 bl_0_27
* net 58 br_0_27
* net 59 bl_0_28
* net 60 br_0_28
* net 61 bl_0_29
* net 62 br_0_29
* net 63 bl_0_30
* net 64 br_0_30
* net 65 bl_0_31
* net 66 br_0_31
* net 67 bl_0_32
* net 68 br_0_32
* net 69 bl_0_33
* net 70 br_0_33
* net 71 bl_0_34
* net 72 br_0_34
* net 73 bl_0_35
* net 74 br_0_35
* net 75 bl_0_36
* net 76 br_0_36
* net 77 bl_0_37
* net 78 br_0_37
* net 79 bl_0_38
* net 80 br_0_38
* net 81 bl_0_39
* net 82 br_0_39
* net 83 bl_0_40
* net 84 br_0_40
* net 85 bl_0_41
* net 86 br_0_41
* net 87 bl_0_42
* net 88 br_0_42
* net 89 bl_0_43
* net 90 br_0_43
* net 91 bl_0_44
* net 92 br_0_44
* net 93 bl_0_45
* net 94 br_0_45
* net 95 bl_0_46
* net 96 br_0_46
* net 97 bl_0_47
* net 98 br_0_47
* net 99 bl_0_48
* net 100 br_0_48
* net 101 bl_0_49
* net 102 br_0_49
* net 103 bl_0_50
* net 104 br_0_50
* net 105 bl_0_51
* net 106 br_0_51
* net 107 bl_0_52
* net 108 br_0_52
* net 109 bl_0_53
* net 110 br_0_53
* net 111 bl_0_54
* net 112 br_0_54
* net 113 bl_0_55
* net 114 br_0_55
* net 115 bl_0_56
* net 116 br_0_56
* net 117 bl_0_57
* net 118 br_0_57
* net 119 bl_0_58
* net 120 br_0_58
* net 121 bl_0_59
* net 122 br_0_59
* net 123 bl_0_60
* net 124 br_0_60
* net 125 bl_0_61
* net 126 br_0_61
* net 127 bl_0_62
* net 128 br_0_62
* net 129 bl_0_63
* net 130 br_0_63
* net 131 bl_0_64
* net 132 br_0_64
* net 133 bl_0_65
* net 134 br_0_65
* net 135 bl_0_66
* net 136 br_0_66
* net 137 bl_0_67
* net 138 br_0_67
* net 139 bl_0_68
* net 140 br_0_68
* net 141 bl_0_69
* net 142 br_0_69
* net 143 bl_0_70
* net 144 br_0_70
* net 145 bl_0_71
* net 146 br_0_71
* net 147 bl_0_72
* net 148 br_0_72
* net 149 bl_0_73
* net 150 br_0_73
* net 151 bl_0_74
* net 152 br_0_74
* net 153 bl_0_75
* net 154 br_0_75
* net 155 bl_0_76
* net 156 br_0_76
* net 157 bl_0_77
* net 158 br_0_77
* net 159 bl_0_78
* net 160 br_0_78
* net 161 bl_0_79
* net 162 br_0_79
* net 163 bl_0_80
* net 164 br_0_80
* net 165 bl_0_81
* net 166 br_0_81
* net 167 bl_0_82
* net 168 br_0_82
* net 169 bl_0_83
* net 170 br_0_83
* net 171 bl_0_84
* net 172 br_0_84
* net 173 bl_0_85
* net 174 br_0_85
* net 175 bl_0_86
* net 176 br_0_86
* net 177 bl_0_87
* net 178 br_0_87
* net 179 bl_0_88
* net 180 br_0_88
* net 181 bl_0_89
* net 182 br_0_89
* net 183 bl_0_90
* net 184 br_0_90
* net 185 bl_0_91
* net 186 br_0_91
* net 187 bl_0_92
* net 188 br_0_92
* net 189 bl_0_93
* net 190 br_0_93
* net 191 bl_0_94
* net 192 br_0_94
* net 193 bl_0_95
* net 194 br_0_95
* net 195 bl_0_96
* net 196 br_0_96
* net 197 bl_0_97
* net 198 br_0_97
* net 199 bl_0_98
* net 200 br_0_98
* net 201 bl_0_99
* net 202 br_0_99
* net 203 bl_0_100
* net 204 br_0_100
* net 205 bl_0_101
* net 206 br_0_101
* net 207 bl_0_102
* net 208 br_0_102
* net 209 bl_0_103
* net 210 br_0_103
* net 211 bl_0_104
* net 212 br_0_104
* net 213 bl_0_105
* net 214 br_0_105
* net 215 bl_0_106
* net 216 br_0_106
* net 217 bl_0_107
* net 218 br_0_107
* net 219 bl_0_108
* net 220 br_0_108
* net 221 bl_0_109
* net 222 br_0_109
* net 223 bl_0_110
* net 224 br_0_110
* net 225 bl_0_111
* net 226 br_0_111
* net 227 bl_0_112
* net 228 br_0_112
* net 229 bl_0_113
* net 230 br_0_113
* net 231 bl_0_114
* net 232 br_0_114
* net 233 bl_0_115
* net 234 br_0_115
* net 235 bl_0_116
* net 236 br_0_116
* net 237 bl_0_117
* net 238 br_0_117
* net 239 bl_0_118
* net 240 br_0_118
* net 241 bl_0_119
* net 242 br_0_119
* net 243 bl_0_120
* net 244 br_0_120
* net 245 bl_0_121
* net 246 br_0_121
* net 247 bl_0_122
* net 248 br_0_122
* net 249 bl_0_123
* net 250 br_0_123
* net 251 bl_0_124
* net 252 br_0_124
* net 253 bl_0_125
* net 254 br_0_125
* net 255 bl_0_126
* net 256 br_0_126
* net 257 bl_0_127
* net 258 br_0_127
* net 259 wl_0_60
* net 260 wl_0_49
* net 261 wl_0_6
* net 262 wl_0_12
* net 263 wl_0_58
* net 264 wl_0_57
* net 265 wl_0_56
* net 266 wl_0_55
* net 267 wl_0_54
* net 268 wl_0_11
* net 269 wl_0_53
* net 270 wl_0_29
* net 271 wl_0_52
* net 272 wl_0_10
* net 273 wl_0_51
* net 274 wl_0_37
* net 275 wl_0_30
* net 276 wl_0_48
* net 277 wl_0_50
* net 278 wl_0_7
* net 279 wl_0_8
* net 280 wl_0_26
* net 281 wl_0_21
* net 282 wl_0_20
* net 283 wl_0_22
* net 284 wl_0_23
* net 285 wl_0_19
* net 286 wl_0_24
* net 287 wl_0_25
* net 288 wl_0_18
* net 289 wl_0_17
* net 290 wl_0_59
* net 291 wl_0_16
* net 292 wl_0_27
* net 293 wl_0_15
* net 294 wl_0_14
* net 295 wl_0_63
* net 296 wl_0_13
* net 297 wl_0_28
* net 298 wl_0_62
* net 299 wl_0_61
* net 300 wl_0_9
* net 301 wl_0_0
* net 302 wl_0_47
* net 303 wl_0_3
* net 304 wl_0_2
* net 305 wl_0_32
* net 306 wl_0_46
* net 307 wl_0_1
* net 308 wl_0_45
* net 309 wl_0_33
* net 310 wl_0_43
* net 311 wl_0_44
* net 312 wl_0_42
* net 313 wl_0_34
* net 314 rbl_wl_0_0
* net 315 wl_0_41
* net 316 wl_0_35
* net 317 wl_0_40
* net 318 wl_0_36
* net 319 wl_0_39
* net 320 wl_0_38
* net 321 wl_0_31
* net 322 wl_0_4
* net 323 wl_0_5
* net 324 bl_0_128
* net 325 br_0_128
* net 326 bl_0_129
* net 327 br_0_129
* net 328 bl_0_130
* net 329 br_0_130
* net 330 bl_0_131
* net 331 br_0_131
* net 332 bl_0_132
* net 333 br_0_132
* net 334 bl_0_133
* net 335 br_0_133
* net 336 bl_0_134
* net 337 br_0_134
* net 338 bl_0_135
* net 339 br_0_135
* net 340 bl_0_136
* net 341 br_0_136
* net 342 bl_0_137
* net 343 br_0_137
* net 344 bl_0_138
* net 345 br_0_138
* net 346 bl_0_139
* net 347 br_0_139
* net 348 bl_0_140
* net 349 br_0_140
* net 350 bl_0_141
* net 351 br_0_141
* net 352 bl_0_142
* net 353 br_0_142
* net 354 bl_0_143
* net 355 br_0_143
* net 356 bl_0_144
* net 357 br_0_144
* net 358 bl_0_145
* net 359 br_0_145
* net 360 bl_0_146
* net 361 br_0_146
* net 362 bl_0_147
* net 363 br_0_147
* net 364 bl_0_148
* net 365 br_0_148
* net 366 bl_0_149
* net 367 br_0_149
* net 368 bl_0_150
* net 369 br_0_150
* net 370 bl_0_151
* net 371 br_0_151
* net 372 bl_0_152
* net 373 br_0_152
* net 374 bl_0_153
* net 375 br_0_153
* net 376 bl_0_154
* net 377 br_0_154
* net 378 bl_0_155
* net 379 br_0_155
* net 380 bl_0_156
* net 381 br_0_156
* net 382 bl_0_157
* net 383 br_0_157
* net 384 bl_0_158
* net 385 br_0_158
* net 386 bl_0_159
* net 387 br_0_159
* net 388 bl_0_160
* net 389 br_0_160
* net 390 bl_0_161
* net 391 br_0_161
* net 392 bl_0_162
* net 393 br_0_162
* net 394 bl_0_163
* net 395 br_0_163
* net 396 bl_0_164
* net 397 br_0_164
* net 398 bl_0_165
* net 399 br_0_165
* net 400 bl_0_166
* net 401 br_0_166
* net 402 bl_0_167
* net 403 br_0_167
* net 404 bl_0_168
* net 405 br_0_168
* net 406 bl_0_169
* net 407 br_0_169
* net 408 bl_0_170
* net 409 br_0_170
* net 410 bl_0_171
* net 411 br_0_171
* net 412 bl_0_172
* net 413 br_0_172
* net 414 bl_0_173
* net 415 br_0_173
* net 416 bl_0_174
* net 417 br_0_174
* net 418 bl_0_175
* net 419 br_0_175
* net 420 bl_0_176
* net 421 br_0_176
* net 422 bl_0_177
* net 423 br_0_177
* net 424 bl_0_178
* net 425 br_0_178
* net 426 bl_0_179
* net 427 br_0_179
* net 428 bl_0_180
* net 429 br_0_180
* net 430 bl_0_181
* net 431 br_0_181
* net 432 bl_0_182
* net 433 br_0_182
* net 434 bl_0_183
* net 435 br_0_183
* net 436 bl_0_184
* net 437 br_0_184
* net 438 bl_0_185
* net 439 br_0_185
* net 440 bl_0_186
* net 441 br_0_186
* net 442 bl_0_187
* net 443 br_0_187
* net 444 bl_0_188
* net 445 br_0_188
* net 446 bl_0_189
* net 447 br_0_189
* net 448 bl_0_190
* net 449 br_0_190
* net 450 bl_0_191
* net 451 br_0_191
* net 452 bl_0_192
* net 453 br_0_192
* net 454 bl_0_193
* net 455 br_0_193
* net 456 bl_0_194
* net 457 br_0_194
* net 458 bl_0_195
* net 459 br_0_195
* net 460 bl_0_196
* net 461 br_0_196
* net 462 bl_0_197
* net 463 br_0_197
* net 464 bl_0_198
* net 465 br_0_198
* net 466 bl_0_199
* net 467 br_0_199
* net 468 bl_0_200
* net 469 br_0_200
* net 470 bl_0_201
* net 471 br_0_201
* net 472 bl_0_202
* net 473 br_0_202
* net 474 bl_0_203
* net 475 br_0_203
* net 476 bl_0_204
* net 477 br_0_204
* net 478 bl_0_205
* net 479 br_0_205
* net 480 bl_0_206
* net 481 br_0_206
* net 482 bl_0_207
* net 483 br_0_207
* net 484 bl_0_208
* net 485 br_0_208
* net 486 bl_0_209
* net 487 br_0_209
* net 488 bl_0_210
* net 489 br_0_210
* net 490 bl_0_211
* net 491 br_0_211
* net 492 bl_0_212
* net 493 br_0_212
* net 494 bl_0_213
* net 495 br_0_213
* net 496 bl_0_214
* net 497 br_0_214
* net 498 bl_0_215
* net 499 br_0_215
* net 500 bl_0_216
* net 501 br_0_216
* net 502 bl_0_217
* net 503 br_0_217
* net 504 bl_0_218
* net 505 br_0_218
* net 506 bl_0_219
* net 507 br_0_219
* net 508 bl_0_220
* net 509 br_0_220
* net 510 bl_0_221
* net 511 br_0_221
* net 512 bl_0_222
* net 513 br_0_222
* net 514 bl_0_223
* net 515 br_0_223
* net 516 bl_0_224
* net 517 br_0_224
* net 518 bl_0_225
* net 519 br_0_225
* net 520 bl_0_226
* net 521 br_0_226
* net 522 bl_0_227
* net 523 br_0_227
* net 524 bl_0_228
* net 525 br_0_228
* net 526 bl_0_229
* net 527 br_0_229
* net 528 bl_0_230
* net 529 br_0_230
* net 530 bl_0_231
* net 531 br_0_231
* net 532 bl_0_232
* net 533 br_0_232
* net 534 bl_0_233
* net 535 br_0_233
* net 536 bl_0_234
* net 537 br_0_234
* net 538 bl_0_235
* net 539 br_0_235
* net 540 bl_0_236
* net 541 br_0_236
* net 542 bl_0_237
* net 543 br_0_237
* net 544 bl_0_238
* net 545 br_0_238
* net 546 bl_0_239
* net 547 br_0_239
* net 548 bl_0_240
* net 549 br_0_240
* net 550 bl_0_241
* net 551 br_0_241
* net 552 bl_0_242
* net 553 br_0_242
* net 554 bl_0_243
* net 555 br_0_243
* net 556 bl_0_244
* net 557 br_0_244
* net 558 bl_0_245
* net 559 br_0_245
* net 560 bl_0_246
* net 561 br_0_246
* net 562 bl_0_247
* net 563 br_0_247
* net 564 bl_0_248
* net 565 br_0_248
* net 566 bl_0_249
* net 567 br_0_249
* net 568 bl_0_250
* net 569 br_0_250
* net 570 bl_0_251
* net 571 br_0_251
* net 572 bl_0_252
* net 573 br_0_252
* net 574 bl_0_253
* net 575 br_0_253
* net 576 bl_0_254
* net 577 br_0_254
* net 578 bl_0_255
* net 579 br_0_255
* net 580 bl_0_256
* net 581 br_0_256
* net 582 wl_0_119
* net 583 wl_0_118
* net 584 wl_0_95
* net 585 wl_0_78
* net 586 wl_0_120
* net 587 wl_0_82
* net 588 wl_0_65
* net 589 wl_0_121
* net 590 wl_0_94
* net 591 wl_0_67
* net 592 wl_0_77
* net 593 wl_0_122
* net 594 wl_0_107
* net 595 wl_0_93
* net 596 wl_0_123
* net 597 wl_0_83
* net 598 wl_0_108
* net 599 wl_0_92
* net 600 wl_0_76
* net 601 wl_0_66
* net 602 wl_0_105
* net 603 wl_0_79
* net 604 wl_0_104
* net 605 wl_0_103
* net 606 wl_0_111
* net 607 wl_0_109
* net 608 wl_0_102
* net 609 wl_0_80
* net 610 wl_0_68
* net 611 wl_0_112
* net 612 wl_0_101
* net 613 wl_0_100
* net 614 wl_0_110
* net 615 wl_0_113
* net 616 wl_0_99
* net 617 wl_0_98
* net 618 wl_0_81
* net 619 wl_0_106
* net 620 wl_0_114
* net 621 wl_0_115
* net 622 wl_0_116
* net 623 wl_0_97
* net 624 wl_0_117
* net 625 wl_0_96
* net 626 wl_0_74
* net 627 wl_0_84
* net 628 wl_0_72
* net 629 wl_0_90
* net 630 wl_0_71
* net 631 wl_0_89
* net 632 wl_0_128
* net 633 wl_0_127
* net 634 wl_0_73
* net 635 wl_0_64
* net 636 wl_0_85
* net 637 wl_0_88
* net 638 wl_0_126
* net 639 wl_0_69
* net 640 wl_0_91
* net 641 wl_0_86
* net 642 wl_0_125
* net 643 wl_0_124
* net 644 wl_0_87
* net 645 wl_0_70
* net 646 wl_0_75
* net 647 vdd
* net 648 gnd
* cell instance $1 r0 *1 1.64,0.25
X$1 648 647 648 freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_1
* cell instance $2 r0 *1 1.64,1.615
X$2 314 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27
+ 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53
+ 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79
+ 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179
+ 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198
+ 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217
+ 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236
+ 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255
+ 256 257 258 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339
+ 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358
+ 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377
+ 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396
+ 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415
+ 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433 434
+ 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452 453
+ 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471 472
+ 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490 491
+ 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509 510
+ 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528 529
+ 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547 548
+ 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566 567
+ 568 569 570 571 572 573 574 575 576 577 578 579 580 581 301 307 304 303 322
+ 323 261 278 279 300 272 268 262 296 294 293 291 289 288 285 282 281 283 284
+ 286 287 280 292 297 270 275 321 305 309 313 316 318 274 320 319 317 315 312
+ 310 311 308 306 302 276 260 277 273 271 269 267 266 265 264 263 290 259 299
+ 298 295 635 588 601 591 610 639 645 630 628 634 626 646 600 592 585 603 609
+ 618 587 597 627 636 641 644 637 631 629 640 599 595 590 584 625 623 617 616
+ 613 612 608 605 604 602 619 594 598 607 614 606 611 615 620 621 622 624 583
+ 582 586 589 593 596 643 642 638 633 632 647 648
+ freepdk45_sram_4kbytes_1rw_32x1024_8_replica_bitcell_array
* cell instance $3 m0 *1 1.64,180.43
X$3 648 647 648 freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_0
* cell instance $4 r0 *1 0.935,0.25
X$4 648 314 301 307 304 303 322 323 261 278 279 300 272 268 262 296 294 293 291
+ 289 288 285 282 281 283 284 286 287 280 292 297 270 275 321 305 309 313 316
+ 318 274 320 319 317 315 312 310 311 308 306 302 276 260 277 273 271 269 267
+ 266 265 264 263 290 259 299 298 295 635 588 601 591 610 639 645 630 628 634
+ 626 646 600 592 585 603 609 618 587 597 627 636 641 644 637 631 629 640 599
+ 595 590 584 625 623 617 616 613 612 608 605 604 602 619 594 598 607 614 606
+ 611 615 620 621 622 624 583 582 586 589 593 596 643 642 638 633 632 648 647
+ 648 freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_2
* cell instance $5 r0 *1 183.53,0.25
X$5 648 314 301 307 304 303 322 323 261 278 279 300 272 268 262 296 294 293 291
+ 289 288 285 282 281 283 284 286 287 280 292 297 270 275 321 305 309 313 316
+ 318 274 320 319 317 315 312 310 311 308 306 302 276 260 277 273 271 269 267
+ 266 265 264 263 290 259 299 298 295 635 588 601 591 610 639 645 630 628 634
+ 626 646 600 592 585 603 609 618 587 597 627 636 641 644 637 631 629 640 599
+ 595 590 584 625 623 617 616 613 612 608 605 604 602 619 594 598 607 614 606
+ 611 615 620 621 622 624 583 582 586 589 593 596 643 642 638 633 632 648 647
+ 648 freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_3
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_capped_replica_bitcell_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_0
* pin Qb
* pin Q
* pin clk
* pin D
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_0 1 2 4 5 6 7
* net 1 Qb
* net 2 Q
* net 4 clk
* net 5 D
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 3.195,0
X$1 3 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_4
* cell instance $2 r0 *1 3.8825,0
X$2 1 2 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_5
* cell instance $5 r0 *1 0,0
X$5 3 5 4 6 7 dff
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dff_buf_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_1
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_1 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_6
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_1

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_1
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_1 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_1

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_19
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_19 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2735 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=7.735U AS=0.87465P AD=0.87465P PS=13.9125U
+ PD=13.9125U
* device instance $27 r0 *1 0.2325,1.8985 PMOS_VTG
M$27 3 1 2 3 PMOS_VTG L=0.05U W=23.205U AS=2.62395P AD=2.62395P PS=29.9775U
+ PD=29.9775U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_19

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_18
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_18 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.27 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.61U AS=0.297975P AD=0.297975P PS=4.955U
+ PD=4.955U
* device instance $10 r0 *1 0.2325,1.91 PMOS_VTG
M$10 3 1 2 3 PMOS_VTG L=0.05U W=7.83U AS=0.893925P AD=0.893925P PS=10.755U
+ PD=10.755U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_18

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_17
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_17 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.275 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.9U AS=0.10575P AD=0.10575P PS=1.905U PD=1.905U
* device instance $4 r0 *1 0.2325,1.895 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=2.7U AS=0.31725P AD=0.31725P PS=4.305U PD=4.305U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_17

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_20

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_5
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_5 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_16
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_5

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_4
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_4 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_15
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_4

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_14
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_14 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2735 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=3.8675U AS=0.43955625P AD=0.43955625P PS=7.12U
+ PD=7.12U
* device instance $14 r0 *1 0.2325,1.8985 PMOS_VTG
M$14 3 1 2 3 PMOS_VTG L=0.05U W=11.6025U AS=1.31866875P AD=1.31866875P
+ PS=15.45U PD=15.45U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_14

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_13
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_13 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.251 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.2625U AS=0.14581875P AD=0.14581875P PS=2.67U
+ PD=2.67U
* device instance $6 r0 *1 0.2325,1.9675 PMOS_VTG
M$6 3 1 2 3 PMOS_VTG L=0.05U W=3.775U AS=0.4360125P AD=0.4360125P PS=5.685U
+ PD=5.685U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_13

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_12
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_12 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2785 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=7.38U AS=0.8348625P AD=0.8348625P PS=13.1175U
+ PD=13.1175U
* device instance $25 r0 *1 0.2325,1.8835 PMOS_VTG
M$25 3 1 2 3 PMOS_VTG L=0.05U W=22.14U AS=2.5045875P AD=2.5045875P PS=28.4925U
+ PD=28.4925U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_12

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_11
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_11 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2775 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.44U AS=0.279075P AD=0.279075P PS=4.575U
+ PD=4.575U
* device instance $9 r0 *1 0.2325,1.89 PMOS_VTG
M$9 3 1 2 3 PMOS_VTG L=0.05U W=7.28U AS=0.83265P AD=0.83265P PS=10.02U PD=10.02U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_11

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_10
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_10 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.81U AS=0.095175P AD=0.095175P PS=1.785U
+ PD=1.785U
* device instance $4 r0 *1 0.2325,1.94 PMOS_VTG
M$4 3 1 2 3 PMOS_VTG L=0.05U W=2.43U AS=0.285525P AD=0.285525P PS=3.945U
+ PD=3.945U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_10

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_9
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_9 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
* device instance $2 r0 *1 0.2325,1.94 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.81U AS=0.103275P AD=0.103275P PS=1.875U
+ PD=1.875U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_9

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8_0
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin in_2
* pin out_2
* pin out_3
* pin out_5
* pin out_4
* pin out_6
* pin out_7
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8_0 1 5 6
+ 7 8 9 10 11 12 13 14 15 16
* net 1 in_0
* net 5 in_1
* net 6 out_0
* net 7 out_1
* net 8 in_2
* net 9 out_2
* net 10 out_3
* net 11 out_5
* net 12 out_4
* net 13 out_6
* net 14 out_7
* net 15 vdd
* net 16 gnd
* cell instance $1 r0 *1 0.7,0
X$1 1 2 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
* cell instance $2 m0 *1 2.5075,19.76
X$2 14 1 5 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $3 m0 *1 2.5075,4.94
X$3 7 1 3 4 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $4 m0 *1 2.5075,9.88
X$4 10 1 5 4 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $5 m0 *1 2.5075,14.82
X$5 11 1 3 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $13 r0 *1 2.5075,0
X$13 6 2 3 4 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $14 r0 *1 2.5075,14.82
X$14 13 2 5 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $15 r0 *1 2.5075,4.94
X$15 9 2 5 4 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $16 r0 *1 2.5075,9.88
X$16 12 2 3 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* cell instance $22 m0 *1 0.7,4.94
X$22 5 3 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
* cell instance $28 r0 *1 0.7,4.94
X$28 8 4 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec_0
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec_0 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.9025,0
X$1 1 2 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_0
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver_array
* pin in_0
* pin wl_0
* pin in_1
* pin wl_1
* pin in_2
* pin wl_2
* pin in_3
* pin wl_3
* pin in_4
* pin wl_4
* pin in_5
* pin wl_5
* pin in_6
* pin wl_6
* pin in_7
* pin wl_7
* pin in_8
* pin wl_8
* pin in_9
* pin wl_9
* pin in_10
* pin wl_10
* pin in_11
* pin wl_11
* pin in_12
* pin wl_12
* pin in_13
* pin wl_13
* pin in_14
* pin wl_14
* pin in_15
* pin wl_15
* pin in_16
* pin wl_16
* pin in_17
* pin wl_17
* pin in_18
* pin wl_18
* pin in_19
* pin wl_19
* pin in_20
* pin wl_20
* pin in_21
* pin wl_21
* pin in_22
* pin wl_22
* pin in_23
* pin wl_23
* pin in_24
* pin wl_24
* pin in_25
* pin wl_25
* pin in_26
* pin wl_26
* pin in_27
* pin wl_27
* pin in_28
* pin wl_28
* pin in_29
* pin wl_29
* pin in_30
* pin wl_30
* pin in_31
* pin wl_31
* pin in_32
* pin wl_32
* pin in_33
* pin wl_33
* pin in_34
* pin wl_34
* pin in_35
* pin wl_35
* pin in_36
* pin wl_36
* pin in_37
* pin wl_37
* pin in_38
* pin wl_38
* pin in_39
* pin wl_39
* pin in_40
* pin wl_40
* pin in_41
* pin wl_41
* pin in_42
* pin wl_42
* pin in_43
* pin wl_43
* pin in_44
* pin wl_44
* pin in_45
* pin wl_45
* pin in_46
* pin wl_46
* pin in_47
* pin wl_47
* pin in_48
* pin wl_48
* pin in_49
* pin wl_49
* pin in_50
* pin wl_50
* pin in_51
* pin wl_51
* pin in_52
* pin wl_52
* pin in_53
* pin wl_53
* pin in_54
* pin wl_54
* pin in_55
* pin wl_55
* pin in_56
* pin wl_56
* pin in_57
* pin wl_57
* pin in_58
* pin wl_58
* pin in_59
* pin wl_59
* pin in_60
* pin wl_60
* pin in_61
* pin wl_61
* pin in_62
* pin wl_62
* pin in_63
* pin wl_63
* pin in_64
* pin wl_64
* pin en
* pin wl_65
* pin in_65
* pin in_66
* pin wl_66
* pin wl_67
* pin in_67
* pin in_68
* pin wl_68
* pin wl_69
* pin in_69
* pin in_70
* pin wl_70
* pin wl_71
* pin in_71
* pin in_72
* pin wl_72
* pin wl_73
* pin in_73
* pin in_74
* pin wl_74
* pin wl_75
* pin in_75
* pin in_76
* pin wl_76
* pin wl_77
* pin in_77
* pin in_78
* pin wl_78
* pin wl_79
* pin in_79
* pin in_80
* pin wl_80
* pin wl_81
* pin in_81
* pin in_82
* pin wl_82
* pin wl_83
* pin in_83
* pin in_84
* pin wl_84
* pin wl_85
* pin in_85
* pin in_86
* pin wl_86
* pin wl_87
* pin in_87
* pin in_88
* pin wl_88
* pin wl_89
* pin in_89
* pin in_90
* pin wl_90
* pin wl_91
* pin in_91
* pin in_92
* pin wl_92
* pin wl_93
* pin in_93
* pin in_94
* pin wl_94
* pin wl_95
* pin in_95
* pin in_96
* pin wl_96
* pin wl_97
* pin in_97
* pin in_98
* pin wl_98
* pin wl_99
* pin in_99
* pin in_100
* pin wl_100
* pin wl_101
* pin in_101
* pin in_102
* pin wl_102
* pin wl_103
* pin in_103
* pin in_104
* pin wl_104
* pin wl_105
* pin in_105
* pin in_106
* pin wl_106
* pin wl_107
* pin in_107
* pin in_108
* pin wl_108
* pin wl_109
* pin in_109
* pin in_110
* pin wl_110
* pin wl_111
* pin in_111
* pin in_112
* pin wl_112
* pin wl_113
* pin in_113
* pin in_114
* pin wl_114
* pin wl_115
* pin in_115
* pin in_116
* pin wl_116
* pin wl_117
* pin in_117
* pin in_118
* pin wl_118
* pin wl_119
* pin in_119
* pin in_120
* pin wl_120
* pin wl_121
* pin in_121
* pin in_122
* pin wl_122
* pin wl_123
* pin in_123
* pin in_124
* pin wl_124
* pin wl_125
* pin in_125
* pin in_126
* pin wl_126
* pin wl_127
* pin in_127
* pin in_128
* pin wl_128
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver_array 1 2 3 4 5 6
+ 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33
+ 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85
+ 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261
* net 1 in_0
* net 2 wl_0
* net 3 in_1
* net 4 wl_1
* net 5 in_2
* net 6 wl_2
* net 7 in_3
* net 8 wl_3
* net 9 in_4
* net 10 wl_4
* net 11 in_5
* net 12 wl_5
* net 13 in_6
* net 14 wl_6
* net 15 in_7
* net 16 wl_7
* net 17 in_8
* net 18 wl_8
* net 19 in_9
* net 20 wl_9
* net 21 in_10
* net 22 wl_10
* net 23 in_11
* net 24 wl_11
* net 25 in_12
* net 26 wl_12
* net 27 in_13
* net 28 wl_13
* net 29 in_14
* net 30 wl_14
* net 31 in_15
* net 32 wl_15
* net 33 in_16
* net 34 wl_16
* net 35 in_17
* net 36 wl_17
* net 37 in_18
* net 38 wl_18
* net 39 in_19
* net 40 wl_19
* net 41 in_20
* net 42 wl_20
* net 43 in_21
* net 44 wl_21
* net 45 in_22
* net 46 wl_22
* net 47 in_23
* net 48 wl_23
* net 49 in_24
* net 50 wl_24
* net 51 in_25
* net 52 wl_25
* net 53 in_26
* net 54 wl_26
* net 55 in_27
* net 56 wl_27
* net 57 in_28
* net 58 wl_28
* net 59 in_29
* net 60 wl_29
* net 61 in_30
* net 62 wl_30
* net 63 in_31
* net 64 wl_31
* net 65 in_32
* net 66 wl_32
* net 67 in_33
* net 68 wl_33
* net 69 in_34
* net 70 wl_34
* net 71 in_35
* net 72 wl_35
* net 73 in_36
* net 74 wl_36
* net 75 in_37
* net 76 wl_37
* net 77 in_38
* net 78 wl_38
* net 79 in_39
* net 80 wl_39
* net 81 in_40
* net 82 wl_40
* net 83 in_41
* net 84 wl_41
* net 85 in_42
* net 86 wl_42
* net 87 in_43
* net 88 wl_43
* net 89 in_44
* net 90 wl_44
* net 91 in_45
* net 92 wl_45
* net 93 in_46
* net 94 wl_46
* net 95 in_47
* net 96 wl_47
* net 97 in_48
* net 98 wl_48
* net 99 in_49
* net 100 wl_49
* net 101 in_50
* net 102 wl_50
* net 103 in_51
* net 104 wl_51
* net 105 in_52
* net 106 wl_52
* net 107 in_53
* net 108 wl_53
* net 109 in_54
* net 110 wl_54
* net 111 in_55
* net 112 wl_55
* net 113 in_56
* net 114 wl_56
* net 115 in_57
* net 116 wl_57
* net 117 in_58
* net 118 wl_58
* net 119 in_59
* net 120 wl_59
* net 121 in_60
* net 122 wl_60
* net 123 in_61
* net 124 wl_61
* net 125 in_62
* net 126 wl_62
* net 127 in_63
* net 128 wl_63
* net 129 in_64
* net 130 wl_64
* net 131 en
* net 132 wl_65
* net 133 in_65
* net 134 in_66
* net 135 wl_66
* net 136 wl_67
* net 137 in_67
* net 138 in_68
* net 139 wl_68
* net 140 wl_69
* net 141 in_69
* net 142 in_70
* net 143 wl_70
* net 144 wl_71
* net 145 in_71
* net 146 in_72
* net 147 wl_72
* net 148 wl_73
* net 149 in_73
* net 150 in_74
* net 151 wl_74
* net 152 wl_75
* net 153 in_75
* net 154 in_76
* net 155 wl_76
* net 156 wl_77
* net 157 in_77
* net 158 in_78
* net 159 wl_78
* net 160 wl_79
* net 161 in_79
* net 162 in_80
* net 163 wl_80
* net 164 wl_81
* net 165 in_81
* net 166 in_82
* net 167 wl_82
* net 168 wl_83
* net 169 in_83
* net 170 in_84
* net 171 wl_84
* net 172 wl_85
* net 173 in_85
* net 174 in_86
* net 175 wl_86
* net 176 wl_87
* net 177 in_87
* net 178 in_88
* net 179 wl_88
* net 180 wl_89
* net 181 in_89
* net 182 in_90
* net 183 wl_90
* net 184 wl_91
* net 185 in_91
* net 186 in_92
* net 187 wl_92
* net 188 wl_93
* net 189 in_93
* net 190 in_94
* net 191 wl_94
* net 192 wl_95
* net 193 in_95
* net 194 in_96
* net 195 wl_96
* net 196 wl_97
* net 197 in_97
* net 198 in_98
* net 199 wl_98
* net 200 wl_99
* net 201 in_99
* net 202 in_100
* net 203 wl_100
* net 204 wl_101
* net 205 in_101
* net 206 in_102
* net 207 wl_102
* net 208 wl_103
* net 209 in_103
* net 210 in_104
* net 211 wl_104
* net 212 wl_105
* net 213 in_105
* net 214 in_106
* net 215 wl_106
* net 216 wl_107
* net 217 in_107
* net 218 in_108
* net 219 wl_108
* net 220 wl_109
* net 221 in_109
* net 222 in_110
* net 223 wl_110
* net 224 wl_111
* net 225 in_111
* net 226 in_112
* net 227 wl_112
* net 228 wl_113
* net 229 in_113
* net 230 in_114
* net 231 wl_114
* net 232 wl_115
* net 233 in_115
* net 234 in_116
* net 235 wl_116
* net 236 wl_117
* net 237 in_117
* net 238 in_118
* net 239 wl_118
* net 240 wl_119
* net 241 in_119
* net 242 in_120
* net 243 wl_120
* net 244 wl_121
* net 245 in_121
* net 246 in_122
* net 247 wl_122
* net 248 wl_123
* net 249 in_123
* net 250 in_124
* net 251 wl_124
* net 252 wl_125
* net 253 in_125
* net 254 in_126
* net 255 wl_126
* net 256 wl_127
* net 257 in_127
* net 258 in_128
* net 259 wl_128
* net 260 vdd
* net 261 gnd
* cell instance $1 r0 *1 0.56,0
X$1 2 1 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $2 m0 *1 0.56,2.73
X$2 4 3 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $3 r0 *1 0.56,2.73
X$3 6 5 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $4 m0 *1 0.56,5.46
X$4 8 7 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $5 r0 *1 0.56,5.46
X$5 10 9 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $6 m0 *1 0.56,8.19
X$6 12 11 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $7 r0 *1 0.56,8.19
X$7 14 13 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $8 m0 *1 0.56,10.92
X$8 16 15 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $9 r0 *1 0.56,10.92
X$9 18 17 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $10 m0 *1 0.56,13.65
X$10 20 19 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $11 r0 *1 0.56,13.65
X$11 22 21 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $12 m0 *1 0.56,16.38
X$12 24 23 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $13 r0 *1 0.56,16.38
X$13 26 25 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $14 m0 *1 0.56,19.11
X$14 28 27 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $15 r0 *1 0.56,19.11
X$15 30 29 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $16 m0 *1 0.56,21.84
X$16 32 31 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $17 r0 *1 0.56,21.84
X$17 34 33 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $18 m0 *1 0.56,24.57
X$18 36 35 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $19 r0 *1 0.56,24.57
X$19 38 37 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $20 m0 *1 0.56,27.3
X$20 40 39 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $21 r0 *1 0.56,27.3
X$21 42 41 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $22 m0 *1 0.56,30.03
X$22 44 43 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $23 r0 *1 0.56,30.03
X$23 46 45 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $24 m0 *1 0.56,32.76
X$24 48 47 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $25 r0 *1 0.56,32.76
X$25 50 49 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $26 m0 *1 0.56,35.49
X$26 52 51 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $27 r0 *1 0.56,35.49
X$27 54 53 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $28 m0 *1 0.56,38.22
X$28 56 55 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $29 r0 *1 0.56,38.22
X$29 58 57 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $30 m0 *1 0.56,40.95
X$30 60 59 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $31 r0 *1 0.56,40.95
X$31 62 61 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $32 m0 *1 0.56,43.68
X$32 64 63 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $33 r0 *1 0.56,43.68
X$33 66 65 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $34 m0 *1 0.56,46.41
X$34 68 67 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $35 r0 *1 0.56,46.41
X$35 70 69 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $36 m0 *1 0.56,49.14
X$36 72 71 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $37 r0 *1 0.56,49.14
X$37 74 73 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $38 m0 *1 0.56,51.87
X$38 76 75 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $39 r0 *1 0.56,51.87
X$39 78 77 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $40 m0 *1 0.56,54.6
X$40 80 79 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $41 r0 *1 0.56,54.6
X$41 82 81 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $42 m0 *1 0.56,57.33
X$42 84 83 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $43 r0 *1 0.56,57.33
X$43 86 85 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $44 m0 *1 0.56,60.06
X$44 88 87 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $45 r0 *1 0.56,60.06
X$45 90 89 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $46 m0 *1 0.56,62.79
X$46 92 91 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $47 r0 *1 0.56,62.79
X$47 94 93 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $48 m0 *1 0.56,65.52
X$48 96 95 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $49 r0 *1 0.56,65.52
X$49 98 97 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $50 m0 *1 0.56,68.25
X$50 100 99 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $51 r0 *1 0.56,68.25
X$51 102 101 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $52 m0 *1 0.56,70.98
X$52 104 103 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $53 r0 *1 0.56,70.98
X$53 106 105 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $54 m0 *1 0.56,73.71
X$54 108 107 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $55 r0 *1 0.56,73.71
X$55 110 109 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $56 m0 *1 0.56,76.44
X$56 112 111 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $57 r0 *1 0.56,76.44
X$57 114 113 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $58 m0 *1 0.56,79.17
X$58 116 115 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $59 r0 *1 0.56,79.17
X$59 118 117 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $60 m0 *1 0.56,81.9
X$60 120 119 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $61 r0 *1 0.56,81.9
X$61 122 121 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $62 m0 *1 0.56,84.63
X$62 124 123 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $63 r0 *1 0.56,84.63
X$63 126 125 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $64 m0 *1 0.56,87.36
X$64 128 127 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $65 r0 *1 0.56,87.36
X$65 130 129 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $67 m0 *1 0.56,166.53
X$67 244 245 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $69 m0 *1 0.56,139.23
X$69 204 205 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $71 r0 *1 0.56,139.23
X$71 207 206 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $73 r0 *1 0.56,163.8
X$73 243 242 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $75 m0 *1 0.56,163.8
X$75 240 241 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $77 m0 *1 0.56,141.96
X$77 208 209 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $79 m0 *1 0.56,171.99
X$79 252 253 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $81 r0 *1 0.56,171.99
X$81 255 254 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $83 r0 *1 0.56,158.34
X$83 235 234 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $85 m0 *1 0.56,174.72
X$85 256 257 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $87 m0 *1 0.56,169.26
X$87 248 249 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $89 r0 *1 0.56,136.5
X$89 203 202 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $91 r0 *1 0.56,166.53
X$91 247 246 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $93 r0 *1 0.56,174.72
X$93 259 258 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $95 r0 *1 0.56,169.26
X$95 251 250 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $97 r0 *1 0.56,147.42
X$97 219 218 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $99 m0 *1 0.56,158.34
X$99 232 233 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $101 r0 *1 0.56,155.61
X$101 231 230 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $103 m0 *1 0.56,155.61
X$103 228 229 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $105 r0 *1 0.56,161.07
X$105 239 238 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $107 r0 *1 0.56,141.96
X$107 211 210 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $109 m0 *1 0.56,147.42
X$109 216 217 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $111 m0 *1 0.56,150.15
X$111 220 221 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $113 r0 *1 0.56,150.15
X$113 223 222 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $115 m0 *1 0.56,152.88
X$115 224 225 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $117 r0 *1 0.56,152.88
X$117 227 226 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $119 m0 *1 0.56,133.77
X$119 196 197 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $121 r0 *1 0.56,133.77
X$121 199 198 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $123 m0 *1 0.56,136.5
X$123 200 201 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $125 m0 *1 0.56,161.07
X$125 236 237 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $127 m0 *1 0.56,144.69
X$127 212 213 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $129 r0 *1 0.56,144.69
X$129 215 214 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $180 m0 *1 0.56,117.39
X$180 172 173 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $182 r0 *1 0.56,114.66
X$182 171 170 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $184 m0 *1 0.56,114.66
X$184 168 169 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $186 m0 *1 0.56,111.93
X$186 164 165 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $188 r0 *1 0.56,111.93
X$188 167 166 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $190 m0 *1 0.56,109.2
X$190 160 161 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $192 r0 *1 0.56,106.47
X$192 159 158 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $194 m0 *1 0.56,106.47
X$194 156 157 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $196 r0 *1 0.56,103.74
X$196 155 154 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $198 m0 *1 0.56,103.74
X$198 152 153 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $200 r0 *1 0.56,101.01
X$200 151 150 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $202 m0 *1 0.56,101.01
X$202 148 149 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $204 r0 *1 0.56,98.28
X$204 147 146 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $206 r0 *1 0.56,95.55
X$206 143 142 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $208 m0 *1 0.56,95.55
X$208 140 141 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $210 r0 *1 0.56,92.82
X$210 139 138 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $212 m0 *1 0.56,92.82
X$212 136 137 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $214 r0 *1 0.56,90.09
X$214 135 134 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $216 m0 *1 0.56,98.28
X$216 144 145 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $218 r0 *1 0.56,117.39
X$218 175 174 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $220 m0 *1 0.56,120.12
X$220 176 177 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $222 m0 *1 0.56,131.04
X$222 192 193 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $224 r0 *1 0.56,128.31
X$224 191 190 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $226 m0 *1 0.56,128.31
X$226 188 189 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $228 r0 *1 0.56,125.58
X$228 187 186 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $230 m0 *1 0.56,125.58
X$230 184 185 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $232 r0 *1 0.56,122.85
X$232 183 182 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $234 m0 *1 0.56,122.85
X$234 180 181 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $236 r0 *1 0.56,120.12
X$236 179 178 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $238 r0 *1 0.56,131.04
X$238 195 194 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $240 r0 *1 0.56,109.2
X$240 163 162 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* cell instance $258 m0 *1 0.56,90.09
X$258 132 133 131 260 261 freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_decoder
* pin decode_1
* pin decode_0
* pin decode_2
* pin addr_0
* pin addr_1
* pin decode_5
* pin decode_3
* pin decode_4
* pin decode_7
* pin decode_6
* pin addr_3
* pin addr_2
* pin decode_8
* pin decode_10
* pin decode_9
* pin addr_4
* pin addr_5
* pin addr_6
* pin addr_7
* pin decode_11
* pin decode_12
* pin decode_13
* pin decode_14
* pin decode_15
* pin decode_17
* pin decode_16
* pin decode_19
* pin decode_18
* pin decode_20
* pin decode_22
* pin decode_21
* pin decode_25
* pin decode_26
* pin decode_23
* pin decode_24
* pin decode_28
* pin decode_29
* pin decode_27
* pin decode_31
* pin decode_32
* pin decode_30
* pin decode_34
* pin decode_35
* pin decode_33
* pin decode_37
* pin decode_38
* pin decode_36
* pin decode_40
* pin decode_41
* pin decode_39
* pin decode_43
* pin decode_42
* pin decode_44
* pin decode_46
* pin decode_47
* pin decode_45
* pin decode_49
* pin decode_48
* pin decode_50
* pin decode_52
* pin decode_53
* pin decode_51
* pin decode_55
* pin decode_56
* pin decode_54
* pin decode_58
* pin decode_59
* pin decode_57
* pin decode_61
* pin decode_60
* pin decode_62
* pin decode_64
* pin decode_63
* pin decode_65
* pin decode_66
* pin decode_67
* pin decode_68
* pin decode_70
* pin decode_71
* pin decode_69
* pin decode_72
* pin decode_73
* pin decode_74
* pin decode_76
* pin decode_75
* pin decode_77
* pin decode_79
* pin decode_78
* pin decode_80
* pin decode_82
* pin decode_83
* pin decode_81
* pin decode_84
* pin decode_85
* pin decode_86
* pin decode_88
* pin decode_87
* pin decode_89
* pin decode_91
* pin decode_90
* pin decode_92
* pin decode_94
* pin decode_93
* pin decode_95
* pin decode_97
* pin decode_96
* pin decode_98
* pin decode_101
* pin decode_100
* pin decode_99
* pin decode_103
* pin decode_104
* pin decode_102
* pin decode_106
* pin decode_107
* pin decode_105
* pin decode_109
* pin decode_108
* pin decode_110
* pin decode_112
* pin decode_113
* pin decode_111
* pin decode_115
* pin decode_114
* pin decode_116
* pin decode_117
* pin decode_119
* pin decode_118
* pin decode_121
* pin decode_122
* pin decode_120
* pin decode_124
* pin decode_125
* pin decode_123
* pin decode_127
* pin decode_126
* pin decode_128
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_decoder 6 7 8 9 10 13
+ 14 15 17 18 19 20 23 24 25 26 27 28 29 32 33 35 36 37 40 41 44 45 46 50 51 52
+ 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78
+ 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159
* net 6 decode_1
* net 7 decode_0
* net 8 decode_2
* net 9 addr_0
* net 10 addr_1
* net 13 decode_5
* net 14 decode_3
* net 15 decode_4
* net 17 decode_7
* net 18 decode_6
* net 19 addr_3
* net 20 addr_2
* net 23 decode_8
* net 24 decode_10
* net 25 decode_9
* net 26 addr_4
* net 27 addr_5
* net 28 addr_6
* net 29 addr_7
* net 32 decode_11
* net 33 decode_12
* net 35 decode_13
* net 36 decode_14
* net 37 decode_15
* net 40 decode_17
* net 41 decode_16
* net 44 decode_19
* net 45 decode_18
* net 46 decode_20
* net 50 decode_22
* net 51 decode_21
* net 52 decode_25
* net 53 decode_26
* net 54 decode_23
* net 55 decode_24
* net 56 decode_28
* net 57 decode_29
* net 58 decode_27
* net 59 decode_31
* net 60 decode_32
* net 61 decode_30
* net 62 decode_34
* net 63 decode_35
* net 64 decode_33
* net 65 decode_37
* net 66 decode_38
* net 67 decode_36
* net 68 decode_40
* net 69 decode_41
* net 70 decode_39
* net 71 decode_43
* net 72 decode_42
* net 73 decode_44
* net 74 decode_46
* net 75 decode_47
* net 76 decode_45
* net 77 decode_49
* net 78 decode_48
* net 79 decode_50
* net 80 decode_52
* net 81 decode_53
* net 82 decode_51
* net 83 decode_55
* net 84 decode_56
* net 85 decode_54
* net 86 decode_58
* net 87 decode_59
* net 88 decode_57
* net 89 decode_61
* net 90 decode_60
* net 91 decode_62
* net 92 decode_64
* net 93 decode_63
* net 94 decode_65
* net 95 decode_66
* net 96 decode_67
* net 97 decode_68
* net 98 decode_70
* net 99 decode_71
* net 100 decode_69
* net 101 decode_72
* net 102 decode_73
* net 103 decode_74
* net 104 decode_76
* net 105 decode_75
* net 106 decode_77
* net 107 decode_79
* net 108 decode_78
* net 109 decode_80
* net 110 decode_82
* net 111 decode_83
* net 112 decode_81
* net 113 decode_84
* net 114 decode_85
* net 115 decode_86
* net 116 decode_88
* net 117 decode_87
* net 118 decode_89
* net 119 decode_91
* net 120 decode_90
* net 121 decode_92
* net 122 decode_94
* net 123 decode_93
* net 124 decode_95
* net 125 decode_97
* net 126 decode_96
* net 127 decode_98
* net 128 decode_101
* net 129 decode_100
* net 130 decode_99
* net 131 decode_103
* net 132 decode_104
* net 133 decode_102
* net 134 decode_106
* net 135 decode_107
* net 136 decode_105
* net 137 decode_109
* net 138 decode_108
* net 139 decode_110
* net 140 decode_112
* net 141 decode_113
* net 142 decode_111
* net 143 decode_115
* net 144 decode_114
* net 145 decode_116
* net 146 decode_117
* net 147 decode_119
* net 148 decode_118
* net 149 decode_121
* net 150 decode_122
* net 151 decode_120
* net 152 decode_124
* net 153 decode_125
* net 154 decode_123
* net 155 decode_127
* net 156 decode_126
* net 157 decode_128
* net 158 vdd
* net 159 gnd
* cell instance $2 r0 *1 8.745,38.22
X$2 56 1 34 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $3 r0 *1 8.745,131.04
X$3 126 1 4 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $4 r0 *1 8.745,70.98
X$4 80 1 31 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $5 r0 *1 8.745,0
X$5 7 1 4 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $6 r0 *1 8.745,49.14
X$6 67 1 12 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $7 r0 *1 8.745,103.74
X$7 104 1 21 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $8 r0 *1 8.745,32.76
X$8 55 1 30 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $9 r0 *1 8.745,98.28
X$9 101 1 16 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $10 r0 *1 8.745,169.26
X$10 152 1 34 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $11 r0 *1 8.745,21.84
X$11 41 1 22 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $12 r0 *1 8.745,163.8
X$12 151 1 30 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $13 r0 *1 8.745,152.88
X$13 140 1 22 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $14 r0 *1 8.745,16.38
X$14 33 1 21 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $15 r0 *1 8.745,120.12
X$15 116 1 30 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $16 r0 *1 8.745,27.3
X$16 46 1 31 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $17 r0 *1 8.745,109.2
X$17 109 1 22 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $18 r0 *1 8.745,87.36
X$18 92 1 4 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $19 r0 *1 8.745,43.68
X$19 60 1 4 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $20 r0 *1 8.745,60.06
X$20 73 1 21 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $21 r0 *1 8.745,65.52
X$21 78 1 22 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $22 r0 *1 8.745,76.44
X$22 84 1 30 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $23 r0 *1 8.745,141.96
X$23 132 1 16 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $24 r0 *1 8.745,136.5
X$24 129 1 12 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $25 r0 *1 8.745,10.92
X$25 23 1 16 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $26 r0 *1 8.745,54.6
X$26 68 1 16 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $27 r0 *1 8.745,147.42
X$27 138 1 21 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $28 r0 *1 8.745,158.34
X$28 145 1 31 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $29 r0 *1 8.745,174.72
X$29 157 1 4 43 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $30 r0 *1 8.745,125.58
X$30 121 1 34 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $31 r0 *1 8.745,5.46
X$31 15 1 12 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $32 r0 *1 8.745,92.82
X$32 97 1 12 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $33 r0 *1 8.745,81.9
X$33 90 1 34 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $34 r0 *1 8.745,114.66
X$34 113 1 31 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $36 r0 *1 1.9875,0
X$36 9 10 1 2 3 11 158 159
+ freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode2x4
* cell instance $72 m0 *1 8.745,144.69
X$72 136 2 16 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $73 m0 *1 8.745,171.99
X$73 153 2 34 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $74 m0 *1 8.745,35.49
X$74 52 2 30 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $75 m0 *1 8.745,128.31
X$75 123 2 34 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $76 m0 *1 8.745,8.19
X$76 13 2 12 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $77 m0 *1 8.745,155.61
X$77 141 2 22 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $78 m0 *1 8.745,84.63
X$78 89 2 34 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $79 m0 *1 8.745,122.85
X$79 118 2 30 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $80 m0 *1 8.745,166.53
X$80 149 2 30 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $81 m0 *1 8.745,161.07
X$81 146 2 31 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $82 m0 *1 8.745,90.09
X$82 94 2 4 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $83 m0 *1 8.745,40.95
X$83 57 2 34 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $84 m0 *1 8.745,79.17
X$84 88 2 30 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $85 m0 *1 8.745,57.33
X$85 69 2 16 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $86 m0 *1 8.745,2.73
X$86 6 2 4 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $87 m0 *1 8.745,46.41
X$87 64 2 4 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $88 m0 *1 8.745,106.47
X$88 106 2 21 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $89 m0 *1 8.745,101.01
X$89 102 2 16 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $90 m0 *1 8.745,51.87
X$90 65 2 12 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $91 m0 *1 8.745,150.15
X$91 137 2 21 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $92 m0 *1 8.745,62.79
X$92 76 2 21 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $93 m0 *1 8.745,117.39
X$93 114 2 31 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $94 m0 *1 8.745,73.71
X$94 81 2 31 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $95 m0 *1 8.745,30.03
X$95 51 2 31 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $96 m0 *1 8.745,68.25
X$96 77 2 22 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $97 m0 *1 8.745,19.11
X$97 35 2 21 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $98 m0 *1 8.745,13.65
X$98 25 2 16 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $99 m0 *1 8.745,139.23
X$99 128 2 12 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $100 m0 *1 8.745,95.55
X$100 100 2 12 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $101 m0 *1 8.745,24.57
X$101 40 2 22 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $102 m0 *1 8.745,133.77
X$102 125 2 4 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $103 m0 *1 8.745,111.93
X$103 112 2 22 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $139 r0 *1 8.745,40.95
X$139 61 3 34 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $140 r0 *1 8.745,2.73
X$140 8 3 4 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $141 r0 *1 8.745,46.41
X$141 62 3 4 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $142 r0 *1 8.745,73.71
X$142 85 3 31 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $143 r0 *1 8.745,106.47
X$143 108 3 21 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $144 r0 *1 8.745,101.01
X$144 103 3 16 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $145 r0 *1 8.745,68.25
X$145 79 3 22 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $146 r0 *1 8.745,166.53
X$146 150 3 30 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $147 r0 *1 8.745,171.99
X$147 156 3 34 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $148 r0 *1 8.745,35.49
X$148 53 3 30 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $149 r0 *1 8.745,51.87
X$149 66 3 12 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $150 r0 *1 8.745,19.11
X$150 36 3 21 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $151 r0 *1 8.745,13.65
X$151 24 3 16 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $152 r0 *1 8.745,30.03
X$152 50 3 31 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $153 r0 *1 8.745,62.79
X$153 74 3 21 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $154 r0 *1 8.745,155.61
X$154 144 3 22 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $155 r0 *1 8.745,133.77
X$155 127 3 4 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $156 r0 *1 8.745,24.57
X$156 45 3 22 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $157 r0 *1 8.745,139.23
X$157 133 3 12 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $158 r0 *1 8.745,144.69
X$158 134 3 16 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $159 r0 *1 8.745,57.33
X$159 72 3 16 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $160 r0 *1 8.745,95.55
X$160 98 3 12 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $161 r0 *1 8.745,90.09
X$161 95 3 4 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $162 r0 *1 8.745,128.31
X$162 122 3 34 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $163 r0 *1 8.745,8.19
X$163 18 3 12 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $164 r0 *1 8.745,122.85
X$164 120 3 30 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $165 r0 *1 8.745,117.39
X$165 115 3 31 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $166 r0 *1 8.745,111.93
X$166 110 3 22 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $167 r0 *1 8.745,161.07
X$167 148 3 31 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $168 r0 *1 8.745,150.15
X$168 139 3 21 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $169 r0 *1 8.745,79.17
X$169 86 3 30 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $170 r0 *1 8.745,84.63
X$170 91 3 34 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $206 m0 *1 8.745,92.82
X$206 96 11 4 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $207 m0 *1 8.745,5.46
X$207 14 11 4 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $208 m0 *1 8.745,49.14
X$208 63 11 4 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $209 m0 *1 8.745,136.5
X$209 130 11 4 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $211 r0 *1 1.2225,8.19
X$211 20 19 4 12 26 16 21 22 31 30 34 158 159
+ freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8
* cell instance $231 m0 *1 8.745,38.22
X$231 58 11 30 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $232 m0 *1 8.745,10.92
X$232 17 11 12 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $233 m0 *1 8.745,32.76
X$233 54 11 31 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $234 m0 *1 8.745,21.84
X$234 37 11 21 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $235 m0 *1 8.745,16.38
X$235 32 11 16 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $236 m0 *1 8.745,43.68
X$236 59 11 34 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $237 m0 *1 8.745,27.3
X$237 44 11 22 5 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $239 r0 *1 1.2225,21.84
X$239 27 28 5 38 29 39 42 43 47 49 48 158 159
+ freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8
* cell instance $278 m0 *1 8.745,81.9
X$278 87 11 30 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $279 m0 *1 8.745,131.04
X$279 124 11 34 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $280 m0 *1 8.745,174.72
X$280 155 11 34 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $281 m0 *1 8.745,125.58
X$281 119 11 30 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $282 m0 *1 8.745,158.34
X$282 143 11 22 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $283 m0 *1 8.745,163.8
X$283 147 11 31 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $284 m0 *1 8.745,87.36
X$284 93 11 34 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $285 m0 *1 8.745,141.96
X$285 131 11 12 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $286 m0 *1 8.745,60.06
X$286 71 11 16 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $287 m0 *1 8.745,109.2
X$287 107 11 21 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $288 m0 *1 8.745,152.88
X$288 142 11 21 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $289 m0 *1 8.745,65.52
X$289 75 11 21 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $290 m0 *1 8.745,98.28
X$290 99 11 12 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $291 m0 *1 8.745,120.12
X$291 117 11 31 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $292 m0 *1 8.745,76.44
X$292 83 11 31 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $293 m0 *1 8.745,169.26
X$293 154 11 30 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $294 m0 *1 8.745,114.66
X$294 111 11 22 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $295 m0 *1 8.745,54.6
X$295 70 11 12 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $296 m0 *1 8.745,103.74
X$296 105 11 16 39 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $297 m0 *1 8.745,70.98
X$297 82 11 22 38 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $298 m0 *1 8.745,147.42
X$298 135 11 16 42 158 159 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_decoder

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux_array
* pin br_out_31
* pin br_out_30
* pin br_out_29
* pin br_out_28
* pin br_out_27
* pin br_out_26
* pin br_out_25
* pin br_out_24
* pin br_out_23
* pin br_out_22
* pin br_out_21
* pin br_out_20
* pin br_out_19
* pin br_out_18
* pin br_out_0
* pin br_out_17
* pin br_out_16
* pin br_out_15
* pin br_out_14
* pin br_out_13
* pin br_out_12
* pin br_out_11
* pin br_out_10
* pin br_out_9
* pin br_out_8
* pin br_out_7
* pin br_out_6
* pin br_out_5
* pin br_out_4
* pin br_out_3
* pin br_out_2
* pin br_out_1
* pin sel_0
* pin sel_1
* pin sel_2
* pin sel_3
* pin bl_out_31
* pin bl_out_30
* pin bl_out_29
* pin bl_out_0
* pin bl_out_28
* pin bl_out_27
* pin bl_out_26
* pin bl_out_1
* pin bl_out_25
* pin bl_out_24
* pin bl_out_23
* pin bl_out_2
* pin bl_out_22
* pin bl_out_21
* pin bl_out_20
* pin bl_out_19
* pin bl_out_3
* pin bl_out_18
* pin bl_out_17
* pin bl_out_16
* pin bl_out_4
* pin bl_out_15
* pin bl_out_14
* pin bl_out_13
* pin bl_out_5
* pin bl_out_12
* pin bl_out_11
* pin bl_out_10
* pin bl_out_6
* pin bl_out_9
* pin bl_out_8
* pin bl_out_7
* pin sel_4
* pin sel_5
* pin sel_6
* pin sel_7
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin bl_128
* pin br_128
* pin bl_129
* pin br_129
* pin bl_130
* pin br_130
* pin bl_131
* pin br_131
* pin bl_132
* pin br_132
* pin bl_133
* pin br_133
* pin bl_134
* pin br_134
* pin bl_135
* pin br_135
* pin bl_136
* pin br_136
* pin bl_137
* pin br_137
* pin bl_138
* pin br_138
* pin bl_139
* pin br_139
* pin bl_140
* pin br_140
* pin bl_141
* pin br_141
* pin bl_142
* pin br_142
* pin bl_143
* pin br_143
* pin bl_144
* pin br_144
* pin bl_145
* pin br_145
* pin bl_146
* pin br_146
* pin bl_147
* pin br_147
* pin bl_148
* pin br_148
* pin bl_149
* pin br_149
* pin bl_150
* pin br_150
* pin bl_151
* pin br_151
* pin bl_152
* pin br_152
* pin bl_153
* pin br_153
* pin bl_154
* pin br_154
* pin bl_155
* pin br_155
* pin bl_156
* pin br_156
* pin bl_157
* pin br_157
* pin bl_158
* pin br_158
* pin bl_159
* pin br_159
* pin bl_160
* pin br_160
* pin bl_161
* pin br_161
* pin bl_162
* pin br_162
* pin bl_163
* pin br_163
* pin bl_164
* pin br_164
* pin bl_165
* pin br_165
* pin bl_166
* pin br_166
* pin bl_167
* pin br_167
* pin bl_168
* pin br_168
* pin bl_169
* pin br_169
* pin bl_170
* pin br_170
* pin bl_171
* pin br_171
* pin bl_172
* pin br_172
* pin bl_173
* pin br_173
* pin bl_174
* pin br_174
* pin bl_175
* pin br_175
* pin bl_176
* pin br_176
* pin bl_177
* pin br_177
* pin bl_178
* pin br_178
* pin bl_179
* pin br_179
* pin bl_180
* pin br_180
* pin bl_181
* pin br_181
* pin bl_182
* pin br_182
* pin bl_183
* pin br_183
* pin bl_184
* pin br_184
* pin bl_185
* pin br_185
* pin bl_186
* pin br_186
* pin bl_187
* pin br_187
* pin bl_188
* pin br_188
* pin bl_189
* pin br_189
* pin bl_190
* pin br_190
* pin bl_191
* pin br_191
* pin bl_192
* pin br_192
* pin bl_193
* pin br_193
* pin bl_194
* pin br_194
* pin bl_195
* pin br_195
* pin bl_196
* pin br_196
* pin bl_197
* pin br_197
* pin bl_198
* pin br_198
* pin bl_199
* pin br_199
* pin bl_200
* pin br_200
* pin bl_201
* pin br_201
* pin bl_202
* pin br_202
* pin bl_203
* pin br_203
* pin bl_204
* pin br_204
* pin bl_205
* pin br_205
* pin bl_206
* pin br_206
* pin bl_207
* pin br_207
* pin bl_208
* pin br_208
* pin bl_209
* pin br_209
* pin bl_210
* pin br_210
* pin bl_211
* pin br_211
* pin bl_212
* pin br_212
* pin bl_213
* pin br_213
* pin bl_214
* pin br_214
* pin bl_215
* pin br_215
* pin bl_216
* pin br_216
* pin bl_217
* pin br_217
* pin bl_218
* pin br_218
* pin bl_219
* pin br_219
* pin bl_220
* pin br_220
* pin bl_221
* pin br_221
* pin bl_222
* pin br_222
* pin bl_223
* pin br_223
* pin bl_224
* pin br_224
* pin bl_225
* pin br_225
* pin bl_226
* pin br_226
* pin bl_227
* pin br_227
* pin bl_228
* pin br_228
* pin bl_229
* pin br_229
* pin bl_230
* pin br_230
* pin bl_231
* pin br_231
* pin bl_232
* pin br_232
* pin bl_233
* pin br_233
* pin bl_234
* pin br_234
* pin bl_235
* pin br_235
* pin bl_236
* pin br_236
* pin bl_237
* pin br_237
* pin bl_238
* pin br_238
* pin bl_239
* pin br_239
* pin bl_240
* pin br_240
* pin bl_241
* pin br_241
* pin bl_242
* pin br_242
* pin bl_243
* pin br_243
* pin bl_244
* pin br_244
* pin bl_245
* pin br_245
* pin bl_246
* pin br_246
* pin bl_247
* pin br_247
* pin bl_248
* pin br_248
* pin bl_249
* pin br_249
* pin bl_250
* pin br_250
* pin bl_251
* pin br_251
* pin bl_252
* pin br_252
* pin bl_253
* pin br_253
* pin bl_254
* pin br_254
* pin bl_255
* pin br_255
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux_array 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147
+ 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166
+ 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299
+ 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318
+ 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337
+ 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356
+ 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375
+ 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394
+ 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413
+ 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432
+ 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451
+ 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489
+ 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508
+ 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527
+ 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546
+ 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565
+ 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584
+ 585
* net 1 br_out_31
* net 2 br_out_30
* net 3 br_out_29
* net 4 br_out_28
* net 5 br_out_27
* net 6 br_out_26
* net 7 br_out_25
* net 8 br_out_24
* net 9 br_out_23
* net 10 br_out_22
* net 11 br_out_21
* net 12 br_out_20
* net 13 br_out_19
* net 14 br_out_18
* net 15 br_out_0
* net 16 br_out_17
* net 17 br_out_16
* net 18 br_out_15
* net 19 br_out_14
* net 20 br_out_13
* net 21 br_out_12
* net 22 br_out_11
* net 23 br_out_10
* net 24 br_out_9
* net 25 br_out_8
* net 26 br_out_7
* net 27 br_out_6
* net 28 br_out_5
* net 29 br_out_4
* net 30 br_out_3
* net 31 br_out_2
* net 32 br_out_1
* net 33 sel_0
* net 34 sel_1
* net 35 sel_2
* net 36 sel_3
* net 37 bl_out_31
* net 38 bl_out_30
* net 39 bl_out_29
* net 40 bl_out_0
* net 41 bl_out_28
* net 42 bl_out_27
* net 43 bl_out_26
* net 44 bl_out_1
* net 45 bl_out_25
* net 46 bl_out_24
* net 47 bl_out_23
* net 48 bl_out_2
* net 49 bl_out_22
* net 50 bl_out_21
* net 51 bl_out_20
* net 52 bl_out_19
* net 53 bl_out_3
* net 54 bl_out_18
* net 55 bl_out_17
* net 56 bl_out_16
* net 57 bl_out_4
* net 58 bl_out_15
* net 59 bl_out_14
* net 60 bl_out_13
* net 61 bl_out_5
* net 62 bl_out_12
* net 63 bl_out_11
* net 64 bl_out_10
* net 65 bl_out_6
* net 66 bl_out_9
* net 67 bl_out_8
* net 68 bl_out_7
* net 69 sel_4
* net 70 sel_5
* net 71 sel_6
* net 72 sel_7
* net 73 bl_0
* net 74 br_0
* net 75 bl_1
* net 76 br_1
* net 77 bl_2
* net 78 br_2
* net 79 bl_3
* net 80 br_3
* net 81 bl_4
* net 82 br_4
* net 83 bl_5
* net 84 br_5
* net 85 bl_6
* net 86 br_6
* net 87 bl_7
* net 88 br_7
* net 89 bl_8
* net 90 br_8
* net 91 bl_9
* net 92 br_9
* net 93 bl_10
* net 94 br_10
* net 95 bl_11
* net 96 br_11
* net 97 bl_12
* net 98 br_12
* net 99 bl_13
* net 100 br_13
* net 101 bl_14
* net 102 br_14
* net 103 bl_15
* net 104 br_15
* net 105 bl_16
* net 106 br_16
* net 107 bl_17
* net 108 br_17
* net 109 bl_18
* net 110 br_18
* net 111 bl_19
* net 112 br_19
* net 113 bl_20
* net 114 br_20
* net 115 bl_21
* net 116 br_21
* net 117 bl_22
* net 118 br_22
* net 119 bl_23
* net 120 br_23
* net 121 bl_24
* net 122 br_24
* net 123 bl_25
* net 124 br_25
* net 125 bl_26
* net 126 br_26
* net 127 bl_27
* net 128 br_27
* net 129 bl_28
* net 130 br_28
* net 131 bl_29
* net 132 br_29
* net 133 bl_30
* net 134 br_30
* net 135 bl_31
* net 136 br_31
* net 137 bl_32
* net 138 br_32
* net 139 bl_33
* net 140 br_33
* net 141 bl_34
* net 142 br_34
* net 143 bl_35
* net 144 br_35
* net 145 bl_36
* net 146 br_36
* net 147 bl_37
* net 148 br_37
* net 149 bl_38
* net 150 br_38
* net 151 bl_39
* net 152 br_39
* net 153 bl_40
* net 154 br_40
* net 155 bl_41
* net 156 br_41
* net 157 bl_42
* net 158 br_42
* net 159 bl_43
* net 160 br_43
* net 161 bl_44
* net 162 br_44
* net 163 bl_45
* net 164 br_45
* net 165 bl_46
* net 166 br_46
* net 167 bl_47
* net 168 br_47
* net 169 bl_48
* net 170 br_48
* net 171 bl_49
* net 172 br_49
* net 173 bl_50
* net 174 br_50
* net 175 bl_51
* net 176 br_51
* net 177 bl_52
* net 178 br_52
* net 179 bl_53
* net 180 br_53
* net 181 bl_54
* net 182 br_54
* net 183 bl_55
* net 184 br_55
* net 185 bl_56
* net 186 br_56
* net 187 bl_57
* net 188 br_57
* net 189 bl_58
* net 190 br_58
* net 191 bl_59
* net 192 br_59
* net 193 bl_60
* net 194 br_60
* net 195 bl_61
* net 196 br_61
* net 197 bl_62
* net 198 br_62
* net 199 bl_63
* net 200 br_63
* net 201 bl_64
* net 202 br_64
* net 203 bl_65
* net 204 br_65
* net 205 bl_66
* net 206 br_66
* net 207 bl_67
* net 208 br_67
* net 209 bl_68
* net 210 br_68
* net 211 bl_69
* net 212 br_69
* net 213 bl_70
* net 214 br_70
* net 215 bl_71
* net 216 br_71
* net 217 bl_72
* net 218 br_72
* net 219 bl_73
* net 220 br_73
* net 221 bl_74
* net 222 br_74
* net 223 bl_75
* net 224 br_75
* net 225 bl_76
* net 226 br_76
* net 227 bl_77
* net 228 br_77
* net 229 bl_78
* net 230 br_78
* net 231 bl_79
* net 232 br_79
* net 233 bl_80
* net 234 br_80
* net 235 bl_81
* net 236 br_81
* net 237 bl_82
* net 238 br_82
* net 239 bl_83
* net 240 br_83
* net 241 bl_84
* net 242 br_84
* net 243 bl_85
* net 244 br_85
* net 245 bl_86
* net 246 br_86
* net 247 bl_87
* net 248 br_87
* net 249 bl_88
* net 250 br_88
* net 251 bl_89
* net 252 br_89
* net 253 bl_90
* net 254 br_90
* net 255 bl_91
* net 256 br_91
* net 257 bl_92
* net 258 br_92
* net 259 bl_93
* net 260 br_93
* net 261 bl_94
* net 262 br_94
* net 263 bl_95
* net 264 br_95
* net 265 bl_96
* net 266 br_96
* net 267 bl_97
* net 268 br_97
* net 269 bl_98
* net 270 br_98
* net 271 bl_99
* net 272 br_99
* net 273 bl_100
* net 274 br_100
* net 275 bl_101
* net 276 br_101
* net 277 bl_102
* net 278 br_102
* net 279 bl_103
* net 280 br_103
* net 281 bl_104
* net 282 br_104
* net 283 bl_105
* net 284 br_105
* net 285 bl_106
* net 286 br_106
* net 287 bl_107
* net 288 br_107
* net 289 bl_108
* net 290 br_108
* net 291 bl_109
* net 292 br_109
* net 293 bl_110
* net 294 br_110
* net 295 bl_111
* net 296 br_111
* net 297 bl_112
* net 298 br_112
* net 299 bl_113
* net 300 br_113
* net 301 bl_114
* net 302 br_114
* net 303 bl_115
* net 304 br_115
* net 305 bl_116
* net 306 br_116
* net 307 bl_117
* net 308 br_117
* net 309 bl_118
* net 310 br_118
* net 311 bl_119
* net 312 br_119
* net 313 bl_120
* net 314 br_120
* net 315 bl_121
* net 316 br_121
* net 317 bl_122
* net 318 br_122
* net 319 bl_123
* net 320 br_123
* net 321 bl_124
* net 322 br_124
* net 323 bl_125
* net 324 br_125
* net 325 bl_126
* net 326 br_126
* net 327 bl_127
* net 328 br_127
* net 329 bl_128
* net 330 br_128
* net 331 bl_129
* net 332 br_129
* net 333 bl_130
* net 334 br_130
* net 335 bl_131
* net 336 br_131
* net 337 bl_132
* net 338 br_132
* net 339 bl_133
* net 340 br_133
* net 341 bl_134
* net 342 br_134
* net 343 bl_135
* net 344 br_135
* net 345 bl_136
* net 346 br_136
* net 347 bl_137
* net 348 br_137
* net 349 bl_138
* net 350 br_138
* net 351 bl_139
* net 352 br_139
* net 353 bl_140
* net 354 br_140
* net 355 bl_141
* net 356 br_141
* net 357 bl_142
* net 358 br_142
* net 359 bl_143
* net 360 br_143
* net 361 bl_144
* net 362 br_144
* net 363 bl_145
* net 364 br_145
* net 365 bl_146
* net 366 br_146
* net 367 bl_147
* net 368 br_147
* net 369 bl_148
* net 370 br_148
* net 371 bl_149
* net 372 br_149
* net 373 bl_150
* net 374 br_150
* net 375 bl_151
* net 376 br_151
* net 377 bl_152
* net 378 br_152
* net 379 bl_153
* net 380 br_153
* net 381 bl_154
* net 382 br_154
* net 383 bl_155
* net 384 br_155
* net 385 bl_156
* net 386 br_156
* net 387 bl_157
* net 388 br_157
* net 389 bl_158
* net 390 br_158
* net 391 bl_159
* net 392 br_159
* net 393 bl_160
* net 394 br_160
* net 395 bl_161
* net 396 br_161
* net 397 bl_162
* net 398 br_162
* net 399 bl_163
* net 400 br_163
* net 401 bl_164
* net 402 br_164
* net 403 bl_165
* net 404 br_165
* net 405 bl_166
* net 406 br_166
* net 407 bl_167
* net 408 br_167
* net 409 bl_168
* net 410 br_168
* net 411 bl_169
* net 412 br_169
* net 413 bl_170
* net 414 br_170
* net 415 bl_171
* net 416 br_171
* net 417 bl_172
* net 418 br_172
* net 419 bl_173
* net 420 br_173
* net 421 bl_174
* net 422 br_174
* net 423 bl_175
* net 424 br_175
* net 425 bl_176
* net 426 br_176
* net 427 bl_177
* net 428 br_177
* net 429 bl_178
* net 430 br_178
* net 431 bl_179
* net 432 br_179
* net 433 bl_180
* net 434 br_180
* net 435 bl_181
* net 436 br_181
* net 437 bl_182
* net 438 br_182
* net 439 bl_183
* net 440 br_183
* net 441 bl_184
* net 442 br_184
* net 443 bl_185
* net 444 br_185
* net 445 bl_186
* net 446 br_186
* net 447 bl_187
* net 448 br_187
* net 449 bl_188
* net 450 br_188
* net 451 bl_189
* net 452 br_189
* net 453 bl_190
* net 454 br_190
* net 455 bl_191
* net 456 br_191
* net 457 bl_192
* net 458 br_192
* net 459 bl_193
* net 460 br_193
* net 461 bl_194
* net 462 br_194
* net 463 bl_195
* net 464 br_195
* net 465 bl_196
* net 466 br_196
* net 467 bl_197
* net 468 br_197
* net 469 bl_198
* net 470 br_198
* net 471 bl_199
* net 472 br_199
* net 473 bl_200
* net 474 br_200
* net 475 bl_201
* net 476 br_201
* net 477 bl_202
* net 478 br_202
* net 479 bl_203
* net 480 br_203
* net 481 bl_204
* net 482 br_204
* net 483 bl_205
* net 484 br_205
* net 485 bl_206
* net 486 br_206
* net 487 bl_207
* net 488 br_207
* net 489 bl_208
* net 490 br_208
* net 491 bl_209
* net 492 br_209
* net 493 bl_210
* net 494 br_210
* net 495 bl_211
* net 496 br_211
* net 497 bl_212
* net 498 br_212
* net 499 bl_213
* net 500 br_213
* net 501 bl_214
* net 502 br_214
* net 503 bl_215
* net 504 br_215
* net 505 bl_216
* net 506 br_216
* net 507 bl_217
* net 508 br_217
* net 509 bl_218
* net 510 br_218
* net 511 bl_219
* net 512 br_219
* net 513 bl_220
* net 514 br_220
* net 515 bl_221
* net 516 br_221
* net 517 bl_222
* net 518 br_222
* net 519 bl_223
* net 520 br_223
* net 521 bl_224
* net 522 br_224
* net 523 bl_225
* net 524 br_225
* net 525 bl_226
* net 526 br_226
* net 527 bl_227
* net 528 br_227
* net 529 bl_228
* net 530 br_228
* net 531 bl_229
* net 532 br_229
* net 533 bl_230
* net 534 br_230
* net 535 bl_231
* net 536 br_231
* net 537 bl_232
* net 538 br_232
* net 539 bl_233
* net 540 br_233
* net 541 bl_234
* net 542 br_234
* net 543 bl_235
* net 544 br_235
* net 545 bl_236
* net 546 br_236
* net 547 bl_237
* net 548 br_237
* net 549 bl_238
* net 550 br_238
* net 551 bl_239
* net 552 br_239
* net 553 bl_240
* net 554 br_240
* net 555 bl_241
* net 556 br_241
* net 557 bl_242
* net 558 br_242
* net 559 bl_243
* net 560 br_243
* net 561 bl_244
* net 562 br_244
* net 563 bl_245
* net 564 br_245
* net 565 bl_246
* net 566 br_246
* net 567 bl_247
* net 568 br_247
* net 569 bl_248
* net 570 br_248
* net 571 bl_249
* net 572 br_249
* net 573 bl_250
* net 574 br_250
* net 575 bl_251
* net 576 br_251
* net 577 bl_252
* net 578 br_252
* net 579 bl_253
* net 580 br_253
* net 581 bl_254
* net 582 br_254
* net 583 bl_255
* net 584 br_255
* net 585 gnd
* cell instance $1 r0 *1 177.185,1.43
X$1 33 569 1 37 570 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $2 r0 *1 177.89,1.43
X$2 34 571 1 37 572 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $3 r0 *1 178.595,1.43
X$3 35 573 1 37 574 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $4 r0 *1 179.3,1.43
X$4 36 575 1 37 576 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $5 r0 *1 180.005,1.43
X$5 69 577 1 37 578 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $6 r0 *1 180.71,1.43
X$6 70 579 1 37 580 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $7 r0 *1 181.415,1.43
X$7 71 581 1 37 582 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $8 r0 *1 182.12,1.43
X$8 72 583 1 37 584 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $17 r0 *1 176.48,1.43
X$17 72 567 2 38 568 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $18 r0 *1 172.25,1.43
X$18 34 555 2 38 556 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $19 r0 *1 171.545,1.43
X$19 33 553 2 38 554 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $20 r0 *1 173.66,1.43
X$20 36 559 2 38 560 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $21 r0 *1 174.365,1.43
X$21 69 561 2 38 562 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $22 r0 *1 175.775,1.43
X$22 71 565 2 38 566 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $23 r0 *1 175.07,1.43
X$23 70 563 2 38 564 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $24 r0 *1 172.955,1.43
X$24 35 557 2 38 558 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $33 r0 *1 170.84,1.43
X$33 72 551 3 39 552 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $34 r0 *1 165.905,1.43
X$34 33 537 3 39 538 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $35 r0 *1 166.61,1.43
X$35 34 539 3 39 540 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $36 r0 *1 167.315,1.43
X$36 35 541 3 39 542 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $37 r0 *1 168.02,1.43
X$37 36 543 3 39 544 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $38 r0 *1 168.725,1.43
X$38 69 545 3 39 546 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $39 r0 *1 169.43,1.43
X$39 70 547 3 39 548 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $40 r0 *1 170.135,1.43
X$40 71 549 3 39 550 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $49 r0 *1 160.97,1.43
X$49 34 523 4 41 524 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $50 r0 *1 161.675,1.43
X$50 35 525 4 41 526 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $51 r0 *1 162.38,1.43
X$51 36 527 4 41 528 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $52 r0 *1 163.085,1.43
X$52 69 529 4 41 530 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $53 r0 *1 163.79,1.43
X$53 70 531 4 41 532 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $54 r0 *1 160.265,1.43
X$54 33 521 4 41 522 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $55 r0 *1 164.495,1.43
X$55 71 533 4 41 534 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $56 r0 *1 165.2,1.43
X$56 72 535 4 41 536 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $65 r0 *1 159.56,1.43
X$65 72 519 5 42 520 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $66 r0 *1 158.855,1.43
X$66 71 517 5 42 518 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $67 r0 *1 154.625,1.43
X$67 33 505 5 42 506 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $68 r0 *1 155.33,1.43
X$68 34 507 5 42 508 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $69 r0 *1 156.035,1.43
X$69 35 509 5 42 510 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $70 r0 *1 156.74,1.43
X$70 36 511 5 42 512 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $71 r0 *1 157.445,1.43
X$71 69 513 5 42 514 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $72 r0 *1 158.15,1.43
X$72 70 515 5 42 516 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $81 r0 *1 148.985,1.43
X$81 33 489 6 43 490 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $82 r0 *1 149.69,1.43
X$82 34 491 6 43 492 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $83 r0 *1 150.395,1.43
X$83 35 493 6 43 494 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $84 r0 *1 151.1,1.43
X$84 36 495 6 43 496 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $85 r0 *1 151.805,1.43
X$85 69 497 6 43 498 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $86 r0 *1 152.51,1.43
X$86 70 499 6 43 500 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $87 r0 *1 153.215,1.43
X$87 71 501 6 43 502 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $88 r0 *1 153.92,1.43
X$88 72 503 6 43 504 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $97 r0 *1 143.345,1.43
X$97 33 473 7 45 474 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $98 r0 *1 144.05,1.43
X$98 34 475 7 45 476 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $99 r0 *1 144.755,1.43
X$99 35 477 7 45 478 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $100 r0 *1 145.46,1.43
X$100 36 479 7 45 480 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $101 r0 *1 146.165,1.43
X$101 69 481 7 45 482 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $102 r0 *1 146.87,1.43
X$102 70 483 7 45 484 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $103 r0 *1 147.575,1.43
X$103 71 485 7 45 486 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $104 r0 *1 148.28,1.43
X$104 72 487 7 45 488 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $113 r0 *1 137.705,1.43
X$113 33 457 8 46 458 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $114 r0 *1 140.525,1.43
X$114 69 465 8 46 466 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $115 r0 *1 141.23,1.43
X$115 70 467 8 46 468 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $116 r0 *1 141.935,1.43
X$116 71 469 8 46 470 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $117 r0 *1 142.64,1.43
X$117 72 471 8 46 472 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $118 r0 *1 138.41,1.43
X$118 34 459 8 46 460 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $119 r0 *1 139.82,1.43
X$119 36 463 8 46 464 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $120 r0 *1 139.115,1.43
X$120 35 461 8 46 462 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $129 r0 *1 132.77,1.43
X$129 34 443 9 47 444 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $130 r0 *1 133.475,1.43
X$130 35 445 9 47 446 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $131 r0 *1 134.18,1.43
X$131 36 447 9 47 448 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $132 r0 *1 134.885,1.43
X$132 69 449 9 47 450 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $133 r0 *1 135.59,1.43
X$133 70 451 9 47 452 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $134 r0 *1 136.295,1.43
X$134 71 453 9 47 454 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $135 r0 *1 132.065,1.43
X$135 33 441 9 47 442 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $136 r0 *1 137,1.43
X$136 72 455 9 47 456 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $145 r0 *1 126.425,1.43
X$145 33 425 10 49 426 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $146 r0 *1 127.835,1.43
X$146 35 429 10 49 430 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $147 r0 *1 128.54,1.43
X$147 36 431 10 49 432 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $148 r0 *1 129.95,1.43
X$148 70 435 10 49 436 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $149 r0 *1 130.655,1.43
X$149 71 437 10 49 438 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $150 r0 *1 131.36,1.43
X$150 72 439 10 49 440 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $151 r0 *1 127.13,1.43
X$151 34 427 10 49 428 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $152 r0 *1 129.245,1.43
X$152 69 433 10 49 434 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $161 r0 *1 125.72,1.43
X$161 72 423 11 50 424 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $162 r0 *1 120.785,1.43
X$162 33 409 11 50 410 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $163 r0 *1 121.49,1.43
X$163 34 411 11 50 412 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $164 r0 *1 123.605,1.43
X$164 69 417 11 50 418 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $165 r0 *1 122.9,1.43
X$165 36 415 11 50 416 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $166 r0 *1 122.195,1.43
X$166 35 413 11 50 414 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $167 r0 *1 125.015,1.43
X$167 71 421 11 50 422 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $168 r0 *1 124.31,1.43
X$168 70 419 11 50 420 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $177 r0 *1 118.67,1.43
X$177 70 403 12 51 404 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $178 r0 *1 119.375,1.43
X$178 71 405 12 51 406 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $179 r0 *1 115.145,1.43
X$179 33 393 12 51 394 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $180 r0 *1 120.08,1.43
X$180 72 407 12 51 408 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $181 r0 *1 117.965,1.43
X$181 69 401 12 51 402 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $182 r0 *1 117.26,1.43
X$182 36 399 12 51 400 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $183 r0 *1 116.555,1.43
X$183 35 397 12 51 398 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $184 r0 *1 115.85,1.43
X$184 34 395 12 51 396 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $193 r0 *1 114.44,1.43
X$193 72 391 13 52 392 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $194 r0 *1 110.21,1.43
X$194 34 379 13 52 380 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $195 r0 *1 109.505,1.43
X$195 33 377 13 52 378 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $196 r0 *1 110.915,1.43
X$196 35 381 13 52 382 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $197 r0 *1 112.325,1.43
X$197 69 385 13 52 386 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $198 r0 *1 113.03,1.43
X$198 70 387 13 52 388 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $199 r0 *1 113.735,1.43
X$199 71 389 13 52 390 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $200 r0 *1 111.62,1.43
X$200 36 383 13 52 384 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $209 r0 *1 103.865,1.43
X$209 33 361 14 54 362 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $210 r0 *1 108.8,1.43
X$210 72 375 14 54 376 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $211 r0 *1 104.57,1.43
X$211 34 363 14 54 364 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $212 r0 *1 105.275,1.43
X$212 35 365 14 54 366 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $213 r0 *1 105.98,1.43
X$213 36 367 14 54 368 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $214 r0 *1 106.685,1.43
X$214 69 369 14 54 370 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $215 r0 *1 107.39,1.43
X$215 70 371 14 54 372 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $216 r0 *1 108.095,1.43
X$216 71 373 14 54 374 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $225 r0 *1 2.345,1.43
X$225 33 73 15 40 74 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $226 r0 *1 3.05,1.43
X$226 34 75 15 40 76 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $227 r0 *1 5.87,1.43
X$227 70 83 15 40 84 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $228 r0 *1 5.165,1.43
X$228 69 81 15 40 82 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $229 r0 *1 4.46,1.43
X$229 36 79 15 40 80 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $230 r0 *1 3.755,1.43
X$230 35 77 15 40 78 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $231 r0 *1 7.28,1.43
X$231 72 87 15 40 88 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $232 r0 *1 6.575,1.43
X$232 71 85 15 40 86 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $241 r0 *1 103.16,1.43
X$241 72 359 16 55 360 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $242 r0 *1 98.225,1.43
X$242 33 345 16 55 346 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $243 r0 *1 98.93,1.43
X$243 34 347 16 55 348 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $244 r0 *1 99.635,1.43
X$244 35 349 16 55 350 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $245 r0 *1 100.34,1.43
X$245 36 351 16 55 352 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $246 r0 *1 102.455,1.43
X$246 71 357 16 55 358 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $247 r0 *1 101.75,1.43
X$247 70 355 16 55 356 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $248 r0 *1 101.045,1.43
X$248 69 353 16 55 354 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $257 r0 *1 92.585,1.43
X$257 33 329 17 56 330 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $258 r0 *1 97.52,1.43
X$258 72 343 17 56 344 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $259 r0 *1 93.995,1.43
X$259 35 333 17 56 334 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $260 r0 *1 93.29,1.43
X$260 34 331 17 56 332 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $261 r0 *1 96.815,1.43
X$261 71 341 17 56 342 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $262 r0 *1 96.11,1.43
X$262 70 339 17 56 340 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $263 r0 *1 95.405,1.43
X$263 69 337 17 56 338 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $264 r0 *1 94.7,1.43
X$264 36 335 17 56 336 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $273 r0 *1 91.88,1.43
X$273 72 327 18 58 328 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $274 r0 *1 86.945,1.43
X$274 33 313 18 58 314 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $275 r0 *1 87.65,1.43
X$275 34 315 18 58 316 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $276 r0 *1 88.355,1.43
X$276 35 317 18 58 318 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $277 r0 *1 89.06,1.43
X$277 36 319 18 58 320 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $278 r0 *1 89.765,1.43
X$278 69 321 18 58 322 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $279 r0 *1 90.47,1.43
X$279 70 323 18 58 324 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $280 r0 *1 91.175,1.43
X$280 71 325 18 58 326 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $289 r0 *1 81.305,1.43
X$289 33 297 19 59 298 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $290 r0 *1 82.715,1.43
X$290 35 301 19 59 302 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $291 r0 *1 83.42,1.43
X$291 36 303 19 59 304 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $292 r0 *1 84.125,1.43
X$292 69 305 19 59 306 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $293 r0 *1 84.83,1.43
X$293 70 307 19 59 308 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $294 r0 *1 85.535,1.43
X$294 71 309 19 59 310 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $295 r0 *1 86.24,1.43
X$295 72 311 19 59 312 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $296 r0 *1 82.01,1.43
X$296 34 299 19 59 300 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $305 r0 *1 80.6,1.43
X$305 72 295 20 60 296 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $306 r0 *1 79.895,1.43
X$306 71 293 20 60 294 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $307 r0 *1 79.19,1.43
X$307 70 291 20 60 292 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $308 r0 *1 78.485,1.43
X$308 69 289 20 60 290 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $309 r0 *1 77.78,1.43
X$309 36 287 20 60 288 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $310 r0 *1 77.075,1.43
X$310 35 285 20 60 286 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $311 r0 *1 76.37,1.43
X$311 34 283 20 60 284 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $312 r0 *1 75.665,1.43
X$312 33 281 20 60 282 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $321 r0 *1 70.025,1.43
X$321 33 265 21 62 266 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $322 r0 *1 71.435,1.43
X$322 35 269 21 62 270 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $323 r0 *1 73.55,1.43
X$323 70 275 21 62 276 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $324 r0 *1 74.255,1.43
X$324 71 277 21 62 278 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $325 r0 *1 74.96,1.43
X$325 72 279 21 62 280 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $326 r0 *1 72.845,1.43
X$326 69 273 21 62 274 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $327 r0 *1 72.14,1.43
X$327 36 271 21 62 272 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $328 r0 *1 70.73,1.43
X$328 34 267 21 62 268 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $337 r0 *1 69.32,1.43
X$337 72 263 22 63 264 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $338 r0 *1 65.795,1.43
X$338 35 253 22 63 254 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $339 r0 *1 66.5,1.43
X$339 36 255 22 63 256 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $340 r0 *1 67.205,1.43
X$340 69 257 22 63 258 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $341 r0 *1 67.91,1.43
X$341 70 259 22 63 260 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $342 r0 *1 68.615,1.43
X$342 71 261 22 63 262 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $343 r0 *1 65.09,1.43
X$343 34 251 22 63 252 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $344 r0 *1 64.385,1.43
X$344 33 249 22 63 250 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $353 r0 *1 59.45,1.43
X$353 34 235 23 64 236 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $354 r0 *1 60.155,1.43
X$354 35 237 23 64 238 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $355 r0 *1 58.745,1.43
X$355 33 233 23 64 234 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $356 r0 *1 60.86,1.43
X$356 36 239 23 64 240 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $357 r0 *1 62.975,1.43
X$357 71 245 23 64 246 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $358 r0 *1 63.68,1.43
X$358 72 247 23 64 248 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $359 r0 *1 61.565,1.43
X$359 69 241 23 64 242 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $360 r0 *1 62.27,1.43
X$360 70 243 23 64 244 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $369 r0 *1 53.105,1.43
X$369 33 217 24 66 218 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $370 r0 *1 53.81,1.43
X$370 34 219 24 66 220 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $371 r0 *1 54.515,1.43
X$371 35 221 24 66 222 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $372 r0 *1 58.04,1.43
X$372 72 231 24 66 232 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $373 r0 *1 57.335,1.43
X$373 71 229 24 66 230 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $374 r0 *1 56.63,1.43
X$374 70 227 24 66 228 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $375 r0 *1 55.925,1.43
X$375 69 225 24 66 226 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $376 r0 *1 55.22,1.43
X$376 36 223 24 66 224 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $385 r0 *1 48.875,1.43
X$385 35 205 25 67 206 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $386 r0 *1 48.17,1.43
X$386 34 203 25 67 204 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $387 r0 *1 52.4,1.43
X$387 72 215 25 67 216 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $388 r0 *1 49.58,1.43
X$388 36 207 25 67 208 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $389 r0 *1 50.285,1.43
X$389 69 209 25 67 210 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $390 r0 *1 50.99,1.43
X$390 70 211 25 67 212 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $391 r0 *1 51.695,1.43
X$391 71 213 25 67 214 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $392 r0 *1 47.465,1.43
X$392 33 201 25 67 202 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $401 r0 *1 41.825,1.43
X$401 33 185 26 68 186 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $402 r0 *1 46.055,1.43
X$402 71 197 26 68 198 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $403 r0 *1 45.35,1.43
X$403 70 195 26 68 196 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $404 r0 *1 44.645,1.43
X$404 69 193 26 68 194 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $405 r0 *1 43.94,1.43
X$405 36 191 26 68 192 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $406 r0 *1 43.235,1.43
X$406 35 189 26 68 190 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $407 r0 *1 42.53,1.43
X$407 34 187 26 68 188 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $408 r0 *1 46.76,1.43
X$408 72 199 26 68 200 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $417 r0 *1 36.89,1.43
X$417 34 171 27 65 172 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $418 r0 *1 37.595,1.43
X$418 35 173 27 65 174 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $419 r0 *1 38.3,1.43
X$419 36 175 27 65 176 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $420 r0 *1 39.005,1.43
X$420 69 177 27 65 178 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $421 r0 *1 40.415,1.43
X$421 71 181 27 65 182 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $422 r0 *1 41.12,1.43
X$422 72 183 27 65 184 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $423 r0 *1 39.71,1.43
X$423 70 179 27 65 180 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $424 r0 *1 36.185,1.43
X$424 33 169 27 65 170 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $433 r0 *1 35.48,1.43
X$433 72 167 28 61 168 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $434 r0 *1 34.775,1.43
X$434 71 165 28 61 166 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $435 r0 *1 34.07,1.43
X$435 70 163 28 61 164 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $436 r0 *1 33.365,1.43
X$436 69 161 28 61 162 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $437 r0 *1 32.66,1.43
X$437 36 159 28 61 160 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $438 r0 *1 31.955,1.43
X$438 35 157 28 61 158 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $439 r0 *1 31.25,1.43
X$439 34 155 28 61 156 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $440 r0 *1 30.545,1.43
X$440 33 153 28 61 154 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $449 r0 *1 24.905,1.43
X$449 33 137 29 57 138 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $450 r0 *1 26.315,1.43
X$450 35 141 29 57 142 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $451 r0 *1 25.61,1.43
X$451 34 139 29 57 140 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $452 r0 *1 29.135,1.43
X$452 71 149 29 57 150 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $453 r0 *1 28.43,1.43
X$453 70 147 29 57 148 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $454 r0 *1 27.725,1.43
X$454 69 145 29 57 146 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $455 r0 *1 27.02,1.43
X$455 36 143 29 57 144 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $456 r0 *1 29.84,1.43
X$456 72 151 29 57 152 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $465 r0 *1 24.2,1.43
X$465 72 135 30 53 136 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $466 r0 *1 23.495,1.43
X$466 71 133 30 53 134 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $467 r0 *1 22.79,1.43
X$467 70 131 30 53 132 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $468 r0 *1 22.085,1.43
X$468 69 129 30 53 130 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $469 r0 *1 21.38,1.43
X$469 36 127 30 53 128 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $470 r0 *1 20.675,1.43
X$470 35 125 30 53 126 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $471 r0 *1 19.97,1.43
X$471 34 123 30 53 124 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $472 r0 *1 19.265,1.43
X$472 33 121 30 53 122 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $481 r0 *1 17.15,1.43
X$481 70 115 31 48 116 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $482 r0 *1 16.445,1.43
X$482 69 113 31 48 114 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $483 r0 *1 15.74,1.43
X$483 36 111 31 48 112 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $484 r0 *1 15.035,1.43
X$484 35 109 31 48 110 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $485 r0 *1 14.33,1.43
X$485 34 107 31 48 108 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $486 r0 *1 17.855,1.43
X$486 71 117 31 48 118 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $487 r0 *1 18.56,1.43
X$487 72 119 31 48 120 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $488 r0 *1 13.625,1.43
X$488 33 105 31 48 106 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $497 r0 *1 12.215,1.43
X$497 71 101 32 44 102 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $498 r0 *1 9.395,1.43
X$498 35 93 32 44 94 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $499 r0 *1 8.69,1.43
X$499 34 91 32 44 92 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $500 r0 *1 7.985,1.43
X$500 33 89 32 44 90 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $501 r0 *1 11.51,1.43
X$501 70 99 32 44 100 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $502 r0 *1 10.805,1.43
X$502 69 97 32 44 98 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $503 r0 *1 10.1,1.43
X$503 36 95 32 44 96 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* cell instance $504 r0 *1 12.92,1.43
X$504 72 103 32 44 104 585 freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_write_mask_and_array
* pin wmask_out_0
* pin wmask_out_1
* pin wmask_out_2
* pin wmask_out_3
* pin wmask_in_0
* pin wmask_in_1
* pin wmask_in_2
* pin wmask_in_3
* pin en
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_write_mask_and_array 1 2 3 4 5 6 7
+ 8 9 10 11
* net 1 wmask_out_0
* net 2 wmask_out_1
* net 3 wmask_out_2
* net 4 wmask_out_3
* net 5 wmask_in_0
* net 6 wmask_in_1
* net 7 wmask_in_2
* net 8 wmask_in_3
* net 9 en
* net 10 vdd
* net 11 gnd
* cell instance $1 r0 *1 2.345,0
X$1 1 5 9 10 11 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2
* cell instance $2 r0 *1 47.465,0
X$2 2 6 9 10 11 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2
* cell instance $3 r0 *1 92.585,0
X$3 3 7 9 10 11 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2
* cell instance $4 r0 *1 137.705,0
X$4 4 8 9 10 11 freepdk45_sram_4kbytes_1rw_32x1024_8_pand2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_write_mask_and_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_write_driver_array
* pin data_0
* pin data_1
* pin data_2
* pin data_3
* pin data_4
* pin data_5
* pin data_6
* pin data_7
* pin data_8
* pin data_9
* pin data_10
* pin data_11
* pin data_12
* pin data_13
* pin data_14
* pin data_15
* pin data_16
* pin data_17
* pin data_18
* pin data_19
* pin data_20
* pin data_21
* pin data_22
* pin data_23
* pin data_24
* pin data_25
* pin data_26
* pin data_27
* pin data_28
* pin data_29
* pin data_30
* pin data_31
* pin data_32
* pin br_0
* pin br_1
* pin br_2
* pin br_3
* pin en_0
* pin br_4
* pin br_5
* pin br_6
* pin br_7
* pin br_8
* pin br_9
* pin br_10
* pin br_11
* pin en_1
* pin br_12
* pin br_13
* pin br_14
* pin br_15
* pin br_16
* pin br_17
* pin br_18
* pin br_19
* pin en_2
* pin br_20
* pin br_21
* pin br_22
* pin br_23
* pin br_24
* pin br_25
* pin br_26
* pin br_27
* pin en_3
* pin br_28
* pin br_29
* pin br_30
* pin br_31
* pin br_32
* pin en_4
* pin bl_0
* pin bl_1
* pin bl_2
* pin bl_3
* pin bl_4
* pin bl_5
* pin bl_6
* pin bl_7
* pin bl_8
* pin bl_9
* pin bl_10
* pin bl_11
* pin bl_12
* pin bl_13
* pin bl_14
* pin bl_15
* pin bl_16
* pin bl_17
* pin bl_18
* pin bl_19
* pin bl_20
* pin bl_21
* pin bl_22
* pin bl_23
* pin bl_24
* pin bl_25
* pin bl_26
* pin bl_27
* pin bl_28
* pin bl_29
* pin bl_30
* pin bl_31
* pin bl_32
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_write_driver_array 1 2 3 4 5 6 7 8
+ 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34
+ 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86
+ 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106
* net 1 data_0
* net 2 data_1
* net 3 data_2
* net 4 data_3
* net 5 data_4
* net 6 data_5
* net 7 data_6
* net 8 data_7
* net 9 data_8
* net 10 data_9
* net 11 data_10
* net 12 data_11
* net 13 data_12
* net 14 data_13
* net 15 data_14
* net 16 data_15
* net 17 data_16
* net 18 data_17
* net 19 data_18
* net 20 data_19
* net 21 data_20
* net 22 data_21
* net 23 data_22
* net 24 data_23
* net 25 data_24
* net 26 data_25
* net 27 data_26
* net 28 data_27
* net 29 data_28
* net 30 data_29
* net 31 data_30
* net 32 data_31
* net 33 data_32
* net 34 br_0
* net 35 br_1
* net 36 br_2
* net 37 br_3
* net 38 en_0
* net 39 br_4
* net 40 br_5
* net 41 br_6
* net 42 br_7
* net 43 br_8
* net 44 br_9
* net 45 br_10
* net 46 br_11
* net 47 en_1
* net 48 br_12
* net 49 br_13
* net 50 br_14
* net 51 br_15
* net 52 br_16
* net 53 br_17
* net 54 br_18
* net 55 br_19
* net 56 en_2
* net 57 br_20
* net 58 br_21
* net 59 br_22
* net 60 br_23
* net 61 br_24
* net 62 br_25
* net 63 br_26
* net 64 br_27
* net 65 en_3
* net 66 br_28
* net 67 br_29
* net 68 br_30
* net 69 br_31
* net 70 br_32
* net 71 en_4
* net 72 bl_0
* net 73 bl_1
* net 74 bl_2
* net 75 bl_3
* net 76 bl_4
* net 77 bl_5
* net 78 bl_6
* net 79 bl_7
* net 80 bl_8
* net 81 bl_9
* net 82 bl_10
* net 83 bl_11
* net 84 bl_12
* net 85 bl_13
* net 86 bl_14
* net 87 bl_15
* net 88 bl_16
* net 89 bl_17
* net 90 bl_18
* net 91 bl_19
* net 92 bl_20
* net 93 bl_21
* net 94 bl_22
* net 95 bl_23
* net 96 bl_24
* net 97 bl_25
* net 98 bl_26
* net 99 bl_27
* net 100 bl_28
* net 101 bl_29
* net 102 bl_30
* net 103 bl_31
* net 104 bl_32
* net 105 vdd
* net 106 gnd
* cell instance $1 r0 *1 2.345,0
X$1 1 38 34 72 105 106 write_driver
* cell instance $2 r0 *1 7.985,0
X$2 2 38 35 73 105 106 write_driver
* cell instance $3 r0 *1 13.625,0
X$3 3 38 36 74 105 106 write_driver
* cell instance $4 r0 *1 19.265,0
X$4 4 38 37 75 105 106 write_driver
* cell instance $5 r0 *1 24.905,0
X$5 5 38 39 76 105 106 write_driver
* cell instance $6 r0 *1 30.545,0
X$6 6 38 40 77 105 106 write_driver
* cell instance $7 r0 *1 36.185,0
X$7 7 38 41 78 105 106 write_driver
* cell instance $8 r0 *1 41.825,0
X$8 8 38 42 79 105 106 write_driver
* cell instance $9 r0 *1 47.465,0
X$9 9 47 43 80 105 106 write_driver
* cell instance $10 r0 *1 53.105,0
X$10 10 47 44 81 105 106 write_driver
* cell instance $11 r0 *1 58.745,0
X$11 11 47 45 82 105 106 write_driver
* cell instance $12 r0 *1 64.385,0
X$12 12 47 46 83 105 106 write_driver
* cell instance $13 r0 *1 70.025,0
X$13 13 47 48 84 105 106 write_driver
* cell instance $14 r0 *1 75.665,0
X$14 14 47 49 85 105 106 write_driver
* cell instance $15 r0 *1 81.305,0
X$15 15 47 50 86 105 106 write_driver
* cell instance $16 r0 *1 86.945,0
X$16 16 47 51 87 105 106 write_driver
* cell instance $17 r0 *1 92.585,0
X$17 17 56 52 88 105 106 write_driver
* cell instance $18 r0 *1 98.225,0
X$18 18 56 53 89 105 106 write_driver
* cell instance $19 r0 *1 103.865,0
X$19 19 56 54 90 105 106 write_driver
* cell instance $20 r0 *1 109.505,0
X$20 20 56 55 91 105 106 write_driver
* cell instance $21 r0 *1 115.145,0
X$21 21 56 57 92 105 106 write_driver
* cell instance $22 r0 *1 120.785,0
X$22 22 56 58 93 105 106 write_driver
* cell instance $23 r0 *1 126.425,0
X$23 23 56 59 94 105 106 write_driver
* cell instance $24 r0 *1 132.065,0
X$24 24 56 60 95 105 106 write_driver
* cell instance $25 r0 *1 137.705,0
X$25 25 65 61 96 105 106 write_driver
* cell instance $26 r0 *1 143.345,0
X$26 26 65 62 97 105 106 write_driver
* cell instance $27 r0 *1 148.985,0
X$27 27 65 63 98 105 106 write_driver
* cell instance $28 r0 *1 154.625,0
X$28 28 65 64 99 105 106 write_driver
* cell instance $29 r0 *1 160.265,0
X$29 29 65 66 100 105 106 write_driver
* cell instance $30 r0 *1 165.905,0
X$30 30 65 67 101 105 106 write_driver
* cell instance $31 r0 *1 171.545,0
X$31 31 65 68 102 105 106 write_driver
* cell instance $32 r0 *1 177.185,0
X$32 32 65 69 103 105 106 write_driver
* cell instance $33 r0 *1 182.825,0
X$33 33 71 70 104 105 106 write_driver
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_write_driver_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_sense_amp_array
* pin data_0
* pin bl_0
* pin br_0
* pin data_1
* pin bl_1
* pin br_1
* pin data_2
* pin bl_2
* pin br_2
* pin data_3
* pin bl_3
* pin br_3
* pin data_4
* pin bl_4
* pin br_4
* pin data_5
* pin bl_5
* pin br_5
* pin data_6
* pin bl_6
* pin br_6
* pin data_7
* pin bl_7
* pin br_7
* pin data_8
* pin bl_8
* pin br_8
* pin data_9
* pin bl_9
* pin br_9
* pin data_10
* pin bl_10
* pin br_10
* pin data_11
* pin bl_11
* pin br_11
* pin data_12
* pin bl_12
* pin br_12
* pin data_13
* pin bl_13
* pin br_13
* pin data_14
* pin bl_14
* pin br_14
* pin data_15
* pin bl_15
* pin br_15
* pin data_16
* pin bl_16
* pin br_16
* pin data_17
* pin bl_17
* pin br_17
* pin data_18
* pin bl_18
* pin br_18
* pin data_19
* pin bl_19
* pin br_19
* pin data_20
* pin bl_20
* pin br_20
* pin data_21
* pin bl_21
* pin br_21
* pin data_22
* pin bl_22
* pin br_22
* pin data_23
* pin bl_23
* pin br_23
* pin data_24
* pin bl_24
* pin br_24
* pin data_25
* pin bl_25
* pin br_25
* pin data_26
* pin bl_26
* pin br_26
* pin data_27
* pin bl_27
* pin br_27
* pin data_28
* pin bl_28
* pin br_28
* pin data_29
* pin bl_29
* pin br_29
* pin data_30
* pin bl_30
* pin br_30
* pin data_31
* pin bl_31
* pin br_31
* pin data_32
* pin bl_32
* pin br_32
* pin en
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_sense_amp_array 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
* net 1 data_0
* net 2 bl_0
* net 3 br_0
* net 4 data_1
* net 5 bl_1
* net 6 br_1
* net 7 data_2
* net 8 bl_2
* net 9 br_2
* net 10 data_3
* net 11 bl_3
* net 12 br_3
* net 13 data_4
* net 14 bl_4
* net 15 br_4
* net 16 data_5
* net 17 bl_5
* net 18 br_5
* net 19 data_6
* net 20 bl_6
* net 21 br_6
* net 22 data_7
* net 23 bl_7
* net 24 br_7
* net 25 data_8
* net 26 bl_8
* net 27 br_8
* net 28 data_9
* net 29 bl_9
* net 30 br_9
* net 31 data_10
* net 32 bl_10
* net 33 br_10
* net 34 data_11
* net 35 bl_11
* net 36 br_11
* net 37 data_12
* net 38 bl_12
* net 39 br_12
* net 40 data_13
* net 41 bl_13
* net 42 br_13
* net 43 data_14
* net 44 bl_14
* net 45 br_14
* net 46 data_15
* net 47 bl_15
* net 48 br_15
* net 49 data_16
* net 50 bl_16
* net 51 br_16
* net 52 data_17
* net 53 bl_17
* net 54 br_17
* net 55 data_18
* net 56 bl_18
* net 57 br_18
* net 58 data_19
* net 59 bl_19
* net 60 br_19
* net 61 data_20
* net 62 bl_20
* net 63 br_20
* net 64 data_21
* net 65 bl_21
* net 66 br_21
* net 67 data_22
* net 68 bl_22
* net 69 br_22
* net 70 data_23
* net 71 bl_23
* net 72 br_23
* net 73 data_24
* net 74 bl_24
* net 75 br_24
* net 76 data_25
* net 77 bl_25
* net 78 br_25
* net 79 data_26
* net 80 bl_26
* net 81 br_26
* net 82 data_27
* net 83 bl_27
* net 84 br_27
* net 85 data_28
* net 86 bl_28
* net 87 br_28
* net 88 data_29
* net 89 bl_29
* net 90 br_29
* net 91 data_30
* net 92 bl_30
* net 93 br_30
* net 94 data_31
* net 95 bl_31
* net 96 br_31
* net 97 data_32
* net 98 bl_32
* net 99 br_32
* net 100 en
* net 101 vdd
* net 102 gnd
* cell instance $1 r0 *1 2.345,0
X$1 3 2 1 100 101 102 sense_amp
* cell instance $2 r0 *1 7.985,0
X$2 6 5 4 100 101 102 sense_amp
* cell instance $3 r0 *1 13.625,0
X$3 9 8 7 100 101 102 sense_amp
* cell instance $4 r0 *1 19.265,0
X$4 12 11 10 100 101 102 sense_amp
* cell instance $5 r0 *1 24.905,0
X$5 15 14 13 100 101 102 sense_amp
* cell instance $6 r0 *1 30.545,0
X$6 18 17 16 100 101 102 sense_amp
* cell instance $7 r0 *1 36.185,0
X$7 21 20 19 100 101 102 sense_amp
* cell instance $8 r0 *1 41.825,0
X$8 24 23 22 100 101 102 sense_amp
* cell instance $9 r0 *1 47.465,0
X$9 27 26 25 100 101 102 sense_amp
* cell instance $10 r0 *1 53.105,0
X$10 30 29 28 100 101 102 sense_amp
* cell instance $11 r0 *1 58.745,0
X$11 33 32 31 100 101 102 sense_amp
* cell instance $12 r0 *1 64.385,0
X$12 36 35 34 100 101 102 sense_amp
* cell instance $13 r0 *1 70.025,0
X$13 39 38 37 100 101 102 sense_amp
* cell instance $14 r0 *1 75.665,0
X$14 42 41 40 100 101 102 sense_amp
* cell instance $15 r0 *1 81.305,0
X$15 45 44 43 100 101 102 sense_amp
* cell instance $16 r0 *1 86.945,0
X$16 48 47 46 100 101 102 sense_amp
* cell instance $17 r0 *1 92.585,0
X$17 51 50 49 100 101 102 sense_amp
* cell instance $18 r0 *1 98.225,0
X$18 54 53 52 100 101 102 sense_amp
* cell instance $19 r0 *1 103.865,0
X$19 57 56 55 100 101 102 sense_amp
* cell instance $20 r0 *1 109.505,0
X$20 60 59 58 100 101 102 sense_amp
* cell instance $21 r0 *1 115.145,0
X$21 63 62 61 100 101 102 sense_amp
* cell instance $22 r0 *1 120.785,0
X$22 66 65 64 100 101 102 sense_amp
* cell instance $23 r0 *1 126.425,0
X$23 69 68 67 100 101 102 sense_amp
* cell instance $24 r0 *1 132.065,0
X$24 72 71 70 100 101 102 sense_amp
* cell instance $25 r0 *1 137.705,0
X$25 75 74 73 100 101 102 sense_amp
* cell instance $26 r0 *1 143.345,0
X$26 78 77 76 100 101 102 sense_amp
* cell instance $27 r0 *1 148.985,0
X$27 81 80 79 100 101 102 sense_amp
* cell instance $28 r0 *1 154.625,0
X$28 84 83 82 100 101 102 sense_amp
* cell instance $29 r0 *1 160.265,0
X$29 87 86 85 100 101 102 sense_amp
* cell instance $30 r0 *1 165.905,0
X$30 90 89 88 100 101 102 sense_amp
* cell instance $31 r0 *1 171.545,0
X$31 93 92 91 100 101 102 sense_amp
* cell instance $32 r0 *1 177.185,0
X$32 96 95 94 100 101 102 sense_amp
* cell instance $33 r0 *1 182.825,0
X$33 99 98 97 100 101 102 sense_amp
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_sense_amp_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_array
* pin en_bar
* pin bl_0
* pin br_0
* pin bl_1
* pin br_1
* pin bl_2
* pin br_2
* pin bl_3
* pin br_3
* pin bl_4
* pin br_4
* pin bl_5
* pin br_5
* pin bl_6
* pin br_6
* pin bl_7
* pin br_7
* pin bl_8
* pin br_8
* pin bl_9
* pin br_9
* pin bl_10
* pin br_10
* pin bl_11
* pin br_11
* pin bl_12
* pin br_12
* pin bl_13
* pin br_13
* pin bl_14
* pin br_14
* pin bl_15
* pin br_15
* pin bl_16
* pin br_16
* pin bl_17
* pin br_17
* pin bl_18
* pin br_18
* pin bl_19
* pin br_19
* pin bl_20
* pin br_20
* pin bl_21
* pin br_21
* pin bl_22
* pin br_22
* pin bl_23
* pin br_23
* pin bl_24
* pin br_24
* pin bl_25
* pin br_25
* pin bl_26
* pin br_26
* pin bl_27
* pin br_27
* pin bl_28
* pin br_28
* pin bl_29
* pin br_29
* pin bl_30
* pin br_30
* pin bl_31
* pin br_31
* pin bl_32
* pin br_32
* pin bl_33
* pin br_33
* pin bl_34
* pin br_34
* pin bl_35
* pin br_35
* pin bl_36
* pin br_36
* pin bl_37
* pin br_37
* pin bl_38
* pin br_38
* pin bl_39
* pin br_39
* pin bl_40
* pin br_40
* pin bl_41
* pin br_41
* pin bl_42
* pin br_42
* pin bl_43
* pin br_43
* pin bl_44
* pin br_44
* pin bl_45
* pin br_45
* pin bl_46
* pin br_46
* pin bl_47
* pin br_47
* pin bl_48
* pin br_48
* pin bl_49
* pin br_49
* pin bl_50
* pin br_50
* pin bl_51
* pin br_51
* pin bl_52
* pin br_52
* pin bl_53
* pin br_53
* pin bl_54
* pin br_54
* pin bl_55
* pin br_55
* pin bl_56
* pin br_56
* pin bl_57
* pin br_57
* pin bl_58
* pin br_58
* pin bl_59
* pin br_59
* pin bl_60
* pin br_60
* pin bl_61
* pin br_61
* pin bl_62
* pin br_62
* pin bl_63
* pin br_63
* pin bl_64
* pin br_64
* pin bl_65
* pin br_65
* pin bl_66
* pin br_66
* pin bl_67
* pin br_67
* pin bl_68
* pin br_68
* pin bl_69
* pin br_69
* pin bl_70
* pin br_70
* pin bl_71
* pin br_71
* pin bl_72
* pin br_72
* pin bl_73
* pin br_73
* pin bl_74
* pin br_74
* pin bl_75
* pin br_75
* pin bl_76
* pin br_76
* pin bl_77
* pin br_77
* pin bl_78
* pin br_78
* pin bl_79
* pin br_79
* pin bl_80
* pin br_80
* pin bl_81
* pin br_81
* pin bl_82
* pin br_82
* pin bl_83
* pin br_83
* pin bl_84
* pin br_84
* pin bl_85
* pin br_85
* pin bl_86
* pin br_86
* pin bl_87
* pin br_87
* pin bl_88
* pin br_88
* pin bl_89
* pin br_89
* pin bl_90
* pin br_90
* pin bl_91
* pin br_91
* pin bl_92
* pin br_92
* pin bl_93
* pin br_93
* pin bl_94
* pin br_94
* pin bl_95
* pin br_95
* pin bl_96
* pin br_96
* pin bl_97
* pin br_97
* pin bl_98
* pin br_98
* pin bl_99
* pin br_99
* pin bl_100
* pin br_100
* pin bl_101
* pin br_101
* pin bl_102
* pin br_102
* pin bl_103
* pin br_103
* pin bl_104
* pin br_104
* pin bl_105
* pin br_105
* pin bl_106
* pin br_106
* pin bl_107
* pin br_107
* pin bl_108
* pin br_108
* pin bl_109
* pin br_109
* pin bl_110
* pin br_110
* pin bl_111
* pin br_111
* pin bl_112
* pin br_112
* pin bl_113
* pin br_113
* pin bl_114
* pin br_114
* pin bl_115
* pin br_115
* pin bl_116
* pin br_116
* pin bl_117
* pin br_117
* pin bl_118
* pin br_118
* pin bl_119
* pin br_119
* pin bl_120
* pin br_120
* pin bl_121
* pin br_121
* pin bl_122
* pin br_122
* pin bl_123
* pin br_123
* pin bl_124
* pin br_124
* pin bl_125
* pin br_125
* pin bl_126
* pin br_126
* pin bl_127
* pin br_127
* pin bl_128
* pin br_128
* pin bl_129
* pin br_129
* pin bl_130
* pin br_130
* pin bl_131
* pin br_131
* pin bl_132
* pin br_132
* pin bl_133
* pin br_133
* pin bl_134
* pin br_134
* pin bl_135
* pin br_135
* pin bl_136
* pin br_136
* pin bl_137
* pin br_137
* pin bl_138
* pin br_138
* pin bl_139
* pin br_139
* pin bl_140
* pin br_140
* pin bl_141
* pin br_141
* pin bl_142
* pin br_142
* pin bl_143
* pin br_143
* pin bl_144
* pin br_144
* pin bl_145
* pin br_145
* pin bl_146
* pin br_146
* pin bl_147
* pin br_147
* pin bl_148
* pin br_148
* pin bl_149
* pin br_149
* pin bl_150
* pin br_150
* pin bl_151
* pin br_151
* pin bl_152
* pin br_152
* pin bl_153
* pin br_153
* pin bl_154
* pin br_154
* pin bl_155
* pin br_155
* pin bl_156
* pin br_156
* pin bl_157
* pin br_157
* pin bl_158
* pin br_158
* pin bl_159
* pin br_159
* pin bl_160
* pin br_160
* pin bl_161
* pin br_161
* pin bl_162
* pin br_162
* pin bl_163
* pin br_163
* pin bl_164
* pin br_164
* pin bl_165
* pin br_165
* pin bl_166
* pin br_166
* pin bl_167
* pin br_167
* pin bl_168
* pin br_168
* pin bl_169
* pin br_169
* pin bl_170
* pin br_170
* pin bl_171
* pin br_171
* pin bl_172
* pin br_172
* pin bl_173
* pin br_173
* pin bl_174
* pin br_174
* pin bl_175
* pin br_175
* pin bl_176
* pin br_176
* pin bl_177
* pin br_177
* pin bl_178
* pin br_178
* pin bl_179
* pin br_179
* pin bl_180
* pin br_180
* pin bl_181
* pin br_181
* pin bl_182
* pin br_182
* pin bl_183
* pin br_183
* pin bl_184
* pin br_184
* pin bl_185
* pin br_185
* pin bl_186
* pin br_186
* pin bl_187
* pin br_187
* pin bl_188
* pin br_188
* pin bl_189
* pin br_189
* pin bl_190
* pin br_190
* pin bl_191
* pin br_191
* pin bl_192
* pin br_192
* pin bl_193
* pin br_193
* pin bl_194
* pin br_194
* pin bl_195
* pin br_195
* pin bl_196
* pin br_196
* pin bl_197
* pin br_197
* pin bl_198
* pin br_198
* pin bl_199
* pin br_199
* pin bl_200
* pin br_200
* pin bl_201
* pin br_201
* pin bl_202
* pin br_202
* pin bl_203
* pin br_203
* pin bl_204
* pin br_204
* pin bl_205
* pin br_205
* pin bl_206
* pin br_206
* pin bl_207
* pin br_207
* pin bl_208
* pin br_208
* pin bl_209
* pin br_209
* pin bl_210
* pin br_210
* pin bl_211
* pin br_211
* pin bl_212
* pin br_212
* pin bl_213
* pin br_213
* pin bl_214
* pin br_214
* pin bl_215
* pin br_215
* pin bl_216
* pin br_216
* pin bl_217
* pin br_217
* pin bl_218
* pin br_218
* pin bl_219
* pin br_219
* pin bl_220
* pin br_220
* pin bl_221
* pin br_221
* pin bl_222
* pin br_222
* pin bl_223
* pin br_223
* pin bl_224
* pin br_224
* pin bl_225
* pin br_225
* pin bl_226
* pin br_226
* pin bl_227
* pin br_227
* pin bl_228
* pin br_228
* pin bl_229
* pin br_229
* pin bl_230
* pin br_230
* pin bl_231
* pin br_231
* pin bl_232
* pin br_232
* pin bl_233
* pin br_233
* pin bl_234
* pin br_234
* pin bl_235
* pin br_235
* pin bl_236
* pin br_236
* pin bl_237
* pin br_237
* pin bl_238
* pin br_238
* pin bl_239
* pin br_239
* pin bl_240
* pin br_240
* pin bl_241
* pin br_241
* pin bl_242
* pin br_242
* pin bl_243
* pin br_243
* pin bl_244
* pin br_244
* pin bl_245
* pin br_245
* pin bl_246
* pin br_246
* pin bl_247
* pin br_247
* pin bl_248
* pin br_248
* pin bl_249
* pin br_249
* pin bl_250
* pin br_250
* pin bl_251
* pin br_251
* pin bl_252
* pin br_252
* pin bl_253
* pin br_253
* pin bl_254
* pin br_254
* pin bl_255
* pin br_255
* pin bl_256
* pin br_256
* pin bl_257
* pin br_257
* pin vdd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_array 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147
+ 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166
+ 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185
+ 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299
+ 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318
+ 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337
+ 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356
+ 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375
+ 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394
+ 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413
+ 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432
+ 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451
+ 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470
+ 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489
+ 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508
+ 509 510 511 512 513 514 515 516 517 518
* net 1 en_bar
* net 2 bl_0
* net 3 br_0
* net 4 bl_1
* net 5 br_1
* net 6 bl_2
* net 7 br_2
* net 8 bl_3
* net 9 br_3
* net 10 bl_4
* net 11 br_4
* net 12 bl_5
* net 13 br_5
* net 14 bl_6
* net 15 br_6
* net 16 bl_7
* net 17 br_7
* net 18 bl_8
* net 19 br_8
* net 20 bl_9
* net 21 br_9
* net 22 bl_10
* net 23 br_10
* net 24 bl_11
* net 25 br_11
* net 26 bl_12
* net 27 br_12
* net 28 bl_13
* net 29 br_13
* net 30 bl_14
* net 31 br_14
* net 32 bl_15
* net 33 br_15
* net 34 bl_16
* net 35 br_16
* net 36 bl_17
* net 37 br_17
* net 38 bl_18
* net 39 br_18
* net 40 bl_19
* net 41 br_19
* net 42 bl_20
* net 43 br_20
* net 44 bl_21
* net 45 br_21
* net 46 bl_22
* net 47 br_22
* net 48 bl_23
* net 49 br_23
* net 50 bl_24
* net 51 br_24
* net 52 bl_25
* net 53 br_25
* net 54 bl_26
* net 55 br_26
* net 56 bl_27
* net 57 br_27
* net 58 bl_28
* net 59 br_28
* net 60 bl_29
* net 61 br_29
* net 62 bl_30
* net 63 br_30
* net 64 bl_31
* net 65 br_31
* net 66 bl_32
* net 67 br_32
* net 68 bl_33
* net 69 br_33
* net 70 bl_34
* net 71 br_34
* net 72 bl_35
* net 73 br_35
* net 74 bl_36
* net 75 br_36
* net 76 bl_37
* net 77 br_37
* net 78 bl_38
* net 79 br_38
* net 80 bl_39
* net 81 br_39
* net 82 bl_40
* net 83 br_40
* net 84 bl_41
* net 85 br_41
* net 86 bl_42
* net 87 br_42
* net 88 bl_43
* net 89 br_43
* net 90 bl_44
* net 91 br_44
* net 92 bl_45
* net 93 br_45
* net 94 bl_46
* net 95 br_46
* net 96 bl_47
* net 97 br_47
* net 98 bl_48
* net 99 br_48
* net 100 bl_49
* net 101 br_49
* net 102 bl_50
* net 103 br_50
* net 104 bl_51
* net 105 br_51
* net 106 bl_52
* net 107 br_52
* net 108 bl_53
* net 109 br_53
* net 110 bl_54
* net 111 br_54
* net 112 bl_55
* net 113 br_55
* net 114 bl_56
* net 115 br_56
* net 116 bl_57
* net 117 br_57
* net 118 bl_58
* net 119 br_58
* net 120 bl_59
* net 121 br_59
* net 122 bl_60
* net 123 br_60
* net 124 bl_61
* net 125 br_61
* net 126 bl_62
* net 127 br_62
* net 128 bl_63
* net 129 br_63
* net 130 bl_64
* net 131 br_64
* net 132 bl_65
* net 133 br_65
* net 134 bl_66
* net 135 br_66
* net 136 bl_67
* net 137 br_67
* net 138 bl_68
* net 139 br_68
* net 140 bl_69
* net 141 br_69
* net 142 bl_70
* net 143 br_70
* net 144 bl_71
* net 145 br_71
* net 146 bl_72
* net 147 br_72
* net 148 bl_73
* net 149 br_73
* net 150 bl_74
* net 151 br_74
* net 152 bl_75
* net 153 br_75
* net 154 bl_76
* net 155 br_76
* net 156 bl_77
* net 157 br_77
* net 158 bl_78
* net 159 br_78
* net 160 bl_79
* net 161 br_79
* net 162 bl_80
* net 163 br_80
* net 164 bl_81
* net 165 br_81
* net 166 bl_82
* net 167 br_82
* net 168 bl_83
* net 169 br_83
* net 170 bl_84
* net 171 br_84
* net 172 bl_85
* net 173 br_85
* net 174 bl_86
* net 175 br_86
* net 176 bl_87
* net 177 br_87
* net 178 bl_88
* net 179 br_88
* net 180 bl_89
* net 181 br_89
* net 182 bl_90
* net 183 br_90
* net 184 bl_91
* net 185 br_91
* net 186 bl_92
* net 187 br_92
* net 188 bl_93
* net 189 br_93
* net 190 bl_94
* net 191 br_94
* net 192 bl_95
* net 193 br_95
* net 194 bl_96
* net 195 br_96
* net 196 bl_97
* net 197 br_97
* net 198 bl_98
* net 199 br_98
* net 200 bl_99
* net 201 br_99
* net 202 bl_100
* net 203 br_100
* net 204 bl_101
* net 205 br_101
* net 206 bl_102
* net 207 br_102
* net 208 bl_103
* net 209 br_103
* net 210 bl_104
* net 211 br_104
* net 212 bl_105
* net 213 br_105
* net 214 bl_106
* net 215 br_106
* net 216 bl_107
* net 217 br_107
* net 218 bl_108
* net 219 br_108
* net 220 bl_109
* net 221 br_109
* net 222 bl_110
* net 223 br_110
* net 224 bl_111
* net 225 br_111
* net 226 bl_112
* net 227 br_112
* net 228 bl_113
* net 229 br_113
* net 230 bl_114
* net 231 br_114
* net 232 bl_115
* net 233 br_115
* net 234 bl_116
* net 235 br_116
* net 236 bl_117
* net 237 br_117
* net 238 bl_118
* net 239 br_118
* net 240 bl_119
* net 241 br_119
* net 242 bl_120
* net 243 br_120
* net 244 bl_121
* net 245 br_121
* net 246 bl_122
* net 247 br_122
* net 248 bl_123
* net 249 br_123
* net 250 bl_124
* net 251 br_124
* net 252 bl_125
* net 253 br_125
* net 254 bl_126
* net 255 br_126
* net 256 bl_127
* net 257 br_127
* net 258 bl_128
* net 259 br_128
* net 260 bl_129
* net 261 br_129
* net 262 bl_130
* net 263 br_130
* net 264 bl_131
* net 265 br_131
* net 266 bl_132
* net 267 br_132
* net 268 bl_133
* net 269 br_133
* net 270 bl_134
* net 271 br_134
* net 272 bl_135
* net 273 br_135
* net 274 bl_136
* net 275 br_136
* net 276 bl_137
* net 277 br_137
* net 278 bl_138
* net 279 br_138
* net 280 bl_139
* net 281 br_139
* net 282 bl_140
* net 283 br_140
* net 284 bl_141
* net 285 br_141
* net 286 bl_142
* net 287 br_142
* net 288 bl_143
* net 289 br_143
* net 290 bl_144
* net 291 br_144
* net 292 bl_145
* net 293 br_145
* net 294 bl_146
* net 295 br_146
* net 296 bl_147
* net 297 br_147
* net 298 bl_148
* net 299 br_148
* net 300 bl_149
* net 301 br_149
* net 302 bl_150
* net 303 br_150
* net 304 bl_151
* net 305 br_151
* net 306 bl_152
* net 307 br_152
* net 308 bl_153
* net 309 br_153
* net 310 bl_154
* net 311 br_154
* net 312 bl_155
* net 313 br_155
* net 314 bl_156
* net 315 br_156
* net 316 bl_157
* net 317 br_157
* net 318 bl_158
* net 319 br_158
* net 320 bl_159
* net 321 br_159
* net 322 bl_160
* net 323 br_160
* net 324 bl_161
* net 325 br_161
* net 326 bl_162
* net 327 br_162
* net 328 bl_163
* net 329 br_163
* net 330 bl_164
* net 331 br_164
* net 332 bl_165
* net 333 br_165
* net 334 bl_166
* net 335 br_166
* net 336 bl_167
* net 337 br_167
* net 338 bl_168
* net 339 br_168
* net 340 bl_169
* net 341 br_169
* net 342 bl_170
* net 343 br_170
* net 344 bl_171
* net 345 br_171
* net 346 bl_172
* net 347 br_172
* net 348 bl_173
* net 349 br_173
* net 350 bl_174
* net 351 br_174
* net 352 bl_175
* net 353 br_175
* net 354 bl_176
* net 355 br_176
* net 356 bl_177
* net 357 br_177
* net 358 bl_178
* net 359 br_178
* net 360 bl_179
* net 361 br_179
* net 362 bl_180
* net 363 br_180
* net 364 bl_181
* net 365 br_181
* net 366 bl_182
* net 367 br_182
* net 368 bl_183
* net 369 br_183
* net 370 bl_184
* net 371 br_184
* net 372 bl_185
* net 373 br_185
* net 374 bl_186
* net 375 br_186
* net 376 bl_187
* net 377 br_187
* net 378 bl_188
* net 379 br_188
* net 380 bl_189
* net 381 br_189
* net 382 bl_190
* net 383 br_190
* net 384 bl_191
* net 385 br_191
* net 386 bl_192
* net 387 br_192
* net 388 bl_193
* net 389 br_193
* net 390 bl_194
* net 391 br_194
* net 392 bl_195
* net 393 br_195
* net 394 bl_196
* net 395 br_196
* net 396 bl_197
* net 397 br_197
* net 398 bl_198
* net 399 br_198
* net 400 bl_199
* net 401 br_199
* net 402 bl_200
* net 403 br_200
* net 404 bl_201
* net 405 br_201
* net 406 bl_202
* net 407 br_202
* net 408 bl_203
* net 409 br_203
* net 410 bl_204
* net 411 br_204
* net 412 bl_205
* net 413 br_205
* net 414 bl_206
* net 415 br_206
* net 416 bl_207
* net 417 br_207
* net 418 bl_208
* net 419 br_208
* net 420 bl_209
* net 421 br_209
* net 422 bl_210
* net 423 br_210
* net 424 bl_211
* net 425 br_211
* net 426 bl_212
* net 427 br_212
* net 428 bl_213
* net 429 br_213
* net 430 bl_214
* net 431 br_214
* net 432 bl_215
* net 433 br_215
* net 434 bl_216
* net 435 br_216
* net 436 bl_217
* net 437 br_217
* net 438 bl_218
* net 439 br_218
* net 440 bl_219
* net 441 br_219
* net 442 bl_220
* net 443 br_220
* net 444 bl_221
* net 445 br_221
* net 446 bl_222
* net 447 br_222
* net 448 bl_223
* net 449 br_223
* net 450 bl_224
* net 451 br_224
* net 452 bl_225
* net 453 br_225
* net 454 bl_226
* net 455 br_226
* net 456 bl_227
* net 457 br_227
* net 458 bl_228
* net 459 br_228
* net 460 bl_229
* net 461 br_229
* net 462 bl_230
* net 463 br_230
* net 464 bl_231
* net 465 br_231
* net 466 bl_232
* net 467 br_232
* net 468 bl_233
* net 469 br_233
* net 470 bl_234
* net 471 br_234
* net 472 bl_235
* net 473 br_235
* net 474 bl_236
* net 475 br_236
* net 476 bl_237
* net 477 br_237
* net 478 bl_238
* net 479 br_238
* net 480 bl_239
* net 481 br_239
* net 482 bl_240
* net 483 br_240
* net 484 bl_241
* net 485 br_241
* net 486 bl_242
* net 487 br_242
* net 488 bl_243
* net 489 br_243
* net 490 bl_244
* net 491 br_244
* net 492 bl_245
* net 493 br_245
* net 494 bl_246
* net 495 br_246
* net 496 bl_247
* net 497 br_247
* net 498 bl_248
* net 499 br_248
* net 500 bl_249
* net 501 br_249
* net 502 bl_250
* net 503 br_250
* net 504 bl_251
* net 505 br_251
* net 506 bl_252
* net 507 br_252
* net 508 bl_253
* net 509 br_253
* net 510 bl_254
* net 511 br_254
* net 512 bl_255
* net 513 br_255
* net 514 bl_256
* net 515 br_256
* net 516 bl_257
* net 517 br_257
* net 518 vdd
* cell instance $1 r0 *1 1.64,0
X$1 1 2 3 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $2 r0 *1 2.345,0
X$2 1 4 5 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $3 r0 *1 3.05,0
X$3 1 6 7 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $4 r0 *1 3.755,0
X$4 1 8 9 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $5 r0 *1 4.46,0
X$5 1 10 11 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $6 r0 *1 5.165,0
X$6 1 12 13 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $7 r0 *1 5.87,0
X$7 1 14 15 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $8 r0 *1 6.575,0
X$8 1 16 17 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $9 r0 *1 7.28,0
X$9 1 18 19 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $10 r0 *1 7.985,0
X$10 1 20 21 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $11 r0 *1 8.69,0
X$11 1 22 23 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $12 r0 *1 9.395,0
X$12 1 24 25 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $13 r0 *1 10.1,0
X$13 1 26 27 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $14 r0 *1 10.805,0
X$14 1 28 29 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $15 r0 *1 11.51,0
X$15 1 30 31 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $16 r0 *1 12.215,0
X$16 1 32 33 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $17 r0 *1 12.92,0
X$17 1 34 35 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $18 r0 *1 13.625,0
X$18 1 36 37 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $19 r0 *1 14.33,0
X$19 1 38 39 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $20 r0 *1 15.035,0
X$20 1 40 41 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $21 r0 *1 15.74,0
X$21 1 42 43 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $22 r0 *1 16.445,0
X$22 1 44 45 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $23 r0 *1 17.15,0
X$23 1 46 47 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $24 r0 *1 17.855,0
X$24 1 48 49 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $25 r0 *1 18.56,0
X$25 1 50 51 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $26 r0 *1 19.265,0
X$26 1 52 53 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $27 r0 *1 19.97,0
X$27 1 54 55 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $28 r0 *1 20.675,0
X$28 1 56 57 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $29 r0 *1 21.38,0
X$29 1 58 59 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $30 r0 *1 22.085,0
X$30 1 60 61 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $31 r0 *1 22.79,0
X$31 1 62 63 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $32 r0 *1 23.495,0
X$32 1 64 65 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $33 r0 *1 24.2,0
X$33 1 66 67 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $34 r0 *1 24.905,0
X$34 1 68 69 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $35 r0 *1 25.61,0
X$35 1 70 71 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $36 r0 *1 26.315,0
X$36 1 72 73 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $37 r0 *1 27.02,0
X$37 1 74 75 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $38 r0 *1 27.725,0
X$38 1 76 77 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $39 r0 *1 28.43,0
X$39 1 78 79 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $40 r0 *1 29.135,0
X$40 1 80 81 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $41 r0 *1 29.84,0
X$41 1 82 83 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $42 r0 *1 30.545,0
X$42 1 84 85 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $43 r0 *1 31.25,0
X$43 1 86 87 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $44 r0 *1 31.955,0
X$44 1 88 89 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $45 r0 *1 32.66,0
X$45 1 90 91 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $46 r0 *1 33.365,0
X$46 1 92 93 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $47 r0 *1 34.07,0
X$47 1 94 95 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $48 r0 *1 34.775,0
X$48 1 96 97 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $49 r0 *1 35.48,0
X$49 1 98 99 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $50 r0 *1 36.185,0
X$50 1 100 101 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $51 r0 *1 36.89,0
X$51 1 102 103 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $52 r0 *1 37.595,0
X$52 1 104 105 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $53 r0 *1 38.3,0
X$53 1 106 107 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $54 r0 *1 39.005,0
X$54 1 108 109 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $55 r0 *1 39.71,0
X$55 1 110 111 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $56 r0 *1 40.415,0
X$56 1 112 113 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $57 r0 *1 41.12,0
X$57 1 114 115 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $58 r0 *1 41.825,0
X$58 1 116 117 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $59 r0 *1 42.53,0
X$59 1 118 119 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $60 r0 *1 43.235,0
X$60 1 120 121 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $61 r0 *1 43.94,0
X$61 1 122 123 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $62 r0 *1 44.645,0
X$62 1 124 125 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $63 r0 *1 45.35,0
X$63 1 126 127 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $64 r0 *1 46.055,0
X$64 1 128 129 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $65 r0 *1 46.76,0
X$65 1 130 131 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $66 r0 *1 47.465,0
X$66 1 132 133 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $67 r0 *1 48.17,0
X$67 1 134 135 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $68 r0 *1 48.875,0
X$68 1 136 137 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $69 r0 *1 49.58,0
X$69 1 138 139 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $70 r0 *1 50.285,0
X$70 1 140 141 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $71 r0 *1 50.99,0
X$71 1 142 143 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $72 r0 *1 51.695,0
X$72 1 144 145 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $73 r0 *1 52.4,0
X$73 1 146 147 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $74 r0 *1 53.105,0
X$74 1 148 149 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $75 r0 *1 53.81,0
X$75 1 150 151 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $76 r0 *1 54.515,0
X$76 1 152 153 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $77 r0 *1 55.22,0
X$77 1 154 155 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $78 r0 *1 55.925,0
X$78 1 156 157 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $79 r0 *1 56.63,0
X$79 1 158 159 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $80 r0 *1 57.335,0
X$80 1 160 161 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $81 r0 *1 58.04,0
X$81 1 162 163 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $82 r0 *1 58.745,0
X$82 1 164 165 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $83 r0 *1 59.45,0
X$83 1 166 167 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $84 r0 *1 60.155,0
X$84 1 168 169 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $85 r0 *1 60.86,0
X$85 1 170 171 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $86 r0 *1 61.565,0
X$86 1 172 173 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $87 r0 *1 62.27,0
X$87 1 174 175 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $88 r0 *1 62.975,0
X$88 1 176 177 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $89 r0 *1 63.68,0
X$89 1 178 179 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $90 r0 *1 64.385,0
X$90 1 180 181 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $91 r0 *1 65.09,0
X$91 1 182 183 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $92 r0 *1 65.795,0
X$92 1 184 185 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $93 r0 *1 66.5,0
X$93 1 186 187 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $94 r0 *1 67.205,0
X$94 1 188 189 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $95 r0 *1 67.91,0
X$95 1 190 191 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $96 r0 *1 68.615,0
X$96 1 192 193 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $97 r0 *1 69.32,0
X$97 1 194 195 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $98 r0 *1 70.025,0
X$98 1 196 197 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $99 r0 *1 70.73,0
X$99 1 198 199 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $100 r0 *1 71.435,0
X$100 1 200 201 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $101 r0 *1 72.14,0
X$101 1 202 203 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $102 r0 *1 72.845,0
X$102 1 204 205 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $103 r0 *1 73.55,0
X$103 1 206 207 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $104 r0 *1 74.255,0
X$104 1 208 209 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $105 r0 *1 74.96,0
X$105 1 210 211 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $106 r0 *1 75.665,0
X$106 1 212 213 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $107 r0 *1 76.37,0
X$107 1 214 215 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $108 r0 *1 77.075,0
X$108 1 216 217 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $109 r0 *1 77.78,0
X$109 1 218 219 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $110 r0 *1 78.485,0
X$110 1 220 221 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $111 r0 *1 79.19,0
X$111 1 222 223 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $112 r0 *1 79.895,0
X$112 1 224 225 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $113 r0 *1 80.6,0
X$113 1 226 227 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $114 r0 *1 81.305,0
X$114 1 228 229 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $115 r0 *1 82.01,0
X$115 1 230 231 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $116 r0 *1 82.715,0
X$116 1 232 233 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $117 r0 *1 83.42,0
X$117 1 234 235 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $118 r0 *1 84.125,0
X$118 1 236 237 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $119 r0 *1 84.83,0
X$119 1 238 239 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $120 r0 *1 85.535,0
X$120 1 240 241 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $121 r0 *1 86.24,0
X$121 1 242 243 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $122 r0 *1 86.945,0
X$122 1 244 245 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $123 r0 *1 87.65,0
X$123 1 246 247 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $124 r0 *1 88.355,0
X$124 1 248 249 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $125 r0 *1 89.06,0
X$125 1 250 251 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $126 r0 *1 89.765,0
X$126 1 252 253 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $127 r0 *1 90.47,0
X$127 1 254 255 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $128 r0 *1 91.175,0
X$128 1 256 257 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $129 r0 *1 91.88,0
X$129 1 258 259 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $130 r0 *1 92.585,0
X$130 1 260 261 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $131 r0 *1 93.29,0
X$131 1 262 263 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $132 r0 *1 93.995,0
X$132 1 264 265 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $133 r0 *1 94.7,0
X$133 1 266 267 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $134 r0 *1 95.405,0
X$134 1 268 269 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $135 r0 *1 96.11,0
X$135 1 270 271 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $136 r0 *1 96.815,0
X$136 1 272 273 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $137 r0 *1 97.52,0
X$137 1 274 275 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $138 r0 *1 98.225,0
X$138 1 276 277 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $139 r0 *1 98.93,0
X$139 1 278 279 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $140 r0 *1 99.635,0
X$140 1 280 281 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $141 r0 *1 100.34,0
X$141 1 282 283 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $142 r0 *1 101.045,0
X$142 1 284 285 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $143 r0 *1 101.75,0
X$143 1 286 287 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $144 r0 *1 102.455,0
X$144 1 288 289 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $145 r0 *1 103.16,0
X$145 1 290 291 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $146 r0 *1 103.865,0
X$146 1 292 293 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $147 r0 *1 104.57,0
X$147 1 294 295 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $148 r0 *1 105.275,0
X$148 1 296 297 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $149 r0 *1 105.98,0
X$149 1 298 299 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $150 r0 *1 106.685,0
X$150 1 300 301 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $151 r0 *1 107.39,0
X$151 1 302 303 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $152 r0 *1 108.095,0
X$152 1 304 305 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $153 r0 *1 108.8,0
X$153 1 306 307 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $154 r0 *1 109.505,0
X$154 1 308 309 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $155 r0 *1 110.21,0
X$155 1 310 311 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $156 r0 *1 110.915,0
X$156 1 312 313 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $157 r0 *1 111.62,0
X$157 1 314 315 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $158 r0 *1 112.325,0
X$158 1 316 317 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $159 r0 *1 113.03,0
X$159 1 318 319 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $160 r0 *1 113.735,0
X$160 1 320 321 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $161 r0 *1 114.44,0
X$161 1 322 323 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $162 r0 *1 115.145,0
X$162 1 324 325 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $163 r0 *1 115.85,0
X$163 1 326 327 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $164 r0 *1 116.555,0
X$164 1 328 329 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $165 r0 *1 117.26,0
X$165 1 330 331 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $166 r0 *1 117.965,0
X$166 1 332 333 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $167 r0 *1 118.67,0
X$167 1 334 335 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $168 r0 *1 119.375,0
X$168 1 336 337 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $169 r0 *1 120.08,0
X$169 1 338 339 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $170 r0 *1 120.785,0
X$170 1 340 341 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $171 r0 *1 121.49,0
X$171 1 342 343 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $172 r0 *1 122.195,0
X$172 1 344 345 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $173 r0 *1 122.9,0
X$173 1 346 347 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $174 r0 *1 123.605,0
X$174 1 348 349 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $175 r0 *1 124.31,0
X$175 1 350 351 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $176 r0 *1 125.015,0
X$176 1 352 353 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $177 r0 *1 125.72,0
X$177 1 354 355 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $178 r0 *1 126.425,0
X$178 1 356 357 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $179 r0 *1 127.13,0
X$179 1 358 359 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $180 r0 *1 127.835,0
X$180 1 360 361 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $181 r0 *1 128.54,0
X$181 1 362 363 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $182 r0 *1 129.245,0
X$182 1 364 365 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $183 r0 *1 129.95,0
X$183 1 366 367 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $184 r0 *1 130.655,0
X$184 1 368 369 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $185 r0 *1 131.36,0
X$185 1 370 371 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $186 r0 *1 132.065,0
X$186 1 372 373 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $187 r0 *1 132.77,0
X$187 1 374 375 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $188 r0 *1 133.475,0
X$188 1 376 377 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $189 r0 *1 134.18,0
X$189 1 378 379 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $190 r0 *1 134.885,0
X$190 1 380 381 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $191 r0 *1 135.59,0
X$191 1 382 383 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $192 r0 *1 136.295,0
X$192 1 384 385 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $193 r0 *1 137,0
X$193 1 386 387 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $194 r0 *1 137.705,0
X$194 1 388 389 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $195 r0 *1 138.41,0
X$195 1 390 391 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $196 r0 *1 139.115,0
X$196 1 392 393 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $197 r0 *1 139.82,0
X$197 1 394 395 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $198 r0 *1 140.525,0
X$198 1 396 397 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $199 r0 *1 141.23,0
X$199 1 398 399 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $200 r0 *1 141.935,0
X$200 1 400 401 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $201 r0 *1 142.64,0
X$201 1 402 403 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $202 r0 *1 143.345,0
X$202 1 404 405 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $203 r0 *1 144.05,0
X$203 1 406 407 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $204 r0 *1 144.755,0
X$204 1 408 409 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $205 r0 *1 145.46,0
X$205 1 410 411 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $206 r0 *1 146.165,0
X$206 1 412 413 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $207 r0 *1 146.87,0
X$207 1 414 415 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $208 r0 *1 147.575,0
X$208 1 416 417 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $209 r0 *1 148.28,0
X$209 1 418 419 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $210 r0 *1 148.985,0
X$210 1 420 421 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $211 r0 *1 149.69,0
X$211 1 422 423 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $212 r0 *1 150.395,0
X$212 1 424 425 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $213 r0 *1 151.1,0
X$213 1 426 427 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $214 r0 *1 151.805,0
X$214 1 428 429 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $215 r0 *1 152.51,0
X$215 1 430 431 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $216 r0 *1 153.215,0
X$216 1 432 433 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $217 r0 *1 153.92,0
X$217 1 434 435 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $218 r0 *1 154.625,0
X$218 1 436 437 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $219 r0 *1 155.33,0
X$219 1 438 439 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $220 r0 *1 156.035,0
X$220 1 440 441 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $221 r0 *1 156.74,0
X$221 1 442 443 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $222 r0 *1 157.445,0
X$222 1 444 445 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $223 r0 *1 158.15,0
X$223 1 446 447 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $224 r0 *1 158.855,0
X$224 1 448 449 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $225 r0 *1 159.56,0
X$225 1 450 451 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $226 r0 *1 160.265,0
X$226 1 452 453 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $227 r0 *1 160.97,0
X$227 1 454 455 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $228 r0 *1 161.675,0
X$228 1 456 457 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $229 r0 *1 162.38,0
X$229 1 458 459 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $230 r0 *1 163.085,0
X$230 1 460 461 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $231 r0 *1 163.79,0
X$231 1 462 463 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $232 r0 *1 164.495,0
X$232 1 464 465 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $233 r0 *1 165.2,0
X$233 1 466 467 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $234 r0 *1 165.905,0
X$234 1 468 469 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $235 r0 *1 166.61,0
X$235 1 470 471 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $236 r0 *1 167.315,0
X$236 1 472 473 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $237 r0 *1 168.02,0
X$237 1 474 475 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $238 r0 *1 168.725,0
X$238 1 476 477 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $239 r0 *1 169.43,0
X$239 1 478 479 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $240 r0 *1 170.135,0
X$240 1 480 481 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $241 r0 *1 170.84,0
X$241 1 482 483 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $242 r0 *1 171.545,0
X$242 1 484 485 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $243 r0 *1 172.25,0
X$243 1 486 487 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $244 r0 *1 172.955,0
X$244 1 488 489 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $245 r0 *1 173.66,0
X$245 1 490 491 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $246 r0 *1 174.365,0
X$246 1 492 493 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $247 r0 *1 175.07,0
X$247 1 494 495 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $248 r0 *1 175.775,0
X$248 1 496 497 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $249 r0 *1 176.48,0
X$249 1 498 499 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $250 r0 *1 177.185,0
X$250 1 500 501 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $251 r0 *1 177.89,0
X$251 1 502 503 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $252 r0 *1 178.595,0
X$252 1 504 505 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $253 r0 *1 179.3,0
X$253 1 506 507 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $254 r0 *1 180.005,0
X$254 1 508 509 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $255 r0 *1 180.71,0
X$255 1 510 511 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $256 r0 *1 181.415,0
X$256 1 512 513 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $257 r0 *1 182.12,0
X$257 1 514 515 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* cell instance $258 r0 *1 182.825,0
X$258 1 516 517 518 freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_3
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_24
* pin wl_0_25
* pin wl_0_26
* pin wl_0_27
* pin wl_0_28
* pin wl_0_29
* pin wl_0_30
* pin wl_0_31
* pin wl_0_32
* pin wl_0_33
* pin wl_0_34
* pin wl_0_35
* pin wl_0_36
* pin wl_0_37
* pin wl_0_38
* pin wl_0_39
* pin wl_0_40
* pin wl_0_41
* pin wl_0_42
* pin wl_0_43
* pin wl_0_44
* pin wl_0_45
* pin wl_0_46
* pin wl_0_47
* pin wl_0_48
* pin wl_0_49
* pin wl_0_50
* pin wl_0_51
* pin wl_0_52
* pin wl_0_53
* pin wl_0_54
* pin wl_0_55
* pin wl_0_56
* pin wl_0_57
* pin wl_0_58
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_62
* pin wl_0_63
* pin wl_0_64
* pin wl_0_65
* pin wl_0_66
* pin wl_0_67
* pin wl_0_68
* pin wl_0_69
* pin wl_0_70
* pin wl_0_71
* pin wl_0_72
* pin wl_0_73
* pin wl_0_74
* pin wl_0_75
* pin wl_0_76
* pin wl_0_77
* pin wl_0_78
* pin wl_0_79
* pin wl_0_80
* pin wl_0_81
* pin wl_0_82
* pin wl_0_83
* pin wl_0_84
* pin wl_0_85
* pin wl_0_86
* pin wl_0_87
* pin wl_0_88
* pin wl_0_89
* pin wl_0_90
* pin wl_0_91
* pin wl_0_92
* pin wl_0_93
* pin wl_0_94
* pin wl_0_95
* pin wl_0_96
* pin wl_0_97
* pin wl_0_98
* pin wl_0_99
* pin wl_0_100
* pin wl_0_101
* pin wl_0_102
* pin wl_0_103
* pin wl_0_104
* pin wl_0_105
* pin wl_0_106
* pin wl_0_107
* pin wl_0_108
* pin wl_0_109
* pin wl_0_110
* pin wl_0_111
* pin wl_0_112
* pin wl_0_113
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_117
* pin wl_0_118
* pin wl_0_119
* pin wl_0_120
* pin wl_0_121
* pin wl_0_122
* pin wl_0_123
* pin wl_0_124
* pin wl_0_125
* pin wl_0_126
* pin wl_0_127
* pin wl_0_128
* pin wl_0_129
* pin wl_0_130
* pin wl_0_131
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_3 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 wl_0_19
* net 21 wl_0_20
* net 22 wl_0_21
* net 23 wl_0_22
* net 24 wl_0_23
* net 25 wl_0_24
* net 26 wl_0_25
* net 27 wl_0_26
* net 28 wl_0_27
* net 29 wl_0_28
* net 30 wl_0_29
* net 31 wl_0_30
* net 32 wl_0_31
* net 33 wl_0_32
* net 34 wl_0_33
* net 35 wl_0_34
* net 36 wl_0_35
* net 37 wl_0_36
* net 38 wl_0_37
* net 39 wl_0_38
* net 40 wl_0_39
* net 41 wl_0_40
* net 42 wl_0_41
* net 43 wl_0_42
* net 44 wl_0_43
* net 45 wl_0_44
* net 46 wl_0_45
* net 47 wl_0_46
* net 48 wl_0_47
* net 49 wl_0_48
* net 50 wl_0_49
* net 51 wl_0_50
* net 52 wl_0_51
* net 53 wl_0_52
* net 54 wl_0_53
* net 55 wl_0_54
* net 56 wl_0_55
* net 57 wl_0_56
* net 58 wl_0_57
* net 59 wl_0_58
* net 60 wl_0_59
* net 61 wl_0_60
* net 62 wl_0_61
* net 63 wl_0_62
* net 64 wl_0_63
* net 65 wl_0_64
* net 66 wl_0_65
* net 67 wl_0_66
* net 68 wl_0_67
* net 69 wl_0_68
* net 70 wl_0_69
* net 71 wl_0_70
* net 72 wl_0_71
* net 73 wl_0_72
* net 74 wl_0_73
* net 75 wl_0_74
* net 76 wl_0_75
* net 77 wl_0_76
* net 78 wl_0_77
* net 79 wl_0_78
* net 80 wl_0_79
* net 81 wl_0_80
* net 82 wl_0_81
* net 83 wl_0_82
* net 84 wl_0_83
* net 85 wl_0_84
* net 86 wl_0_85
* net 87 wl_0_86
* net 88 wl_0_87
* net 89 wl_0_88
* net 90 wl_0_89
* net 91 wl_0_90
* net 92 wl_0_91
* net 93 wl_0_92
* net 94 wl_0_93
* net 95 wl_0_94
* net 96 wl_0_95
* net 97 wl_0_96
* net 98 wl_0_97
* net 99 wl_0_98
* net 100 wl_0_99
* net 101 wl_0_100
* net 102 wl_0_101
* net 103 wl_0_102
* net 104 wl_0_103
* net 105 wl_0_104
* net 106 wl_0_105
* net 107 wl_0_106
* net 108 wl_0_107
* net 109 wl_0_108
* net 110 wl_0_109
* net 111 wl_0_110
* net 112 wl_0_111
* net 113 wl_0_112
* net 114 wl_0_113
* net 115 wl_0_114
* net 116 wl_0_115
* net 117 wl_0_116
* net 118 wl_0_117
* net 119 wl_0_118
* net 120 wl_0_119
* net 121 wl_0_120
* net 122 wl_0_121
* net 123 wl_0_122
* net 124 wl_0_123
* net 125 wl_0_124
* net 126 wl_0_125
* net 127 wl_0_126
* net 128 wl_0_127
* net 129 wl_0_128
* net 130 wl_0_129
* net 131 wl_0_130
* net 132 wl_0_131
* net 133 vdd
* net 134 gnd
* cell instance $1 r0 *1 0,0
X$1 1 133 134 dummy_cell_1rw
* cell instance $2 m0 *1 0,2.73
X$2 2 133 134 dummy_cell_1rw
* cell instance $3 r0 *1 0,2.73
X$3 3 133 134 dummy_cell_1rw
* cell instance $4 m0 *1 0,5.46
X$4 4 133 134 dummy_cell_1rw
* cell instance $5 r0 *1 0,5.46
X$5 5 133 134 dummy_cell_1rw
* cell instance $6 m0 *1 0,8.19
X$6 6 133 134 dummy_cell_1rw
* cell instance $7 r0 *1 0,8.19
X$7 7 133 134 dummy_cell_1rw
* cell instance $8 m0 *1 0,10.92
X$8 8 133 134 dummy_cell_1rw
* cell instance $9 r0 *1 0,10.92
X$9 9 133 134 dummy_cell_1rw
* cell instance $10 m0 *1 0,13.65
X$10 10 133 134 dummy_cell_1rw
* cell instance $11 r0 *1 0,13.65
X$11 11 133 134 dummy_cell_1rw
* cell instance $12 m0 *1 0,16.38
X$12 12 133 134 dummy_cell_1rw
* cell instance $13 r0 *1 0,16.38
X$13 13 133 134 dummy_cell_1rw
* cell instance $14 m0 *1 0,19.11
X$14 14 133 134 dummy_cell_1rw
* cell instance $15 r0 *1 0,19.11
X$15 15 133 134 dummy_cell_1rw
* cell instance $16 m0 *1 0,21.84
X$16 16 133 134 dummy_cell_1rw
* cell instance $17 r0 *1 0,21.84
X$17 17 133 134 dummy_cell_1rw
* cell instance $18 m0 *1 0,24.57
X$18 18 133 134 dummy_cell_1rw
* cell instance $19 r0 *1 0,24.57
X$19 19 133 134 dummy_cell_1rw
* cell instance $20 m0 *1 0,27.3
X$20 20 133 134 dummy_cell_1rw
* cell instance $21 r0 *1 0,27.3
X$21 21 133 134 dummy_cell_1rw
* cell instance $22 m0 *1 0,30.03
X$22 22 133 134 dummy_cell_1rw
* cell instance $23 r0 *1 0,30.03
X$23 23 133 134 dummy_cell_1rw
* cell instance $24 m0 *1 0,32.76
X$24 24 133 134 dummy_cell_1rw
* cell instance $25 r0 *1 0,32.76
X$25 25 133 134 dummy_cell_1rw
* cell instance $26 m0 *1 0,35.49
X$26 26 133 134 dummy_cell_1rw
* cell instance $27 r0 *1 0,35.49
X$27 27 133 134 dummy_cell_1rw
* cell instance $28 m0 *1 0,38.22
X$28 28 133 134 dummy_cell_1rw
* cell instance $29 r0 *1 0,38.22
X$29 29 133 134 dummy_cell_1rw
* cell instance $30 m0 *1 0,40.95
X$30 30 133 134 dummy_cell_1rw
* cell instance $31 r0 *1 0,40.95
X$31 31 133 134 dummy_cell_1rw
* cell instance $32 m0 *1 0,43.68
X$32 32 133 134 dummy_cell_1rw
* cell instance $33 r0 *1 0,43.68
X$33 33 133 134 dummy_cell_1rw
* cell instance $34 m0 *1 0,46.41
X$34 34 133 134 dummy_cell_1rw
* cell instance $35 r0 *1 0,46.41
X$35 35 133 134 dummy_cell_1rw
* cell instance $36 m0 *1 0,49.14
X$36 36 133 134 dummy_cell_1rw
* cell instance $37 r0 *1 0,49.14
X$37 37 133 134 dummy_cell_1rw
* cell instance $38 m0 *1 0,51.87
X$38 38 133 134 dummy_cell_1rw
* cell instance $39 r0 *1 0,51.87
X$39 39 133 134 dummy_cell_1rw
* cell instance $40 m0 *1 0,54.6
X$40 40 133 134 dummy_cell_1rw
* cell instance $41 r0 *1 0,54.6
X$41 41 133 134 dummy_cell_1rw
* cell instance $42 m0 *1 0,57.33
X$42 42 133 134 dummy_cell_1rw
* cell instance $43 r0 *1 0,57.33
X$43 43 133 134 dummy_cell_1rw
* cell instance $44 m0 *1 0,60.06
X$44 44 133 134 dummy_cell_1rw
* cell instance $45 r0 *1 0,60.06
X$45 45 133 134 dummy_cell_1rw
* cell instance $46 m0 *1 0,62.79
X$46 46 133 134 dummy_cell_1rw
* cell instance $47 r0 *1 0,62.79
X$47 47 133 134 dummy_cell_1rw
* cell instance $48 m0 *1 0,65.52
X$48 48 133 134 dummy_cell_1rw
* cell instance $49 r0 *1 0,65.52
X$49 49 133 134 dummy_cell_1rw
* cell instance $50 m0 *1 0,68.25
X$50 50 133 134 dummy_cell_1rw
* cell instance $51 r0 *1 0,68.25
X$51 51 133 134 dummy_cell_1rw
* cell instance $52 m0 *1 0,70.98
X$52 52 133 134 dummy_cell_1rw
* cell instance $53 r0 *1 0,70.98
X$53 53 133 134 dummy_cell_1rw
* cell instance $54 m0 *1 0,73.71
X$54 54 133 134 dummy_cell_1rw
* cell instance $55 r0 *1 0,73.71
X$55 55 133 134 dummy_cell_1rw
* cell instance $56 m0 *1 0,76.44
X$56 56 133 134 dummy_cell_1rw
* cell instance $57 r0 *1 0,76.44
X$57 57 133 134 dummy_cell_1rw
* cell instance $58 m0 *1 0,79.17
X$58 58 133 134 dummy_cell_1rw
* cell instance $59 r0 *1 0,79.17
X$59 59 133 134 dummy_cell_1rw
* cell instance $60 m0 *1 0,81.9
X$60 60 133 134 dummy_cell_1rw
* cell instance $61 r0 *1 0,81.9
X$61 61 133 134 dummy_cell_1rw
* cell instance $62 m0 *1 0,84.63
X$62 62 133 134 dummy_cell_1rw
* cell instance $63 r0 *1 0,84.63
X$63 63 133 134 dummy_cell_1rw
* cell instance $64 m0 *1 0,87.36
X$64 64 133 134 dummy_cell_1rw
* cell instance $65 r0 *1 0,87.36
X$65 65 133 134 dummy_cell_1rw
* cell instance $66 m0 *1 0,90.09
X$66 66 133 134 dummy_cell_1rw
* cell instance $67 r0 *1 0,90.09
X$67 67 133 134 dummy_cell_1rw
* cell instance $68 m0 *1 0,92.82
X$68 68 133 134 dummy_cell_1rw
* cell instance $69 r0 *1 0,92.82
X$69 69 133 134 dummy_cell_1rw
* cell instance $70 m0 *1 0,95.55
X$70 70 133 134 dummy_cell_1rw
* cell instance $71 r0 *1 0,95.55
X$71 71 133 134 dummy_cell_1rw
* cell instance $72 m0 *1 0,98.28
X$72 72 133 134 dummy_cell_1rw
* cell instance $73 r0 *1 0,98.28
X$73 73 133 134 dummy_cell_1rw
* cell instance $74 m0 *1 0,101.01
X$74 74 133 134 dummy_cell_1rw
* cell instance $75 r0 *1 0,101.01
X$75 75 133 134 dummy_cell_1rw
* cell instance $76 m0 *1 0,103.74
X$76 76 133 134 dummy_cell_1rw
* cell instance $77 r0 *1 0,103.74
X$77 77 133 134 dummy_cell_1rw
* cell instance $78 m0 *1 0,106.47
X$78 78 133 134 dummy_cell_1rw
* cell instance $79 r0 *1 0,106.47
X$79 79 133 134 dummy_cell_1rw
* cell instance $80 m0 *1 0,109.2
X$80 80 133 134 dummy_cell_1rw
* cell instance $81 r0 *1 0,109.2
X$81 81 133 134 dummy_cell_1rw
* cell instance $82 m0 *1 0,111.93
X$82 82 133 134 dummy_cell_1rw
* cell instance $83 r0 *1 0,111.93
X$83 83 133 134 dummy_cell_1rw
* cell instance $84 m0 *1 0,114.66
X$84 84 133 134 dummy_cell_1rw
* cell instance $85 r0 *1 0,114.66
X$85 85 133 134 dummy_cell_1rw
* cell instance $86 m0 *1 0,117.39
X$86 86 133 134 dummy_cell_1rw
* cell instance $87 r0 *1 0,117.39
X$87 87 133 134 dummy_cell_1rw
* cell instance $88 m0 *1 0,120.12
X$88 88 133 134 dummy_cell_1rw
* cell instance $89 r0 *1 0,120.12
X$89 89 133 134 dummy_cell_1rw
* cell instance $90 m0 *1 0,122.85
X$90 90 133 134 dummy_cell_1rw
* cell instance $91 r0 *1 0,122.85
X$91 91 133 134 dummy_cell_1rw
* cell instance $92 m0 *1 0,125.58
X$92 92 133 134 dummy_cell_1rw
* cell instance $93 r0 *1 0,125.58
X$93 93 133 134 dummy_cell_1rw
* cell instance $94 m0 *1 0,128.31
X$94 94 133 134 dummy_cell_1rw
* cell instance $95 r0 *1 0,128.31
X$95 95 133 134 dummy_cell_1rw
* cell instance $96 m0 *1 0,131.04
X$96 96 133 134 dummy_cell_1rw
* cell instance $97 r0 *1 0,131.04
X$97 97 133 134 dummy_cell_1rw
* cell instance $98 m0 *1 0,133.77
X$98 98 133 134 dummy_cell_1rw
* cell instance $99 r0 *1 0,133.77
X$99 99 133 134 dummy_cell_1rw
* cell instance $100 m0 *1 0,136.5
X$100 100 133 134 dummy_cell_1rw
* cell instance $101 r0 *1 0,136.5
X$101 101 133 134 dummy_cell_1rw
* cell instance $102 m0 *1 0,139.23
X$102 102 133 134 dummy_cell_1rw
* cell instance $103 r0 *1 0,139.23
X$103 103 133 134 dummy_cell_1rw
* cell instance $104 m0 *1 0,141.96
X$104 104 133 134 dummy_cell_1rw
* cell instance $105 r0 *1 0,141.96
X$105 105 133 134 dummy_cell_1rw
* cell instance $106 m0 *1 0,144.69
X$106 106 133 134 dummy_cell_1rw
* cell instance $107 r0 *1 0,144.69
X$107 107 133 134 dummy_cell_1rw
* cell instance $108 m0 *1 0,147.42
X$108 108 133 134 dummy_cell_1rw
* cell instance $109 r0 *1 0,147.42
X$109 109 133 134 dummy_cell_1rw
* cell instance $110 m0 *1 0,150.15
X$110 110 133 134 dummy_cell_1rw
* cell instance $111 r0 *1 0,150.15
X$111 111 133 134 dummy_cell_1rw
* cell instance $112 m0 *1 0,152.88
X$112 112 133 134 dummy_cell_1rw
* cell instance $113 r0 *1 0,152.88
X$113 113 133 134 dummy_cell_1rw
* cell instance $114 m0 *1 0,155.61
X$114 114 133 134 dummy_cell_1rw
* cell instance $115 r0 *1 0,155.61
X$115 115 133 134 dummy_cell_1rw
* cell instance $116 m0 *1 0,158.34
X$116 116 133 134 dummy_cell_1rw
* cell instance $117 r0 *1 0,158.34
X$117 117 133 134 dummy_cell_1rw
* cell instance $118 m0 *1 0,161.07
X$118 118 133 134 dummy_cell_1rw
* cell instance $119 r0 *1 0,161.07
X$119 119 133 134 dummy_cell_1rw
* cell instance $120 m0 *1 0,163.8
X$120 120 133 134 dummy_cell_1rw
* cell instance $121 r0 *1 0,163.8
X$121 121 133 134 dummy_cell_1rw
* cell instance $122 m0 *1 0,166.53
X$122 122 133 134 dummy_cell_1rw
* cell instance $123 r0 *1 0,166.53
X$123 123 133 134 dummy_cell_1rw
* cell instance $124 m0 *1 0,169.26
X$124 124 133 134 dummy_cell_1rw
* cell instance $125 r0 *1 0,169.26
X$125 125 133 134 dummy_cell_1rw
* cell instance $126 m0 *1 0,171.99
X$126 126 133 134 dummy_cell_1rw
* cell instance $127 r0 *1 0,171.99
X$127 127 133 134 dummy_cell_1rw
* cell instance $128 m0 *1 0,174.72
X$128 128 133 134 dummy_cell_1rw
* cell instance $129 r0 *1 0,174.72
X$129 129 133 134 dummy_cell_1rw
* cell instance $130 m0 *1 0,177.45
X$130 130 133 134 dummy_cell_1rw
* cell instance $131 r0 *1 0,177.45
X$131 131 133 134 dummy_cell_1rw
* cell instance $132 m0 *1 0,180.18
X$132 132 133 134 dummy_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_3

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_2
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_24
* pin wl_0_25
* pin wl_0_26
* pin wl_0_27
* pin wl_0_28
* pin wl_0_29
* pin wl_0_30
* pin wl_0_31
* pin wl_0_32
* pin wl_0_33
* pin wl_0_34
* pin wl_0_35
* pin wl_0_36
* pin wl_0_37
* pin wl_0_38
* pin wl_0_39
* pin wl_0_40
* pin wl_0_41
* pin wl_0_42
* pin wl_0_43
* pin wl_0_44
* pin wl_0_45
* pin wl_0_46
* pin wl_0_47
* pin wl_0_48
* pin wl_0_49
* pin wl_0_50
* pin wl_0_51
* pin wl_0_52
* pin wl_0_53
* pin wl_0_54
* pin wl_0_55
* pin wl_0_56
* pin wl_0_57
* pin wl_0_58
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_62
* pin wl_0_63
* pin wl_0_64
* pin wl_0_65
* pin wl_0_66
* pin wl_0_67
* pin wl_0_68
* pin wl_0_69
* pin wl_0_70
* pin wl_0_71
* pin wl_0_72
* pin wl_0_73
* pin wl_0_74
* pin wl_0_75
* pin wl_0_76
* pin wl_0_77
* pin wl_0_78
* pin wl_0_79
* pin wl_0_80
* pin wl_0_81
* pin wl_0_82
* pin wl_0_83
* pin wl_0_84
* pin wl_0_85
* pin wl_0_86
* pin wl_0_87
* pin wl_0_88
* pin wl_0_89
* pin wl_0_90
* pin wl_0_91
* pin wl_0_92
* pin wl_0_93
* pin wl_0_94
* pin wl_0_95
* pin wl_0_96
* pin wl_0_97
* pin wl_0_98
* pin wl_0_99
* pin wl_0_100
* pin wl_0_101
* pin wl_0_102
* pin wl_0_103
* pin wl_0_104
* pin wl_0_105
* pin wl_0_106
* pin wl_0_107
* pin wl_0_108
* pin wl_0_109
* pin wl_0_110
* pin wl_0_111
* pin wl_0_112
* pin wl_0_113
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_117
* pin wl_0_118
* pin wl_0_119
* pin wl_0_120
* pin wl_0_121
* pin wl_0_122
* pin wl_0_123
* pin wl_0_124
* pin wl_0_125
* pin wl_0_126
* pin wl_0_127
* pin wl_0_128
* pin wl_0_129
* pin wl_0_130
* pin wl_0_131
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_2 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 wl_0_19
* net 21 wl_0_20
* net 22 wl_0_21
* net 23 wl_0_22
* net 24 wl_0_23
* net 25 wl_0_24
* net 26 wl_0_25
* net 27 wl_0_26
* net 28 wl_0_27
* net 29 wl_0_28
* net 30 wl_0_29
* net 31 wl_0_30
* net 32 wl_0_31
* net 33 wl_0_32
* net 34 wl_0_33
* net 35 wl_0_34
* net 36 wl_0_35
* net 37 wl_0_36
* net 38 wl_0_37
* net 39 wl_0_38
* net 40 wl_0_39
* net 41 wl_0_40
* net 42 wl_0_41
* net 43 wl_0_42
* net 44 wl_0_43
* net 45 wl_0_44
* net 46 wl_0_45
* net 47 wl_0_46
* net 48 wl_0_47
* net 49 wl_0_48
* net 50 wl_0_49
* net 51 wl_0_50
* net 52 wl_0_51
* net 53 wl_0_52
* net 54 wl_0_53
* net 55 wl_0_54
* net 56 wl_0_55
* net 57 wl_0_56
* net 58 wl_0_57
* net 59 wl_0_58
* net 60 wl_0_59
* net 61 wl_0_60
* net 62 wl_0_61
* net 63 wl_0_62
* net 64 wl_0_63
* net 65 wl_0_64
* net 66 wl_0_65
* net 67 wl_0_66
* net 68 wl_0_67
* net 69 wl_0_68
* net 70 wl_0_69
* net 71 wl_0_70
* net 72 wl_0_71
* net 73 wl_0_72
* net 74 wl_0_73
* net 75 wl_0_74
* net 76 wl_0_75
* net 77 wl_0_76
* net 78 wl_0_77
* net 79 wl_0_78
* net 80 wl_0_79
* net 81 wl_0_80
* net 82 wl_0_81
* net 83 wl_0_82
* net 84 wl_0_83
* net 85 wl_0_84
* net 86 wl_0_85
* net 87 wl_0_86
* net 88 wl_0_87
* net 89 wl_0_88
* net 90 wl_0_89
* net 91 wl_0_90
* net 92 wl_0_91
* net 93 wl_0_92
* net 94 wl_0_93
* net 95 wl_0_94
* net 96 wl_0_95
* net 97 wl_0_96
* net 98 wl_0_97
* net 99 wl_0_98
* net 100 wl_0_99
* net 101 wl_0_100
* net 102 wl_0_101
* net 103 wl_0_102
* net 104 wl_0_103
* net 105 wl_0_104
* net 106 wl_0_105
* net 107 wl_0_106
* net 108 wl_0_107
* net 109 wl_0_108
* net 110 wl_0_109
* net 111 wl_0_110
* net 112 wl_0_111
* net 113 wl_0_112
* net 114 wl_0_113
* net 115 wl_0_114
* net 116 wl_0_115
* net 117 wl_0_116
* net 118 wl_0_117
* net 119 wl_0_118
* net 120 wl_0_119
* net 121 wl_0_120
* net 122 wl_0_121
* net 123 wl_0_122
* net 124 wl_0_123
* net 125 wl_0_124
* net 126 wl_0_125
* net 127 wl_0_126
* net 128 wl_0_127
* net 129 wl_0_128
* net 130 wl_0_129
* net 131 wl_0_130
* net 132 wl_0_131
* net 133 vdd
* net 134 gnd
* cell instance $1 r0 *1 0,0
X$1 1 133 134 dummy_cell_1rw
* cell instance $2 m0 *1 0,2.73
X$2 2 133 134 dummy_cell_1rw
* cell instance $3 r0 *1 0,2.73
X$3 3 133 134 dummy_cell_1rw
* cell instance $4 m0 *1 0,5.46
X$4 4 133 134 dummy_cell_1rw
* cell instance $5 r0 *1 0,5.46
X$5 5 133 134 dummy_cell_1rw
* cell instance $6 m0 *1 0,8.19
X$6 6 133 134 dummy_cell_1rw
* cell instance $7 r0 *1 0,8.19
X$7 7 133 134 dummy_cell_1rw
* cell instance $8 m0 *1 0,10.92
X$8 8 133 134 dummy_cell_1rw
* cell instance $9 r0 *1 0,10.92
X$9 9 133 134 dummy_cell_1rw
* cell instance $10 m0 *1 0,13.65
X$10 10 133 134 dummy_cell_1rw
* cell instance $11 r0 *1 0,13.65
X$11 11 133 134 dummy_cell_1rw
* cell instance $12 m0 *1 0,16.38
X$12 12 133 134 dummy_cell_1rw
* cell instance $13 r0 *1 0,16.38
X$13 13 133 134 dummy_cell_1rw
* cell instance $14 m0 *1 0,19.11
X$14 14 133 134 dummy_cell_1rw
* cell instance $15 r0 *1 0,19.11
X$15 15 133 134 dummy_cell_1rw
* cell instance $16 m0 *1 0,21.84
X$16 16 133 134 dummy_cell_1rw
* cell instance $17 r0 *1 0,21.84
X$17 17 133 134 dummy_cell_1rw
* cell instance $18 m0 *1 0,24.57
X$18 18 133 134 dummy_cell_1rw
* cell instance $19 r0 *1 0,24.57
X$19 19 133 134 dummy_cell_1rw
* cell instance $20 m0 *1 0,27.3
X$20 20 133 134 dummy_cell_1rw
* cell instance $21 r0 *1 0,27.3
X$21 21 133 134 dummy_cell_1rw
* cell instance $22 m0 *1 0,30.03
X$22 22 133 134 dummy_cell_1rw
* cell instance $23 r0 *1 0,30.03
X$23 23 133 134 dummy_cell_1rw
* cell instance $24 m0 *1 0,32.76
X$24 24 133 134 dummy_cell_1rw
* cell instance $25 r0 *1 0,32.76
X$25 25 133 134 dummy_cell_1rw
* cell instance $26 m0 *1 0,35.49
X$26 26 133 134 dummy_cell_1rw
* cell instance $27 r0 *1 0,35.49
X$27 27 133 134 dummy_cell_1rw
* cell instance $28 m0 *1 0,38.22
X$28 28 133 134 dummy_cell_1rw
* cell instance $29 r0 *1 0,38.22
X$29 29 133 134 dummy_cell_1rw
* cell instance $30 m0 *1 0,40.95
X$30 30 133 134 dummy_cell_1rw
* cell instance $31 r0 *1 0,40.95
X$31 31 133 134 dummy_cell_1rw
* cell instance $32 m0 *1 0,43.68
X$32 32 133 134 dummy_cell_1rw
* cell instance $33 r0 *1 0,43.68
X$33 33 133 134 dummy_cell_1rw
* cell instance $34 m0 *1 0,46.41
X$34 34 133 134 dummy_cell_1rw
* cell instance $35 r0 *1 0,46.41
X$35 35 133 134 dummy_cell_1rw
* cell instance $36 m0 *1 0,49.14
X$36 36 133 134 dummy_cell_1rw
* cell instance $37 r0 *1 0,49.14
X$37 37 133 134 dummy_cell_1rw
* cell instance $38 m0 *1 0,51.87
X$38 38 133 134 dummy_cell_1rw
* cell instance $39 r0 *1 0,51.87
X$39 39 133 134 dummy_cell_1rw
* cell instance $40 m0 *1 0,54.6
X$40 40 133 134 dummy_cell_1rw
* cell instance $41 r0 *1 0,54.6
X$41 41 133 134 dummy_cell_1rw
* cell instance $42 m0 *1 0,57.33
X$42 42 133 134 dummy_cell_1rw
* cell instance $43 r0 *1 0,57.33
X$43 43 133 134 dummy_cell_1rw
* cell instance $44 m0 *1 0,60.06
X$44 44 133 134 dummy_cell_1rw
* cell instance $45 r0 *1 0,60.06
X$45 45 133 134 dummy_cell_1rw
* cell instance $46 m0 *1 0,62.79
X$46 46 133 134 dummy_cell_1rw
* cell instance $47 r0 *1 0,62.79
X$47 47 133 134 dummy_cell_1rw
* cell instance $48 m0 *1 0,65.52
X$48 48 133 134 dummy_cell_1rw
* cell instance $49 r0 *1 0,65.52
X$49 49 133 134 dummy_cell_1rw
* cell instance $50 m0 *1 0,68.25
X$50 50 133 134 dummy_cell_1rw
* cell instance $51 r0 *1 0,68.25
X$51 51 133 134 dummy_cell_1rw
* cell instance $52 m0 *1 0,70.98
X$52 52 133 134 dummy_cell_1rw
* cell instance $53 r0 *1 0,70.98
X$53 53 133 134 dummy_cell_1rw
* cell instance $54 m0 *1 0,73.71
X$54 54 133 134 dummy_cell_1rw
* cell instance $55 r0 *1 0,73.71
X$55 55 133 134 dummy_cell_1rw
* cell instance $56 m0 *1 0,76.44
X$56 56 133 134 dummy_cell_1rw
* cell instance $57 r0 *1 0,76.44
X$57 57 133 134 dummy_cell_1rw
* cell instance $58 m0 *1 0,79.17
X$58 58 133 134 dummy_cell_1rw
* cell instance $59 r0 *1 0,79.17
X$59 59 133 134 dummy_cell_1rw
* cell instance $60 m0 *1 0,81.9
X$60 60 133 134 dummy_cell_1rw
* cell instance $61 r0 *1 0,81.9
X$61 61 133 134 dummy_cell_1rw
* cell instance $62 m0 *1 0,84.63
X$62 62 133 134 dummy_cell_1rw
* cell instance $63 r0 *1 0,84.63
X$63 63 133 134 dummy_cell_1rw
* cell instance $64 m0 *1 0,87.36
X$64 64 133 134 dummy_cell_1rw
* cell instance $65 r0 *1 0,87.36
X$65 65 133 134 dummy_cell_1rw
* cell instance $66 m0 *1 0,90.09
X$66 66 133 134 dummy_cell_1rw
* cell instance $67 r0 *1 0,90.09
X$67 67 133 134 dummy_cell_1rw
* cell instance $68 m0 *1 0,92.82
X$68 68 133 134 dummy_cell_1rw
* cell instance $69 r0 *1 0,92.82
X$69 69 133 134 dummy_cell_1rw
* cell instance $70 m0 *1 0,95.55
X$70 70 133 134 dummy_cell_1rw
* cell instance $71 r0 *1 0,95.55
X$71 71 133 134 dummy_cell_1rw
* cell instance $72 m0 *1 0,98.28
X$72 72 133 134 dummy_cell_1rw
* cell instance $73 r0 *1 0,98.28
X$73 73 133 134 dummy_cell_1rw
* cell instance $74 m0 *1 0,101.01
X$74 74 133 134 dummy_cell_1rw
* cell instance $75 r0 *1 0,101.01
X$75 75 133 134 dummy_cell_1rw
* cell instance $76 m0 *1 0,103.74
X$76 76 133 134 dummy_cell_1rw
* cell instance $77 r0 *1 0,103.74
X$77 77 133 134 dummy_cell_1rw
* cell instance $78 m0 *1 0,106.47
X$78 78 133 134 dummy_cell_1rw
* cell instance $79 r0 *1 0,106.47
X$79 79 133 134 dummy_cell_1rw
* cell instance $80 m0 *1 0,109.2
X$80 80 133 134 dummy_cell_1rw
* cell instance $81 r0 *1 0,109.2
X$81 81 133 134 dummy_cell_1rw
* cell instance $82 m0 *1 0,111.93
X$82 82 133 134 dummy_cell_1rw
* cell instance $83 r0 *1 0,111.93
X$83 83 133 134 dummy_cell_1rw
* cell instance $84 m0 *1 0,114.66
X$84 84 133 134 dummy_cell_1rw
* cell instance $85 r0 *1 0,114.66
X$85 85 133 134 dummy_cell_1rw
* cell instance $86 m0 *1 0,117.39
X$86 86 133 134 dummy_cell_1rw
* cell instance $87 r0 *1 0,117.39
X$87 87 133 134 dummy_cell_1rw
* cell instance $88 m0 *1 0,120.12
X$88 88 133 134 dummy_cell_1rw
* cell instance $89 r0 *1 0,120.12
X$89 89 133 134 dummy_cell_1rw
* cell instance $90 m0 *1 0,122.85
X$90 90 133 134 dummy_cell_1rw
* cell instance $91 r0 *1 0,122.85
X$91 91 133 134 dummy_cell_1rw
* cell instance $92 m0 *1 0,125.58
X$92 92 133 134 dummy_cell_1rw
* cell instance $93 r0 *1 0,125.58
X$93 93 133 134 dummy_cell_1rw
* cell instance $94 m0 *1 0,128.31
X$94 94 133 134 dummy_cell_1rw
* cell instance $95 r0 *1 0,128.31
X$95 95 133 134 dummy_cell_1rw
* cell instance $96 m0 *1 0,131.04
X$96 96 133 134 dummy_cell_1rw
* cell instance $97 r0 *1 0,131.04
X$97 97 133 134 dummy_cell_1rw
* cell instance $98 m0 *1 0,133.77
X$98 98 133 134 dummy_cell_1rw
* cell instance $99 r0 *1 0,133.77
X$99 99 133 134 dummy_cell_1rw
* cell instance $100 m0 *1 0,136.5
X$100 100 133 134 dummy_cell_1rw
* cell instance $101 r0 *1 0,136.5
X$101 101 133 134 dummy_cell_1rw
* cell instance $102 m0 *1 0,139.23
X$102 102 133 134 dummy_cell_1rw
* cell instance $103 r0 *1 0,139.23
X$103 103 133 134 dummy_cell_1rw
* cell instance $104 m0 *1 0,141.96
X$104 104 133 134 dummy_cell_1rw
* cell instance $105 r0 *1 0,141.96
X$105 105 133 134 dummy_cell_1rw
* cell instance $106 m0 *1 0,144.69
X$106 106 133 134 dummy_cell_1rw
* cell instance $107 r0 *1 0,144.69
X$107 107 133 134 dummy_cell_1rw
* cell instance $108 m0 *1 0,147.42
X$108 108 133 134 dummy_cell_1rw
* cell instance $109 r0 *1 0,147.42
X$109 109 133 134 dummy_cell_1rw
* cell instance $110 m0 *1 0,150.15
X$110 110 133 134 dummy_cell_1rw
* cell instance $111 r0 *1 0,150.15
X$111 111 133 134 dummy_cell_1rw
* cell instance $112 m0 *1 0,152.88
X$112 112 133 134 dummy_cell_1rw
* cell instance $113 r0 *1 0,152.88
X$113 113 133 134 dummy_cell_1rw
* cell instance $114 m0 *1 0,155.61
X$114 114 133 134 dummy_cell_1rw
* cell instance $115 r0 *1 0,155.61
X$115 115 133 134 dummy_cell_1rw
* cell instance $116 m0 *1 0,158.34
X$116 116 133 134 dummy_cell_1rw
* cell instance $117 r0 *1 0,158.34
X$117 117 133 134 dummy_cell_1rw
* cell instance $118 m0 *1 0,161.07
X$118 118 133 134 dummy_cell_1rw
* cell instance $119 r0 *1 0,161.07
X$119 119 133 134 dummy_cell_1rw
* cell instance $120 m0 *1 0,163.8
X$120 120 133 134 dummy_cell_1rw
* cell instance $121 r0 *1 0,163.8
X$121 121 133 134 dummy_cell_1rw
* cell instance $122 m0 *1 0,166.53
X$122 122 133 134 dummy_cell_1rw
* cell instance $123 r0 *1 0,166.53
X$123 123 133 134 dummy_cell_1rw
* cell instance $124 m0 *1 0,169.26
X$124 124 133 134 dummy_cell_1rw
* cell instance $125 r0 *1 0,169.26
X$125 125 133 134 dummy_cell_1rw
* cell instance $126 m0 *1 0,171.99
X$126 126 133 134 dummy_cell_1rw
* cell instance $127 r0 *1 0,171.99
X$127 127 133 134 dummy_cell_1rw
* cell instance $128 m0 *1 0,174.72
X$128 128 133 134 dummy_cell_1rw
* cell instance $129 r0 *1 0,174.72
X$129 129 133 134 dummy_cell_1rw
* cell instance $130 m0 *1 0,177.45
X$130 130 133 134 dummy_cell_1rw
* cell instance $131 r0 *1 0,177.45
X$131 131 133 134 dummy_cell_1rw
* cell instance $132 m0 *1 0,180.18
X$132 132 133 134 dummy_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_2

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_0
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_0 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 1 2 3 dummy_cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 1 2 3 dummy_cell_1rw
* cell instance $4 r0 *1 2.115,0
X$4 1 2 3 dummy_cell_1rw
* cell instance $5 r0 *1 2.82,0
X$5 1 2 3 dummy_cell_1rw
* cell instance $6 r0 *1 3.525,0
X$6 1 2 3 dummy_cell_1rw
* cell instance $7 r0 *1 4.23,0
X$7 1 2 3 dummy_cell_1rw
* cell instance $8 r0 *1 4.935,0
X$8 1 2 3 dummy_cell_1rw
* cell instance $9 r0 *1 5.64,0
X$9 1 2 3 dummy_cell_1rw
* cell instance $10 r0 *1 6.345,0
X$10 1 2 3 dummy_cell_1rw
* cell instance $11 r0 *1 7.05,0
X$11 1 2 3 dummy_cell_1rw
* cell instance $12 r0 *1 7.755,0
X$12 1 2 3 dummy_cell_1rw
* cell instance $13 r0 *1 8.46,0
X$13 1 2 3 dummy_cell_1rw
* cell instance $14 r0 *1 9.165,0
X$14 1 2 3 dummy_cell_1rw
* cell instance $15 r0 *1 9.87,0
X$15 1 2 3 dummy_cell_1rw
* cell instance $16 r0 *1 10.575,0
X$16 1 2 3 dummy_cell_1rw
* cell instance $17 r0 *1 11.28,0
X$17 1 2 3 dummy_cell_1rw
* cell instance $18 r0 *1 11.985,0
X$18 1 2 3 dummy_cell_1rw
* cell instance $19 r0 *1 12.69,0
X$19 1 2 3 dummy_cell_1rw
* cell instance $20 r0 *1 13.395,0
X$20 1 2 3 dummy_cell_1rw
* cell instance $21 r0 *1 14.1,0
X$21 1 2 3 dummy_cell_1rw
* cell instance $22 r0 *1 14.805,0
X$22 1 2 3 dummy_cell_1rw
* cell instance $23 r0 *1 15.51,0
X$23 1 2 3 dummy_cell_1rw
* cell instance $24 r0 *1 16.215,0
X$24 1 2 3 dummy_cell_1rw
* cell instance $25 r0 *1 16.92,0
X$25 1 2 3 dummy_cell_1rw
* cell instance $26 r0 *1 17.625,0
X$26 1 2 3 dummy_cell_1rw
* cell instance $27 r0 *1 18.33,0
X$27 1 2 3 dummy_cell_1rw
* cell instance $28 r0 *1 19.035,0
X$28 1 2 3 dummy_cell_1rw
* cell instance $29 r0 *1 19.74,0
X$29 1 2 3 dummy_cell_1rw
* cell instance $30 r0 *1 20.445,0
X$30 1 2 3 dummy_cell_1rw
* cell instance $31 r0 *1 21.15,0
X$31 1 2 3 dummy_cell_1rw
* cell instance $32 r0 *1 21.855,0
X$32 1 2 3 dummy_cell_1rw
* cell instance $33 r0 *1 22.56,0
X$33 1 2 3 dummy_cell_1rw
* cell instance $34 r0 *1 23.265,0
X$34 1 2 3 dummy_cell_1rw
* cell instance $35 r0 *1 23.97,0
X$35 1 2 3 dummy_cell_1rw
* cell instance $36 r0 *1 24.675,0
X$36 1 2 3 dummy_cell_1rw
* cell instance $37 r0 *1 25.38,0
X$37 1 2 3 dummy_cell_1rw
* cell instance $38 r0 *1 26.085,0
X$38 1 2 3 dummy_cell_1rw
* cell instance $39 r0 *1 26.79,0
X$39 1 2 3 dummy_cell_1rw
* cell instance $40 r0 *1 27.495,0
X$40 1 2 3 dummy_cell_1rw
* cell instance $41 r0 *1 28.2,0
X$41 1 2 3 dummy_cell_1rw
* cell instance $42 r0 *1 28.905,0
X$42 1 2 3 dummy_cell_1rw
* cell instance $43 r0 *1 29.61,0
X$43 1 2 3 dummy_cell_1rw
* cell instance $44 r0 *1 30.315,0
X$44 1 2 3 dummy_cell_1rw
* cell instance $45 r0 *1 31.02,0
X$45 1 2 3 dummy_cell_1rw
* cell instance $46 r0 *1 31.725,0
X$46 1 2 3 dummy_cell_1rw
* cell instance $47 r0 *1 32.43,0
X$47 1 2 3 dummy_cell_1rw
* cell instance $48 r0 *1 33.135,0
X$48 1 2 3 dummy_cell_1rw
* cell instance $49 r0 *1 33.84,0
X$49 1 2 3 dummy_cell_1rw
* cell instance $50 r0 *1 34.545,0
X$50 1 2 3 dummy_cell_1rw
* cell instance $51 r0 *1 35.25,0
X$51 1 2 3 dummy_cell_1rw
* cell instance $52 r0 *1 35.955,0
X$52 1 2 3 dummy_cell_1rw
* cell instance $53 r0 *1 36.66,0
X$53 1 2 3 dummy_cell_1rw
* cell instance $54 r0 *1 37.365,0
X$54 1 2 3 dummy_cell_1rw
* cell instance $55 r0 *1 38.07,0
X$55 1 2 3 dummy_cell_1rw
* cell instance $56 r0 *1 38.775,0
X$56 1 2 3 dummy_cell_1rw
* cell instance $57 r0 *1 39.48,0
X$57 1 2 3 dummy_cell_1rw
* cell instance $58 r0 *1 40.185,0
X$58 1 2 3 dummy_cell_1rw
* cell instance $59 r0 *1 40.89,0
X$59 1 2 3 dummy_cell_1rw
* cell instance $60 r0 *1 41.595,0
X$60 1 2 3 dummy_cell_1rw
* cell instance $61 r0 *1 42.3,0
X$61 1 2 3 dummy_cell_1rw
* cell instance $62 r0 *1 43.005,0
X$62 1 2 3 dummy_cell_1rw
* cell instance $63 r0 *1 43.71,0
X$63 1 2 3 dummy_cell_1rw
* cell instance $64 r0 *1 44.415,0
X$64 1 2 3 dummy_cell_1rw
* cell instance $65 r0 *1 45.12,0
X$65 1 2 3 dummy_cell_1rw
* cell instance $66 r0 *1 45.825,0
X$66 1 2 3 dummy_cell_1rw
* cell instance $67 r0 *1 46.53,0
X$67 1 2 3 dummy_cell_1rw
* cell instance $68 r0 *1 47.235,0
X$68 1 2 3 dummy_cell_1rw
* cell instance $69 r0 *1 47.94,0
X$69 1 2 3 dummy_cell_1rw
* cell instance $70 r0 *1 48.645,0
X$70 1 2 3 dummy_cell_1rw
* cell instance $71 r0 *1 49.35,0
X$71 1 2 3 dummy_cell_1rw
* cell instance $72 r0 *1 50.055,0
X$72 1 2 3 dummy_cell_1rw
* cell instance $73 r0 *1 50.76,0
X$73 1 2 3 dummy_cell_1rw
* cell instance $74 r0 *1 51.465,0
X$74 1 2 3 dummy_cell_1rw
* cell instance $75 r0 *1 52.17,0
X$75 1 2 3 dummy_cell_1rw
* cell instance $76 r0 *1 52.875,0
X$76 1 2 3 dummy_cell_1rw
* cell instance $77 r0 *1 53.58,0
X$77 1 2 3 dummy_cell_1rw
* cell instance $78 r0 *1 54.285,0
X$78 1 2 3 dummy_cell_1rw
* cell instance $79 r0 *1 54.99,0
X$79 1 2 3 dummy_cell_1rw
* cell instance $80 r0 *1 55.695,0
X$80 1 2 3 dummy_cell_1rw
* cell instance $81 r0 *1 56.4,0
X$81 1 2 3 dummy_cell_1rw
* cell instance $82 r0 *1 57.105,0
X$82 1 2 3 dummy_cell_1rw
* cell instance $83 r0 *1 57.81,0
X$83 1 2 3 dummy_cell_1rw
* cell instance $84 r0 *1 58.515,0
X$84 1 2 3 dummy_cell_1rw
* cell instance $85 r0 *1 59.22,0
X$85 1 2 3 dummy_cell_1rw
* cell instance $86 r0 *1 59.925,0
X$86 1 2 3 dummy_cell_1rw
* cell instance $87 r0 *1 60.63,0
X$87 1 2 3 dummy_cell_1rw
* cell instance $88 r0 *1 61.335,0
X$88 1 2 3 dummy_cell_1rw
* cell instance $89 r0 *1 62.04,0
X$89 1 2 3 dummy_cell_1rw
* cell instance $90 r0 *1 62.745,0
X$90 1 2 3 dummy_cell_1rw
* cell instance $91 r0 *1 63.45,0
X$91 1 2 3 dummy_cell_1rw
* cell instance $92 r0 *1 64.155,0
X$92 1 2 3 dummy_cell_1rw
* cell instance $93 r0 *1 64.86,0
X$93 1 2 3 dummy_cell_1rw
* cell instance $94 r0 *1 65.565,0
X$94 1 2 3 dummy_cell_1rw
* cell instance $95 r0 *1 66.27,0
X$95 1 2 3 dummy_cell_1rw
* cell instance $96 r0 *1 66.975,0
X$96 1 2 3 dummy_cell_1rw
* cell instance $97 r0 *1 67.68,0
X$97 1 2 3 dummy_cell_1rw
* cell instance $98 r0 *1 68.385,0
X$98 1 2 3 dummy_cell_1rw
* cell instance $99 r0 *1 69.09,0
X$99 1 2 3 dummy_cell_1rw
* cell instance $100 r0 *1 69.795,0
X$100 1 2 3 dummy_cell_1rw
* cell instance $101 r0 *1 70.5,0
X$101 1 2 3 dummy_cell_1rw
* cell instance $102 r0 *1 71.205,0
X$102 1 2 3 dummy_cell_1rw
* cell instance $103 r0 *1 71.91,0
X$103 1 2 3 dummy_cell_1rw
* cell instance $104 r0 *1 72.615,0
X$104 1 2 3 dummy_cell_1rw
* cell instance $105 r0 *1 73.32,0
X$105 1 2 3 dummy_cell_1rw
* cell instance $106 r0 *1 74.025,0
X$106 1 2 3 dummy_cell_1rw
* cell instance $107 r0 *1 74.73,0
X$107 1 2 3 dummy_cell_1rw
* cell instance $108 r0 *1 75.435,0
X$108 1 2 3 dummy_cell_1rw
* cell instance $109 r0 *1 76.14,0
X$109 1 2 3 dummy_cell_1rw
* cell instance $110 r0 *1 76.845,0
X$110 1 2 3 dummy_cell_1rw
* cell instance $111 r0 *1 77.55,0
X$111 1 2 3 dummy_cell_1rw
* cell instance $112 r0 *1 78.255,0
X$112 1 2 3 dummy_cell_1rw
* cell instance $113 r0 *1 78.96,0
X$113 1 2 3 dummy_cell_1rw
* cell instance $114 r0 *1 79.665,0
X$114 1 2 3 dummy_cell_1rw
* cell instance $115 r0 *1 80.37,0
X$115 1 2 3 dummy_cell_1rw
* cell instance $116 r0 *1 81.075,0
X$116 1 2 3 dummy_cell_1rw
* cell instance $117 r0 *1 81.78,0
X$117 1 2 3 dummy_cell_1rw
* cell instance $118 r0 *1 82.485,0
X$118 1 2 3 dummy_cell_1rw
* cell instance $119 r0 *1 83.19,0
X$119 1 2 3 dummy_cell_1rw
* cell instance $120 r0 *1 83.895,0
X$120 1 2 3 dummy_cell_1rw
* cell instance $121 r0 *1 84.6,0
X$121 1 2 3 dummy_cell_1rw
* cell instance $122 r0 *1 85.305,0
X$122 1 2 3 dummy_cell_1rw
* cell instance $123 r0 *1 86.01,0
X$123 1 2 3 dummy_cell_1rw
* cell instance $124 r0 *1 86.715,0
X$124 1 2 3 dummy_cell_1rw
* cell instance $125 r0 *1 87.42,0
X$125 1 2 3 dummy_cell_1rw
* cell instance $126 r0 *1 88.125,0
X$126 1 2 3 dummy_cell_1rw
* cell instance $127 r0 *1 88.83,0
X$127 1 2 3 dummy_cell_1rw
* cell instance $128 r0 *1 89.535,0
X$128 1 2 3 dummy_cell_1rw
* cell instance $129 r0 *1 90.24,0
X$129 1 2 3 dummy_cell_1rw
* cell instance $130 r0 *1 90.945,0
X$130 1 2 3 dummy_cell_1rw
* cell instance $131 r0 *1 91.65,0
X$131 1 2 3 dummy_cell_1rw
* cell instance $132 r0 *1 92.355,0
X$132 1 2 3 dummy_cell_1rw
* cell instance $133 r0 *1 93.06,0
X$133 1 2 3 dummy_cell_1rw
* cell instance $134 r0 *1 93.765,0
X$134 1 2 3 dummy_cell_1rw
* cell instance $135 r0 *1 94.47,0
X$135 1 2 3 dummy_cell_1rw
* cell instance $136 r0 *1 95.175,0
X$136 1 2 3 dummy_cell_1rw
* cell instance $137 r0 *1 95.88,0
X$137 1 2 3 dummy_cell_1rw
* cell instance $138 r0 *1 96.585,0
X$138 1 2 3 dummy_cell_1rw
* cell instance $139 r0 *1 97.29,0
X$139 1 2 3 dummy_cell_1rw
* cell instance $140 r0 *1 97.995,0
X$140 1 2 3 dummy_cell_1rw
* cell instance $141 r0 *1 98.7,0
X$141 1 2 3 dummy_cell_1rw
* cell instance $142 r0 *1 99.405,0
X$142 1 2 3 dummy_cell_1rw
* cell instance $143 r0 *1 100.11,0
X$143 1 2 3 dummy_cell_1rw
* cell instance $144 r0 *1 100.815,0
X$144 1 2 3 dummy_cell_1rw
* cell instance $145 r0 *1 101.52,0
X$145 1 2 3 dummy_cell_1rw
* cell instance $146 r0 *1 102.225,0
X$146 1 2 3 dummy_cell_1rw
* cell instance $147 r0 *1 102.93,0
X$147 1 2 3 dummy_cell_1rw
* cell instance $148 r0 *1 103.635,0
X$148 1 2 3 dummy_cell_1rw
* cell instance $149 r0 *1 104.34,0
X$149 1 2 3 dummy_cell_1rw
* cell instance $150 r0 *1 105.045,0
X$150 1 2 3 dummy_cell_1rw
* cell instance $151 r0 *1 105.75,0
X$151 1 2 3 dummy_cell_1rw
* cell instance $152 r0 *1 106.455,0
X$152 1 2 3 dummy_cell_1rw
* cell instance $153 r0 *1 107.16,0
X$153 1 2 3 dummy_cell_1rw
* cell instance $154 r0 *1 107.865,0
X$154 1 2 3 dummy_cell_1rw
* cell instance $155 r0 *1 108.57,0
X$155 1 2 3 dummy_cell_1rw
* cell instance $156 r0 *1 109.275,0
X$156 1 2 3 dummy_cell_1rw
* cell instance $157 r0 *1 109.98,0
X$157 1 2 3 dummy_cell_1rw
* cell instance $158 r0 *1 110.685,0
X$158 1 2 3 dummy_cell_1rw
* cell instance $159 r0 *1 111.39,0
X$159 1 2 3 dummy_cell_1rw
* cell instance $160 r0 *1 112.095,0
X$160 1 2 3 dummy_cell_1rw
* cell instance $161 r0 *1 112.8,0
X$161 1 2 3 dummy_cell_1rw
* cell instance $162 r0 *1 113.505,0
X$162 1 2 3 dummy_cell_1rw
* cell instance $163 r0 *1 114.21,0
X$163 1 2 3 dummy_cell_1rw
* cell instance $164 r0 *1 114.915,0
X$164 1 2 3 dummy_cell_1rw
* cell instance $165 r0 *1 115.62,0
X$165 1 2 3 dummy_cell_1rw
* cell instance $166 r0 *1 116.325,0
X$166 1 2 3 dummy_cell_1rw
* cell instance $167 r0 *1 117.03,0
X$167 1 2 3 dummy_cell_1rw
* cell instance $168 r0 *1 117.735,0
X$168 1 2 3 dummy_cell_1rw
* cell instance $169 r0 *1 118.44,0
X$169 1 2 3 dummy_cell_1rw
* cell instance $170 r0 *1 119.145,0
X$170 1 2 3 dummy_cell_1rw
* cell instance $171 r0 *1 119.85,0
X$171 1 2 3 dummy_cell_1rw
* cell instance $172 r0 *1 120.555,0
X$172 1 2 3 dummy_cell_1rw
* cell instance $173 r0 *1 121.26,0
X$173 1 2 3 dummy_cell_1rw
* cell instance $174 r0 *1 121.965,0
X$174 1 2 3 dummy_cell_1rw
* cell instance $175 r0 *1 122.67,0
X$175 1 2 3 dummy_cell_1rw
* cell instance $176 r0 *1 123.375,0
X$176 1 2 3 dummy_cell_1rw
* cell instance $177 r0 *1 124.08,0
X$177 1 2 3 dummy_cell_1rw
* cell instance $178 r0 *1 124.785,0
X$178 1 2 3 dummy_cell_1rw
* cell instance $179 r0 *1 125.49,0
X$179 1 2 3 dummy_cell_1rw
* cell instance $180 r0 *1 126.195,0
X$180 1 2 3 dummy_cell_1rw
* cell instance $181 r0 *1 126.9,0
X$181 1 2 3 dummy_cell_1rw
* cell instance $182 r0 *1 127.605,0
X$182 1 2 3 dummy_cell_1rw
* cell instance $183 r0 *1 128.31,0
X$183 1 2 3 dummy_cell_1rw
* cell instance $184 r0 *1 129.015,0
X$184 1 2 3 dummy_cell_1rw
* cell instance $185 r0 *1 129.72,0
X$185 1 2 3 dummy_cell_1rw
* cell instance $186 r0 *1 130.425,0
X$186 1 2 3 dummy_cell_1rw
* cell instance $187 r0 *1 131.13,0
X$187 1 2 3 dummy_cell_1rw
* cell instance $188 r0 *1 131.835,0
X$188 1 2 3 dummy_cell_1rw
* cell instance $189 r0 *1 132.54,0
X$189 1 2 3 dummy_cell_1rw
* cell instance $190 r0 *1 133.245,0
X$190 1 2 3 dummy_cell_1rw
* cell instance $191 r0 *1 133.95,0
X$191 1 2 3 dummy_cell_1rw
* cell instance $192 r0 *1 134.655,0
X$192 1 2 3 dummy_cell_1rw
* cell instance $193 r0 *1 135.36,0
X$193 1 2 3 dummy_cell_1rw
* cell instance $194 r0 *1 136.065,0
X$194 1 2 3 dummy_cell_1rw
* cell instance $195 r0 *1 136.77,0
X$195 1 2 3 dummy_cell_1rw
* cell instance $196 r0 *1 137.475,0
X$196 1 2 3 dummy_cell_1rw
* cell instance $197 r0 *1 138.18,0
X$197 1 2 3 dummy_cell_1rw
* cell instance $198 r0 *1 138.885,0
X$198 1 2 3 dummy_cell_1rw
* cell instance $199 r0 *1 139.59,0
X$199 1 2 3 dummy_cell_1rw
* cell instance $200 r0 *1 140.295,0
X$200 1 2 3 dummy_cell_1rw
* cell instance $201 r0 *1 141,0
X$201 1 2 3 dummy_cell_1rw
* cell instance $202 r0 *1 141.705,0
X$202 1 2 3 dummy_cell_1rw
* cell instance $203 r0 *1 142.41,0
X$203 1 2 3 dummy_cell_1rw
* cell instance $204 r0 *1 143.115,0
X$204 1 2 3 dummy_cell_1rw
* cell instance $205 r0 *1 143.82,0
X$205 1 2 3 dummy_cell_1rw
* cell instance $206 r0 *1 144.525,0
X$206 1 2 3 dummy_cell_1rw
* cell instance $207 r0 *1 145.23,0
X$207 1 2 3 dummy_cell_1rw
* cell instance $208 r0 *1 145.935,0
X$208 1 2 3 dummy_cell_1rw
* cell instance $209 r0 *1 146.64,0
X$209 1 2 3 dummy_cell_1rw
* cell instance $210 r0 *1 147.345,0
X$210 1 2 3 dummy_cell_1rw
* cell instance $211 r0 *1 148.05,0
X$211 1 2 3 dummy_cell_1rw
* cell instance $212 r0 *1 148.755,0
X$212 1 2 3 dummy_cell_1rw
* cell instance $213 r0 *1 149.46,0
X$213 1 2 3 dummy_cell_1rw
* cell instance $214 r0 *1 150.165,0
X$214 1 2 3 dummy_cell_1rw
* cell instance $215 r0 *1 150.87,0
X$215 1 2 3 dummy_cell_1rw
* cell instance $216 r0 *1 151.575,0
X$216 1 2 3 dummy_cell_1rw
* cell instance $217 r0 *1 152.28,0
X$217 1 2 3 dummy_cell_1rw
* cell instance $218 r0 *1 152.985,0
X$218 1 2 3 dummy_cell_1rw
* cell instance $219 r0 *1 153.69,0
X$219 1 2 3 dummy_cell_1rw
* cell instance $220 r0 *1 154.395,0
X$220 1 2 3 dummy_cell_1rw
* cell instance $221 r0 *1 155.1,0
X$221 1 2 3 dummy_cell_1rw
* cell instance $222 r0 *1 155.805,0
X$222 1 2 3 dummy_cell_1rw
* cell instance $223 r0 *1 156.51,0
X$223 1 2 3 dummy_cell_1rw
* cell instance $224 r0 *1 157.215,0
X$224 1 2 3 dummy_cell_1rw
* cell instance $225 r0 *1 157.92,0
X$225 1 2 3 dummy_cell_1rw
* cell instance $226 r0 *1 158.625,0
X$226 1 2 3 dummy_cell_1rw
* cell instance $227 r0 *1 159.33,0
X$227 1 2 3 dummy_cell_1rw
* cell instance $228 r0 *1 160.035,0
X$228 1 2 3 dummy_cell_1rw
* cell instance $229 r0 *1 160.74,0
X$229 1 2 3 dummy_cell_1rw
* cell instance $230 r0 *1 161.445,0
X$230 1 2 3 dummy_cell_1rw
* cell instance $231 r0 *1 162.15,0
X$231 1 2 3 dummy_cell_1rw
* cell instance $232 r0 *1 162.855,0
X$232 1 2 3 dummy_cell_1rw
* cell instance $233 r0 *1 163.56,0
X$233 1 2 3 dummy_cell_1rw
* cell instance $234 r0 *1 164.265,0
X$234 1 2 3 dummy_cell_1rw
* cell instance $235 r0 *1 164.97,0
X$235 1 2 3 dummy_cell_1rw
* cell instance $236 r0 *1 165.675,0
X$236 1 2 3 dummy_cell_1rw
* cell instance $237 r0 *1 166.38,0
X$237 1 2 3 dummy_cell_1rw
* cell instance $238 r0 *1 167.085,0
X$238 1 2 3 dummy_cell_1rw
* cell instance $239 r0 *1 167.79,0
X$239 1 2 3 dummy_cell_1rw
* cell instance $240 r0 *1 168.495,0
X$240 1 2 3 dummy_cell_1rw
* cell instance $241 r0 *1 169.2,0
X$241 1 2 3 dummy_cell_1rw
* cell instance $242 r0 *1 169.905,0
X$242 1 2 3 dummy_cell_1rw
* cell instance $243 r0 *1 170.61,0
X$243 1 2 3 dummy_cell_1rw
* cell instance $244 r0 *1 171.315,0
X$244 1 2 3 dummy_cell_1rw
* cell instance $245 r0 *1 172.02,0
X$245 1 2 3 dummy_cell_1rw
* cell instance $246 r0 *1 172.725,0
X$246 1 2 3 dummy_cell_1rw
* cell instance $247 r0 *1 173.43,0
X$247 1 2 3 dummy_cell_1rw
* cell instance $248 r0 *1 174.135,0
X$248 1 2 3 dummy_cell_1rw
* cell instance $249 r0 *1 174.84,0
X$249 1 2 3 dummy_cell_1rw
* cell instance $250 r0 *1 175.545,0
X$250 1 2 3 dummy_cell_1rw
* cell instance $251 r0 *1 176.25,0
X$251 1 2 3 dummy_cell_1rw
* cell instance $252 r0 *1 176.955,0
X$252 1 2 3 dummy_cell_1rw
* cell instance $253 r0 *1 177.66,0
X$253 1 2 3 dummy_cell_1rw
* cell instance $254 r0 *1 178.365,0
X$254 1 2 3 dummy_cell_1rw
* cell instance $255 r0 *1 179.07,0
X$255 1 2 3 dummy_cell_1rw
* cell instance $256 r0 *1 179.775,0
X$256 1 2 3 dummy_cell_1rw
* cell instance $257 r0 *1 180.48,0
X$257 1 2 3 dummy_cell_1rw
* cell instance $258 r0 *1 181.185,0
X$258 1 2 3 dummy_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_1
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_1 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 1 2 3 dummy_cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 1 2 3 dummy_cell_1rw
* cell instance $4 r0 *1 2.115,0
X$4 1 2 3 dummy_cell_1rw
* cell instance $5 r0 *1 2.82,0
X$5 1 2 3 dummy_cell_1rw
* cell instance $6 r0 *1 3.525,0
X$6 1 2 3 dummy_cell_1rw
* cell instance $7 r0 *1 4.23,0
X$7 1 2 3 dummy_cell_1rw
* cell instance $8 r0 *1 4.935,0
X$8 1 2 3 dummy_cell_1rw
* cell instance $9 r0 *1 5.64,0
X$9 1 2 3 dummy_cell_1rw
* cell instance $10 r0 *1 6.345,0
X$10 1 2 3 dummy_cell_1rw
* cell instance $11 r0 *1 7.05,0
X$11 1 2 3 dummy_cell_1rw
* cell instance $12 r0 *1 7.755,0
X$12 1 2 3 dummy_cell_1rw
* cell instance $13 r0 *1 8.46,0
X$13 1 2 3 dummy_cell_1rw
* cell instance $14 r0 *1 9.165,0
X$14 1 2 3 dummy_cell_1rw
* cell instance $15 r0 *1 9.87,0
X$15 1 2 3 dummy_cell_1rw
* cell instance $16 r0 *1 10.575,0
X$16 1 2 3 dummy_cell_1rw
* cell instance $17 r0 *1 11.28,0
X$17 1 2 3 dummy_cell_1rw
* cell instance $18 r0 *1 11.985,0
X$18 1 2 3 dummy_cell_1rw
* cell instance $19 r0 *1 12.69,0
X$19 1 2 3 dummy_cell_1rw
* cell instance $20 r0 *1 13.395,0
X$20 1 2 3 dummy_cell_1rw
* cell instance $21 r0 *1 14.1,0
X$21 1 2 3 dummy_cell_1rw
* cell instance $22 r0 *1 14.805,0
X$22 1 2 3 dummy_cell_1rw
* cell instance $23 r0 *1 15.51,0
X$23 1 2 3 dummy_cell_1rw
* cell instance $24 r0 *1 16.215,0
X$24 1 2 3 dummy_cell_1rw
* cell instance $25 r0 *1 16.92,0
X$25 1 2 3 dummy_cell_1rw
* cell instance $26 r0 *1 17.625,0
X$26 1 2 3 dummy_cell_1rw
* cell instance $27 r0 *1 18.33,0
X$27 1 2 3 dummy_cell_1rw
* cell instance $28 r0 *1 19.035,0
X$28 1 2 3 dummy_cell_1rw
* cell instance $29 r0 *1 19.74,0
X$29 1 2 3 dummy_cell_1rw
* cell instance $30 r0 *1 20.445,0
X$30 1 2 3 dummy_cell_1rw
* cell instance $31 r0 *1 21.15,0
X$31 1 2 3 dummy_cell_1rw
* cell instance $32 r0 *1 21.855,0
X$32 1 2 3 dummy_cell_1rw
* cell instance $33 r0 *1 22.56,0
X$33 1 2 3 dummy_cell_1rw
* cell instance $34 r0 *1 23.265,0
X$34 1 2 3 dummy_cell_1rw
* cell instance $35 r0 *1 23.97,0
X$35 1 2 3 dummy_cell_1rw
* cell instance $36 r0 *1 24.675,0
X$36 1 2 3 dummy_cell_1rw
* cell instance $37 r0 *1 25.38,0
X$37 1 2 3 dummy_cell_1rw
* cell instance $38 r0 *1 26.085,0
X$38 1 2 3 dummy_cell_1rw
* cell instance $39 r0 *1 26.79,0
X$39 1 2 3 dummy_cell_1rw
* cell instance $40 r0 *1 27.495,0
X$40 1 2 3 dummy_cell_1rw
* cell instance $41 r0 *1 28.2,0
X$41 1 2 3 dummy_cell_1rw
* cell instance $42 r0 *1 28.905,0
X$42 1 2 3 dummy_cell_1rw
* cell instance $43 r0 *1 29.61,0
X$43 1 2 3 dummy_cell_1rw
* cell instance $44 r0 *1 30.315,0
X$44 1 2 3 dummy_cell_1rw
* cell instance $45 r0 *1 31.02,0
X$45 1 2 3 dummy_cell_1rw
* cell instance $46 r0 *1 31.725,0
X$46 1 2 3 dummy_cell_1rw
* cell instance $47 r0 *1 32.43,0
X$47 1 2 3 dummy_cell_1rw
* cell instance $48 r0 *1 33.135,0
X$48 1 2 3 dummy_cell_1rw
* cell instance $49 r0 *1 33.84,0
X$49 1 2 3 dummy_cell_1rw
* cell instance $50 r0 *1 34.545,0
X$50 1 2 3 dummy_cell_1rw
* cell instance $51 r0 *1 35.25,0
X$51 1 2 3 dummy_cell_1rw
* cell instance $52 r0 *1 35.955,0
X$52 1 2 3 dummy_cell_1rw
* cell instance $53 r0 *1 36.66,0
X$53 1 2 3 dummy_cell_1rw
* cell instance $54 r0 *1 37.365,0
X$54 1 2 3 dummy_cell_1rw
* cell instance $55 r0 *1 38.07,0
X$55 1 2 3 dummy_cell_1rw
* cell instance $56 r0 *1 38.775,0
X$56 1 2 3 dummy_cell_1rw
* cell instance $57 r0 *1 39.48,0
X$57 1 2 3 dummy_cell_1rw
* cell instance $58 r0 *1 40.185,0
X$58 1 2 3 dummy_cell_1rw
* cell instance $59 r0 *1 40.89,0
X$59 1 2 3 dummy_cell_1rw
* cell instance $60 r0 *1 41.595,0
X$60 1 2 3 dummy_cell_1rw
* cell instance $61 r0 *1 42.3,0
X$61 1 2 3 dummy_cell_1rw
* cell instance $62 r0 *1 43.005,0
X$62 1 2 3 dummy_cell_1rw
* cell instance $63 r0 *1 43.71,0
X$63 1 2 3 dummy_cell_1rw
* cell instance $64 r0 *1 44.415,0
X$64 1 2 3 dummy_cell_1rw
* cell instance $65 r0 *1 45.12,0
X$65 1 2 3 dummy_cell_1rw
* cell instance $66 r0 *1 45.825,0
X$66 1 2 3 dummy_cell_1rw
* cell instance $67 r0 *1 46.53,0
X$67 1 2 3 dummy_cell_1rw
* cell instance $68 r0 *1 47.235,0
X$68 1 2 3 dummy_cell_1rw
* cell instance $69 r0 *1 47.94,0
X$69 1 2 3 dummy_cell_1rw
* cell instance $70 r0 *1 48.645,0
X$70 1 2 3 dummy_cell_1rw
* cell instance $71 r0 *1 49.35,0
X$71 1 2 3 dummy_cell_1rw
* cell instance $72 r0 *1 50.055,0
X$72 1 2 3 dummy_cell_1rw
* cell instance $73 r0 *1 50.76,0
X$73 1 2 3 dummy_cell_1rw
* cell instance $74 r0 *1 51.465,0
X$74 1 2 3 dummy_cell_1rw
* cell instance $75 r0 *1 52.17,0
X$75 1 2 3 dummy_cell_1rw
* cell instance $76 r0 *1 52.875,0
X$76 1 2 3 dummy_cell_1rw
* cell instance $77 r0 *1 53.58,0
X$77 1 2 3 dummy_cell_1rw
* cell instance $78 r0 *1 54.285,0
X$78 1 2 3 dummy_cell_1rw
* cell instance $79 r0 *1 54.99,0
X$79 1 2 3 dummy_cell_1rw
* cell instance $80 r0 *1 55.695,0
X$80 1 2 3 dummy_cell_1rw
* cell instance $81 r0 *1 56.4,0
X$81 1 2 3 dummy_cell_1rw
* cell instance $82 r0 *1 57.105,0
X$82 1 2 3 dummy_cell_1rw
* cell instance $83 r0 *1 57.81,0
X$83 1 2 3 dummy_cell_1rw
* cell instance $84 r0 *1 58.515,0
X$84 1 2 3 dummy_cell_1rw
* cell instance $85 r0 *1 59.22,0
X$85 1 2 3 dummy_cell_1rw
* cell instance $86 r0 *1 59.925,0
X$86 1 2 3 dummy_cell_1rw
* cell instance $87 r0 *1 60.63,0
X$87 1 2 3 dummy_cell_1rw
* cell instance $88 r0 *1 61.335,0
X$88 1 2 3 dummy_cell_1rw
* cell instance $89 r0 *1 62.04,0
X$89 1 2 3 dummy_cell_1rw
* cell instance $90 r0 *1 62.745,0
X$90 1 2 3 dummy_cell_1rw
* cell instance $91 r0 *1 63.45,0
X$91 1 2 3 dummy_cell_1rw
* cell instance $92 r0 *1 64.155,0
X$92 1 2 3 dummy_cell_1rw
* cell instance $93 r0 *1 64.86,0
X$93 1 2 3 dummy_cell_1rw
* cell instance $94 r0 *1 65.565,0
X$94 1 2 3 dummy_cell_1rw
* cell instance $95 r0 *1 66.27,0
X$95 1 2 3 dummy_cell_1rw
* cell instance $96 r0 *1 66.975,0
X$96 1 2 3 dummy_cell_1rw
* cell instance $97 r0 *1 67.68,0
X$97 1 2 3 dummy_cell_1rw
* cell instance $98 r0 *1 68.385,0
X$98 1 2 3 dummy_cell_1rw
* cell instance $99 r0 *1 69.09,0
X$99 1 2 3 dummy_cell_1rw
* cell instance $100 r0 *1 69.795,0
X$100 1 2 3 dummy_cell_1rw
* cell instance $101 r0 *1 70.5,0
X$101 1 2 3 dummy_cell_1rw
* cell instance $102 r0 *1 71.205,0
X$102 1 2 3 dummy_cell_1rw
* cell instance $103 r0 *1 71.91,0
X$103 1 2 3 dummy_cell_1rw
* cell instance $104 r0 *1 72.615,0
X$104 1 2 3 dummy_cell_1rw
* cell instance $105 r0 *1 73.32,0
X$105 1 2 3 dummy_cell_1rw
* cell instance $106 r0 *1 74.025,0
X$106 1 2 3 dummy_cell_1rw
* cell instance $107 r0 *1 74.73,0
X$107 1 2 3 dummy_cell_1rw
* cell instance $108 r0 *1 75.435,0
X$108 1 2 3 dummy_cell_1rw
* cell instance $109 r0 *1 76.14,0
X$109 1 2 3 dummy_cell_1rw
* cell instance $110 r0 *1 76.845,0
X$110 1 2 3 dummy_cell_1rw
* cell instance $111 r0 *1 77.55,0
X$111 1 2 3 dummy_cell_1rw
* cell instance $112 r0 *1 78.255,0
X$112 1 2 3 dummy_cell_1rw
* cell instance $113 r0 *1 78.96,0
X$113 1 2 3 dummy_cell_1rw
* cell instance $114 r0 *1 79.665,0
X$114 1 2 3 dummy_cell_1rw
* cell instance $115 r0 *1 80.37,0
X$115 1 2 3 dummy_cell_1rw
* cell instance $116 r0 *1 81.075,0
X$116 1 2 3 dummy_cell_1rw
* cell instance $117 r0 *1 81.78,0
X$117 1 2 3 dummy_cell_1rw
* cell instance $118 r0 *1 82.485,0
X$118 1 2 3 dummy_cell_1rw
* cell instance $119 r0 *1 83.19,0
X$119 1 2 3 dummy_cell_1rw
* cell instance $120 r0 *1 83.895,0
X$120 1 2 3 dummy_cell_1rw
* cell instance $121 r0 *1 84.6,0
X$121 1 2 3 dummy_cell_1rw
* cell instance $122 r0 *1 85.305,0
X$122 1 2 3 dummy_cell_1rw
* cell instance $123 r0 *1 86.01,0
X$123 1 2 3 dummy_cell_1rw
* cell instance $124 r0 *1 86.715,0
X$124 1 2 3 dummy_cell_1rw
* cell instance $125 r0 *1 87.42,0
X$125 1 2 3 dummy_cell_1rw
* cell instance $126 r0 *1 88.125,0
X$126 1 2 3 dummy_cell_1rw
* cell instance $127 r0 *1 88.83,0
X$127 1 2 3 dummy_cell_1rw
* cell instance $128 r0 *1 89.535,0
X$128 1 2 3 dummy_cell_1rw
* cell instance $129 r0 *1 90.24,0
X$129 1 2 3 dummy_cell_1rw
* cell instance $130 r0 *1 90.945,0
X$130 1 2 3 dummy_cell_1rw
* cell instance $131 r0 *1 91.65,0
X$131 1 2 3 dummy_cell_1rw
* cell instance $132 r0 *1 92.355,0
X$132 1 2 3 dummy_cell_1rw
* cell instance $133 r0 *1 93.06,0
X$133 1 2 3 dummy_cell_1rw
* cell instance $134 r0 *1 93.765,0
X$134 1 2 3 dummy_cell_1rw
* cell instance $135 r0 *1 94.47,0
X$135 1 2 3 dummy_cell_1rw
* cell instance $136 r0 *1 95.175,0
X$136 1 2 3 dummy_cell_1rw
* cell instance $137 r0 *1 95.88,0
X$137 1 2 3 dummy_cell_1rw
* cell instance $138 r0 *1 96.585,0
X$138 1 2 3 dummy_cell_1rw
* cell instance $139 r0 *1 97.29,0
X$139 1 2 3 dummy_cell_1rw
* cell instance $140 r0 *1 97.995,0
X$140 1 2 3 dummy_cell_1rw
* cell instance $141 r0 *1 98.7,0
X$141 1 2 3 dummy_cell_1rw
* cell instance $142 r0 *1 99.405,0
X$142 1 2 3 dummy_cell_1rw
* cell instance $143 r0 *1 100.11,0
X$143 1 2 3 dummy_cell_1rw
* cell instance $144 r0 *1 100.815,0
X$144 1 2 3 dummy_cell_1rw
* cell instance $145 r0 *1 101.52,0
X$145 1 2 3 dummy_cell_1rw
* cell instance $146 r0 *1 102.225,0
X$146 1 2 3 dummy_cell_1rw
* cell instance $147 r0 *1 102.93,0
X$147 1 2 3 dummy_cell_1rw
* cell instance $148 r0 *1 103.635,0
X$148 1 2 3 dummy_cell_1rw
* cell instance $149 r0 *1 104.34,0
X$149 1 2 3 dummy_cell_1rw
* cell instance $150 r0 *1 105.045,0
X$150 1 2 3 dummy_cell_1rw
* cell instance $151 r0 *1 105.75,0
X$151 1 2 3 dummy_cell_1rw
* cell instance $152 r0 *1 106.455,0
X$152 1 2 3 dummy_cell_1rw
* cell instance $153 r0 *1 107.16,0
X$153 1 2 3 dummy_cell_1rw
* cell instance $154 r0 *1 107.865,0
X$154 1 2 3 dummy_cell_1rw
* cell instance $155 r0 *1 108.57,0
X$155 1 2 3 dummy_cell_1rw
* cell instance $156 r0 *1 109.275,0
X$156 1 2 3 dummy_cell_1rw
* cell instance $157 r0 *1 109.98,0
X$157 1 2 3 dummy_cell_1rw
* cell instance $158 r0 *1 110.685,0
X$158 1 2 3 dummy_cell_1rw
* cell instance $159 r0 *1 111.39,0
X$159 1 2 3 dummy_cell_1rw
* cell instance $160 r0 *1 112.095,0
X$160 1 2 3 dummy_cell_1rw
* cell instance $161 r0 *1 112.8,0
X$161 1 2 3 dummy_cell_1rw
* cell instance $162 r0 *1 113.505,0
X$162 1 2 3 dummy_cell_1rw
* cell instance $163 r0 *1 114.21,0
X$163 1 2 3 dummy_cell_1rw
* cell instance $164 r0 *1 114.915,0
X$164 1 2 3 dummy_cell_1rw
* cell instance $165 r0 *1 115.62,0
X$165 1 2 3 dummy_cell_1rw
* cell instance $166 r0 *1 116.325,0
X$166 1 2 3 dummy_cell_1rw
* cell instance $167 r0 *1 117.03,0
X$167 1 2 3 dummy_cell_1rw
* cell instance $168 r0 *1 117.735,0
X$168 1 2 3 dummy_cell_1rw
* cell instance $169 r0 *1 118.44,0
X$169 1 2 3 dummy_cell_1rw
* cell instance $170 r0 *1 119.145,0
X$170 1 2 3 dummy_cell_1rw
* cell instance $171 r0 *1 119.85,0
X$171 1 2 3 dummy_cell_1rw
* cell instance $172 r0 *1 120.555,0
X$172 1 2 3 dummy_cell_1rw
* cell instance $173 r0 *1 121.26,0
X$173 1 2 3 dummy_cell_1rw
* cell instance $174 r0 *1 121.965,0
X$174 1 2 3 dummy_cell_1rw
* cell instance $175 r0 *1 122.67,0
X$175 1 2 3 dummy_cell_1rw
* cell instance $176 r0 *1 123.375,0
X$176 1 2 3 dummy_cell_1rw
* cell instance $177 r0 *1 124.08,0
X$177 1 2 3 dummy_cell_1rw
* cell instance $178 r0 *1 124.785,0
X$178 1 2 3 dummy_cell_1rw
* cell instance $179 r0 *1 125.49,0
X$179 1 2 3 dummy_cell_1rw
* cell instance $180 r0 *1 126.195,0
X$180 1 2 3 dummy_cell_1rw
* cell instance $181 r0 *1 126.9,0
X$181 1 2 3 dummy_cell_1rw
* cell instance $182 r0 *1 127.605,0
X$182 1 2 3 dummy_cell_1rw
* cell instance $183 r0 *1 128.31,0
X$183 1 2 3 dummy_cell_1rw
* cell instance $184 r0 *1 129.015,0
X$184 1 2 3 dummy_cell_1rw
* cell instance $185 r0 *1 129.72,0
X$185 1 2 3 dummy_cell_1rw
* cell instance $186 r0 *1 130.425,0
X$186 1 2 3 dummy_cell_1rw
* cell instance $187 r0 *1 131.13,0
X$187 1 2 3 dummy_cell_1rw
* cell instance $188 r0 *1 131.835,0
X$188 1 2 3 dummy_cell_1rw
* cell instance $189 r0 *1 132.54,0
X$189 1 2 3 dummy_cell_1rw
* cell instance $190 r0 *1 133.245,0
X$190 1 2 3 dummy_cell_1rw
* cell instance $191 r0 *1 133.95,0
X$191 1 2 3 dummy_cell_1rw
* cell instance $192 r0 *1 134.655,0
X$192 1 2 3 dummy_cell_1rw
* cell instance $193 r0 *1 135.36,0
X$193 1 2 3 dummy_cell_1rw
* cell instance $194 r0 *1 136.065,0
X$194 1 2 3 dummy_cell_1rw
* cell instance $195 r0 *1 136.77,0
X$195 1 2 3 dummy_cell_1rw
* cell instance $196 r0 *1 137.475,0
X$196 1 2 3 dummy_cell_1rw
* cell instance $197 r0 *1 138.18,0
X$197 1 2 3 dummy_cell_1rw
* cell instance $198 r0 *1 138.885,0
X$198 1 2 3 dummy_cell_1rw
* cell instance $199 r0 *1 139.59,0
X$199 1 2 3 dummy_cell_1rw
* cell instance $200 r0 *1 140.295,0
X$200 1 2 3 dummy_cell_1rw
* cell instance $201 r0 *1 141,0
X$201 1 2 3 dummy_cell_1rw
* cell instance $202 r0 *1 141.705,0
X$202 1 2 3 dummy_cell_1rw
* cell instance $203 r0 *1 142.41,0
X$203 1 2 3 dummy_cell_1rw
* cell instance $204 r0 *1 143.115,0
X$204 1 2 3 dummy_cell_1rw
* cell instance $205 r0 *1 143.82,0
X$205 1 2 3 dummy_cell_1rw
* cell instance $206 r0 *1 144.525,0
X$206 1 2 3 dummy_cell_1rw
* cell instance $207 r0 *1 145.23,0
X$207 1 2 3 dummy_cell_1rw
* cell instance $208 r0 *1 145.935,0
X$208 1 2 3 dummy_cell_1rw
* cell instance $209 r0 *1 146.64,0
X$209 1 2 3 dummy_cell_1rw
* cell instance $210 r0 *1 147.345,0
X$210 1 2 3 dummy_cell_1rw
* cell instance $211 r0 *1 148.05,0
X$211 1 2 3 dummy_cell_1rw
* cell instance $212 r0 *1 148.755,0
X$212 1 2 3 dummy_cell_1rw
* cell instance $213 r0 *1 149.46,0
X$213 1 2 3 dummy_cell_1rw
* cell instance $214 r0 *1 150.165,0
X$214 1 2 3 dummy_cell_1rw
* cell instance $215 r0 *1 150.87,0
X$215 1 2 3 dummy_cell_1rw
* cell instance $216 r0 *1 151.575,0
X$216 1 2 3 dummy_cell_1rw
* cell instance $217 r0 *1 152.28,0
X$217 1 2 3 dummy_cell_1rw
* cell instance $218 r0 *1 152.985,0
X$218 1 2 3 dummy_cell_1rw
* cell instance $219 r0 *1 153.69,0
X$219 1 2 3 dummy_cell_1rw
* cell instance $220 r0 *1 154.395,0
X$220 1 2 3 dummy_cell_1rw
* cell instance $221 r0 *1 155.1,0
X$221 1 2 3 dummy_cell_1rw
* cell instance $222 r0 *1 155.805,0
X$222 1 2 3 dummy_cell_1rw
* cell instance $223 r0 *1 156.51,0
X$223 1 2 3 dummy_cell_1rw
* cell instance $224 r0 *1 157.215,0
X$224 1 2 3 dummy_cell_1rw
* cell instance $225 r0 *1 157.92,0
X$225 1 2 3 dummy_cell_1rw
* cell instance $226 r0 *1 158.625,0
X$226 1 2 3 dummy_cell_1rw
* cell instance $227 r0 *1 159.33,0
X$227 1 2 3 dummy_cell_1rw
* cell instance $228 r0 *1 160.035,0
X$228 1 2 3 dummy_cell_1rw
* cell instance $229 r0 *1 160.74,0
X$229 1 2 3 dummy_cell_1rw
* cell instance $230 r0 *1 161.445,0
X$230 1 2 3 dummy_cell_1rw
* cell instance $231 r0 *1 162.15,0
X$231 1 2 3 dummy_cell_1rw
* cell instance $232 r0 *1 162.855,0
X$232 1 2 3 dummy_cell_1rw
* cell instance $233 r0 *1 163.56,0
X$233 1 2 3 dummy_cell_1rw
* cell instance $234 r0 *1 164.265,0
X$234 1 2 3 dummy_cell_1rw
* cell instance $235 r0 *1 164.97,0
X$235 1 2 3 dummy_cell_1rw
* cell instance $236 r0 *1 165.675,0
X$236 1 2 3 dummy_cell_1rw
* cell instance $237 r0 *1 166.38,0
X$237 1 2 3 dummy_cell_1rw
* cell instance $238 r0 *1 167.085,0
X$238 1 2 3 dummy_cell_1rw
* cell instance $239 r0 *1 167.79,0
X$239 1 2 3 dummy_cell_1rw
* cell instance $240 r0 *1 168.495,0
X$240 1 2 3 dummy_cell_1rw
* cell instance $241 r0 *1 169.2,0
X$241 1 2 3 dummy_cell_1rw
* cell instance $242 r0 *1 169.905,0
X$242 1 2 3 dummy_cell_1rw
* cell instance $243 r0 *1 170.61,0
X$243 1 2 3 dummy_cell_1rw
* cell instance $244 r0 *1 171.315,0
X$244 1 2 3 dummy_cell_1rw
* cell instance $245 r0 *1 172.02,0
X$245 1 2 3 dummy_cell_1rw
* cell instance $246 r0 *1 172.725,0
X$246 1 2 3 dummy_cell_1rw
* cell instance $247 r0 *1 173.43,0
X$247 1 2 3 dummy_cell_1rw
* cell instance $248 r0 *1 174.135,0
X$248 1 2 3 dummy_cell_1rw
* cell instance $249 r0 *1 174.84,0
X$249 1 2 3 dummy_cell_1rw
* cell instance $250 r0 *1 175.545,0
X$250 1 2 3 dummy_cell_1rw
* cell instance $251 r0 *1 176.25,0
X$251 1 2 3 dummy_cell_1rw
* cell instance $252 r0 *1 176.955,0
X$252 1 2 3 dummy_cell_1rw
* cell instance $253 r0 *1 177.66,0
X$253 1 2 3 dummy_cell_1rw
* cell instance $254 r0 *1 178.365,0
X$254 1 2 3 dummy_cell_1rw
* cell instance $255 r0 *1 179.07,0
X$255 1 2 3 dummy_cell_1rw
* cell instance $256 r0 *1 179.775,0
X$256 1 2 3 dummy_cell_1rw
* cell instance $257 r0 *1 180.48,0
X$257 1 2 3 dummy_cell_1rw
* cell instance $258 r0 *1 181.185,0
X$258 1 2 3 dummy_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array_1

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_replica_bitcell_array
* pin rbl_wl_0_0
* pin rbl_bl_0_0
* pin rbl_br_0_0
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin bl_0_2
* pin br_0_2
* pin bl_0_3
* pin br_0_3
* pin bl_0_4
* pin br_0_4
* pin bl_0_5
* pin br_0_5
* pin bl_0_6
* pin br_0_6
* pin bl_0_7
* pin br_0_7
* pin bl_0_8
* pin br_0_8
* pin bl_0_9
* pin br_0_9
* pin bl_0_10
* pin br_0_10
* pin bl_0_11
* pin br_0_11
* pin bl_0_12
* pin br_0_12
* pin bl_0_13
* pin br_0_13
* pin bl_0_14
* pin br_0_14
* pin bl_0_15
* pin br_0_15
* pin bl_0_16
* pin br_0_16
* pin bl_0_17
* pin br_0_17
* pin bl_0_18
* pin br_0_18
* pin bl_0_19
* pin br_0_19
* pin bl_0_20
* pin br_0_20
* pin bl_0_21
* pin br_0_21
* pin bl_0_22
* pin br_0_22
* pin bl_0_23
* pin br_0_23
* pin bl_0_24
* pin br_0_24
* pin bl_0_25
* pin br_0_25
* pin bl_0_26
* pin br_0_26
* pin bl_0_27
* pin br_0_27
* pin bl_0_28
* pin br_0_28
* pin bl_0_29
* pin br_0_29
* pin bl_0_30
* pin br_0_30
* pin bl_0_31
* pin br_0_31
* pin bl_0_32
* pin br_0_32
* pin bl_0_33
* pin br_0_33
* pin bl_0_34
* pin br_0_34
* pin bl_0_35
* pin br_0_35
* pin bl_0_36
* pin br_0_36
* pin bl_0_37
* pin br_0_37
* pin bl_0_38
* pin br_0_38
* pin bl_0_39
* pin br_0_39
* pin bl_0_40
* pin br_0_40
* pin bl_0_41
* pin br_0_41
* pin bl_0_42
* pin br_0_42
* pin bl_0_43
* pin br_0_43
* pin bl_0_44
* pin br_0_44
* pin bl_0_45
* pin br_0_45
* pin bl_0_46
* pin br_0_46
* pin bl_0_47
* pin br_0_47
* pin bl_0_48
* pin br_0_48
* pin bl_0_49
* pin br_0_49
* pin bl_0_50
* pin br_0_50
* pin bl_0_51
* pin br_0_51
* pin bl_0_52
* pin br_0_52
* pin bl_0_53
* pin br_0_53
* pin bl_0_54
* pin br_0_54
* pin bl_0_55
* pin br_0_55
* pin bl_0_56
* pin br_0_56
* pin bl_0_57
* pin br_0_57
* pin bl_0_58
* pin br_0_58
* pin bl_0_59
* pin br_0_59
* pin bl_0_60
* pin br_0_60
* pin bl_0_61
* pin br_0_61
* pin bl_0_62
* pin br_0_62
* pin bl_0_63
* pin br_0_63
* pin bl_0_64
* pin br_0_64
* pin bl_0_65
* pin br_0_65
* pin bl_0_66
* pin br_0_66
* pin bl_0_67
* pin br_0_67
* pin bl_0_68
* pin br_0_68
* pin bl_0_69
* pin br_0_69
* pin bl_0_70
* pin br_0_70
* pin bl_0_71
* pin br_0_71
* pin bl_0_72
* pin br_0_72
* pin bl_0_73
* pin br_0_73
* pin bl_0_74
* pin br_0_74
* pin bl_0_75
* pin br_0_75
* pin bl_0_76
* pin br_0_76
* pin bl_0_77
* pin br_0_77
* pin bl_0_78
* pin br_0_78
* pin bl_0_79
* pin br_0_79
* pin bl_0_80
* pin br_0_80
* pin bl_0_81
* pin br_0_81
* pin bl_0_82
* pin br_0_82
* pin bl_0_83
* pin br_0_83
* pin bl_0_84
* pin br_0_84
* pin bl_0_85
* pin br_0_85
* pin bl_0_86
* pin br_0_86
* pin bl_0_87
* pin br_0_87
* pin bl_0_88
* pin br_0_88
* pin bl_0_89
* pin br_0_89
* pin bl_0_90
* pin br_0_90
* pin bl_0_91
* pin br_0_91
* pin bl_0_92
* pin br_0_92
* pin bl_0_93
* pin br_0_93
* pin bl_0_94
* pin br_0_94
* pin bl_0_95
* pin br_0_95
* pin bl_0_96
* pin br_0_96
* pin bl_0_97
* pin br_0_97
* pin bl_0_98
* pin br_0_98
* pin bl_0_99
* pin br_0_99
* pin bl_0_100
* pin br_0_100
* pin bl_0_101
* pin br_0_101
* pin bl_0_102
* pin br_0_102
* pin bl_0_103
* pin br_0_103
* pin bl_0_104
* pin br_0_104
* pin bl_0_105
* pin br_0_105
* pin bl_0_106
* pin br_0_106
* pin bl_0_107
* pin br_0_107
* pin bl_0_108
* pin br_0_108
* pin bl_0_109
* pin br_0_109
* pin bl_0_110
* pin br_0_110
* pin bl_0_111
* pin br_0_111
* pin bl_0_112
* pin br_0_112
* pin bl_0_113
* pin br_0_113
* pin bl_0_114
* pin br_0_114
* pin bl_0_115
* pin br_0_115
* pin bl_0_116
* pin br_0_116
* pin bl_0_117
* pin br_0_117
* pin bl_0_118
* pin br_0_118
* pin bl_0_119
* pin br_0_119
* pin bl_0_120
* pin br_0_120
* pin bl_0_121
* pin br_0_121
* pin bl_0_122
* pin br_0_122
* pin bl_0_123
* pin br_0_123
* pin bl_0_124
* pin br_0_124
* pin bl_0_125
* pin br_0_125
* pin bl_0_126
* pin br_0_126
* pin bl_0_127
* pin br_0_127
* pin bl_0_128
* pin br_0_128
* pin bl_0_129
* pin br_0_129
* pin bl_0_130
* pin br_0_130
* pin bl_0_131
* pin br_0_131
* pin bl_0_132
* pin br_0_132
* pin bl_0_133
* pin br_0_133
* pin bl_0_134
* pin br_0_134
* pin bl_0_135
* pin br_0_135
* pin bl_0_136
* pin br_0_136
* pin bl_0_137
* pin br_0_137
* pin bl_0_138
* pin br_0_138
* pin bl_0_139
* pin br_0_139
* pin bl_0_140
* pin br_0_140
* pin bl_0_141
* pin br_0_141
* pin bl_0_142
* pin br_0_142
* pin bl_0_143
* pin br_0_143
* pin bl_0_144
* pin br_0_144
* pin bl_0_145
* pin br_0_145
* pin bl_0_146
* pin br_0_146
* pin bl_0_147
* pin br_0_147
* pin bl_0_148
* pin br_0_148
* pin bl_0_149
* pin br_0_149
* pin bl_0_150
* pin br_0_150
* pin bl_0_151
* pin br_0_151
* pin bl_0_152
* pin br_0_152
* pin bl_0_153
* pin br_0_153
* pin bl_0_154
* pin br_0_154
* pin bl_0_155
* pin br_0_155
* pin bl_0_156
* pin br_0_156
* pin bl_0_157
* pin br_0_157
* pin bl_0_158
* pin br_0_158
* pin bl_0_159
* pin br_0_159
* pin bl_0_160
* pin br_0_160
* pin bl_0_161
* pin br_0_161
* pin bl_0_162
* pin br_0_162
* pin bl_0_163
* pin br_0_163
* pin bl_0_164
* pin br_0_164
* pin bl_0_165
* pin br_0_165
* pin bl_0_166
* pin br_0_166
* pin bl_0_167
* pin br_0_167
* pin bl_0_168
* pin br_0_168
* pin bl_0_169
* pin br_0_169
* pin bl_0_170
* pin br_0_170
* pin bl_0_171
* pin br_0_171
* pin bl_0_172
* pin br_0_172
* pin bl_0_173
* pin br_0_173
* pin bl_0_174
* pin br_0_174
* pin bl_0_175
* pin br_0_175
* pin bl_0_176
* pin br_0_176
* pin bl_0_177
* pin br_0_177
* pin bl_0_178
* pin br_0_178
* pin bl_0_179
* pin br_0_179
* pin bl_0_180
* pin br_0_180
* pin bl_0_181
* pin br_0_181
* pin bl_0_182
* pin br_0_182
* pin bl_0_183
* pin br_0_183
* pin bl_0_184
* pin br_0_184
* pin bl_0_185
* pin br_0_185
* pin bl_0_186
* pin br_0_186
* pin bl_0_187
* pin br_0_187
* pin bl_0_188
* pin br_0_188
* pin bl_0_189
* pin br_0_189
* pin bl_0_190
* pin br_0_190
* pin bl_0_191
* pin br_0_191
* pin bl_0_192
* pin br_0_192
* pin bl_0_193
* pin br_0_193
* pin bl_0_194
* pin br_0_194
* pin bl_0_195
* pin br_0_195
* pin bl_0_196
* pin br_0_196
* pin bl_0_197
* pin br_0_197
* pin bl_0_198
* pin br_0_198
* pin bl_0_199
* pin br_0_199
* pin bl_0_200
* pin br_0_200
* pin bl_0_201
* pin br_0_201
* pin bl_0_202
* pin br_0_202
* pin bl_0_203
* pin br_0_203
* pin bl_0_204
* pin br_0_204
* pin bl_0_205
* pin br_0_205
* pin bl_0_206
* pin br_0_206
* pin bl_0_207
* pin br_0_207
* pin bl_0_208
* pin br_0_208
* pin bl_0_209
* pin br_0_209
* pin bl_0_210
* pin br_0_210
* pin bl_0_211
* pin br_0_211
* pin bl_0_212
* pin br_0_212
* pin bl_0_213
* pin br_0_213
* pin bl_0_214
* pin br_0_214
* pin bl_0_215
* pin br_0_215
* pin bl_0_216
* pin br_0_216
* pin bl_0_217
* pin br_0_217
* pin bl_0_218
* pin br_0_218
* pin bl_0_219
* pin br_0_219
* pin bl_0_220
* pin br_0_220
* pin bl_0_221
* pin br_0_221
* pin bl_0_222
* pin br_0_222
* pin bl_0_223
* pin br_0_223
* pin bl_0_224
* pin br_0_224
* pin bl_0_225
* pin br_0_225
* pin bl_0_226
* pin br_0_226
* pin bl_0_227
* pin br_0_227
* pin bl_0_228
* pin br_0_228
* pin bl_0_229
* pin br_0_229
* pin bl_0_230
* pin br_0_230
* pin bl_0_231
* pin br_0_231
* pin bl_0_232
* pin br_0_232
* pin bl_0_233
* pin br_0_233
* pin bl_0_234
* pin br_0_234
* pin bl_0_235
* pin br_0_235
* pin bl_0_236
* pin br_0_236
* pin bl_0_237
* pin br_0_237
* pin bl_0_238
* pin br_0_238
* pin bl_0_239
* pin br_0_239
* pin bl_0_240
* pin br_0_240
* pin bl_0_241
* pin br_0_241
* pin bl_0_242
* pin br_0_242
* pin bl_0_243
* pin br_0_243
* pin bl_0_244
* pin br_0_244
* pin bl_0_245
* pin br_0_245
* pin bl_0_246
* pin br_0_246
* pin bl_0_247
* pin br_0_247
* pin bl_0_248
* pin br_0_248
* pin bl_0_249
* pin br_0_249
* pin bl_0_250
* pin br_0_250
* pin bl_0_251
* pin br_0_251
* pin bl_0_252
* pin br_0_252
* pin bl_0_253
* pin br_0_253
* pin bl_0_254
* pin br_0_254
* pin bl_0_255
* pin br_0_255
* pin bl_0_256
* pin br_0_256
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_24
* pin wl_0_25
* pin wl_0_26
* pin wl_0_27
* pin wl_0_28
* pin wl_0_29
* pin wl_0_30
* pin wl_0_31
* pin wl_0_32
* pin wl_0_33
* pin wl_0_34
* pin wl_0_35
* pin wl_0_36
* pin wl_0_37
* pin wl_0_38
* pin wl_0_39
* pin wl_0_40
* pin wl_0_41
* pin wl_0_42
* pin wl_0_43
* pin wl_0_44
* pin wl_0_45
* pin wl_0_46
* pin wl_0_47
* pin wl_0_48
* pin wl_0_49
* pin wl_0_50
* pin wl_0_51
* pin wl_0_52
* pin wl_0_53
* pin wl_0_54
* pin wl_0_55
* pin wl_0_56
* pin wl_0_57
* pin wl_0_58
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_62
* pin wl_0_63
* pin wl_0_64
* pin wl_0_65
* pin wl_0_66
* pin wl_0_67
* pin wl_0_68
* pin wl_0_69
* pin wl_0_70
* pin wl_0_71
* pin wl_0_72
* pin wl_0_73
* pin wl_0_74
* pin wl_0_75
* pin wl_0_76
* pin wl_0_77
* pin wl_0_78
* pin wl_0_79
* pin wl_0_80
* pin wl_0_81
* pin wl_0_82
* pin wl_0_83
* pin wl_0_84
* pin wl_0_85
* pin wl_0_86
* pin wl_0_87
* pin wl_0_88
* pin wl_0_89
* pin wl_0_90
* pin wl_0_91
* pin wl_0_92
* pin wl_0_93
* pin wl_0_94
* pin wl_0_95
* pin wl_0_96
* pin wl_0_97
* pin wl_0_98
* pin wl_0_99
* pin wl_0_100
* pin wl_0_101
* pin wl_0_102
* pin wl_0_103
* pin wl_0_104
* pin wl_0_105
* pin wl_0_106
* pin wl_0_107
* pin wl_0_108
* pin wl_0_109
* pin wl_0_110
* pin wl_0_111
* pin wl_0_112
* pin wl_0_113
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_117
* pin wl_0_118
* pin wl_0_119
* pin wl_0_120
* pin wl_0_121
* pin wl_0_122
* pin wl_0_123
* pin wl_0_124
* pin wl_0_125
* pin wl_0_126
* pin wl_0_127
* pin wl_0_128
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_replica_bitcell_array 1 2 3 4 5 6
+ 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33
+ 34 35 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59
+ 60 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85
+ 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108
+ 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127
+ 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146
+ 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165
+ 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279
+ 280 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298
+ 299 300 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317
+ 318 319 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336
+ 337 338 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355
+ 356 357 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374
+ 375 376 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393
+ 394 395 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412
+ 413 414 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431
+ 432 433 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450
+ 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469
+ 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488
+ 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507
+ 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526
+ 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545
+ 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564
+ 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583
+ 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621
+ 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640
+ 641 642 643 644 645 646 647 648
* net 1 rbl_wl_0_0
* net 2 rbl_bl_0_0
* net 3 rbl_br_0_0
* net 4 bl_0_0
* net 5 br_0_0
* net 6 bl_0_1
* net 7 br_0_1
* net 8 bl_0_2
* net 9 br_0_2
* net 10 bl_0_3
* net 11 br_0_3
* net 12 bl_0_4
* net 13 br_0_4
* net 14 bl_0_5
* net 15 br_0_5
* net 16 bl_0_6
* net 17 br_0_6
* net 18 bl_0_7
* net 19 br_0_7
* net 20 bl_0_8
* net 21 br_0_8
* net 22 bl_0_9
* net 23 br_0_9
* net 24 bl_0_10
* net 25 br_0_10
* net 26 bl_0_11
* net 27 br_0_11
* net 28 bl_0_12
* net 29 br_0_12
* net 30 bl_0_13
* net 31 br_0_13
* net 32 bl_0_14
* net 33 br_0_14
* net 34 bl_0_15
* net 35 br_0_15
* net 36 bl_0_16
* net 37 br_0_16
* net 38 bl_0_17
* net 39 br_0_17
* net 40 bl_0_18
* net 41 br_0_18
* net 42 bl_0_19
* net 43 br_0_19
* net 44 bl_0_20
* net 45 br_0_20
* net 46 bl_0_21
* net 47 br_0_21
* net 48 bl_0_22
* net 49 br_0_22
* net 50 bl_0_23
* net 51 br_0_23
* net 52 bl_0_24
* net 53 br_0_24
* net 54 bl_0_25
* net 55 br_0_25
* net 56 bl_0_26
* net 57 br_0_26
* net 58 bl_0_27
* net 59 br_0_27
* net 60 bl_0_28
* net 61 br_0_28
* net 62 bl_0_29
* net 63 br_0_29
* net 64 bl_0_30
* net 65 br_0_30
* net 66 bl_0_31
* net 67 br_0_31
* net 68 bl_0_32
* net 69 br_0_32
* net 70 bl_0_33
* net 71 br_0_33
* net 72 bl_0_34
* net 73 br_0_34
* net 74 bl_0_35
* net 75 br_0_35
* net 76 bl_0_36
* net 77 br_0_36
* net 78 bl_0_37
* net 79 br_0_37
* net 80 bl_0_38
* net 81 br_0_38
* net 82 bl_0_39
* net 83 br_0_39
* net 84 bl_0_40
* net 85 br_0_40
* net 86 bl_0_41
* net 87 br_0_41
* net 88 bl_0_42
* net 89 br_0_42
* net 90 bl_0_43
* net 91 br_0_43
* net 92 bl_0_44
* net 93 br_0_44
* net 94 bl_0_45
* net 95 br_0_45
* net 96 bl_0_46
* net 97 br_0_46
* net 98 bl_0_47
* net 99 br_0_47
* net 100 bl_0_48
* net 101 br_0_48
* net 102 bl_0_49
* net 103 br_0_49
* net 104 bl_0_50
* net 105 br_0_50
* net 106 bl_0_51
* net 107 br_0_51
* net 108 bl_0_52
* net 109 br_0_52
* net 110 bl_0_53
* net 111 br_0_53
* net 112 bl_0_54
* net 113 br_0_54
* net 114 bl_0_55
* net 115 br_0_55
* net 116 bl_0_56
* net 117 br_0_56
* net 118 bl_0_57
* net 119 br_0_57
* net 120 bl_0_58
* net 121 br_0_58
* net 122 bl_0_59
* net 123 br_0_59
* net 124 bl_0_60
* net 125 br_0_60
* net 126 bl_0_61
* net 127 br_0_61
* net 128 bl_0_62
* net 129 br_0_62
* net 130 bl_0_63
* net 131 br_0_63
* net 132 bl_0_64
* net 133 br_0_64
* net 134 bl_0_65
* net 135 br_0_65
* net 136 bl_0_66
* net 137 br_0_66
* net 138 bl_0_67
* net 139 br_0_67
* net 140 bl_0_68
* net 141 br_0_68
* net 142 bl_0_69
* net 143 br_0_69
* net 144 bl_0_70
* net 145 br_0_70
* net 146 bl_0_71
* net 147 br_0_71
* net 148 bl_0_72
* net 149 br_0_72
* net 150 bl_0_73
* net 151 br_0_73
* net 152 bl_0_74
* net 153 br_0_74
* net 154 bl_0_75
* net 155 br_0_75
* net 156 bl_0_76
* net 157 br_0_76
* net 158 bl_0_77
* net 159 br_0_77
* net 160 bl_0_78
* net 161 br_0_78
* net 162 bl_0_79
* net 163 br_0_79
* net 164 bl_0_80
* net 165 br_0_80
* net 166 bl_0_81
* net 167 br_0_81
* net 168 bl_0_82
* net 169 br_0_82
* net 170 bl_0_83
* net 171 br_0_83
* net 172 bl_0_84
* net 173 br_0_84
* net 174 bl_0_85
* net 175 br_0_85
* net 176 bl_0_86
* net 177 br_0_86
* net 178 bl_0_87
* net 179 br_0_87
* net 180 bl_0_88
* net 181 br_0_88
* net 182 bl_0_89
* net 183 br_0_89
* net 184 bl_0_90
* net 185 br_0_90
* net 186 bl_0_91
* net 187 br_0_91
* net 188 bl_0_92
* net 189 br_0_92
* net 190 bl_0_93
* net 191 br_0_93
* net 192 bl_0_94
* net 193 br_0_94
* net 194 bl_0_95
* net 195 br_0_95
* net 196 bl_0_96
* net 197 br_0_96
* net 198 bl_0_97
* net 199 br_0_97
* net 200 bl_0_98
* net 201 br_0_98
* net 202 bl_0_99
* net 203 br_0_99
* net 204 bl_0_100
* net 205 br_0_100
* net 206 bl_0_101
* net 207 br_0_101
* net 208 bl_0_102
* net 209 br_0_102
* net 210 bl_0_103
* net 211 br_0_103
* net 212 bl_0_104
* net 213 br_0_104
* net 214 bl_0_105
* net 215 br_0_105
* net 216 bl_0_106
* net 217 br_0_106
* net 218 bl_0_107
* net 219 br_0_107
* net 220 bl_0_108
* net 221 br_0_108
* net 222 bl_0_109
* net 223 br_0_109
* net 224 bl_0_110
* net 225 br_0_110
* net 226 bl_0_111
* net 227 br_0_111
* net 228 bl_0_112
* net 229 br_0_112
* net 230 bl_0_113
* net 231 br_0_113
* net 232 bl_0_114
* net 233 br_0_114
* net 234 bl_0_115
* net 235 br_0_115
* net 236 bl_0_116
* net 237 br_0_116
* net 238 bl_0_117
* net 239 br_0_117
* net 240 bl_0_118
* net 241 br_0_118
* net 242 bl_0_119
* net 243 br_0_119
* net 244 bl_0_120
* net 245 br_0_120
* net 246 bl_0_121
* net 247 br_0_121
* net 248 bl_0_122
* net 249 br_0_122
* net 250 bl_0_123
* net 251 br_0_123
* net 252 bl_0_124
* net 253 br_0_124
* net 254 bl_0_125
* net 255 br_0_125
* net 256 bl_0_126
* net 257 br_0_126
* net 258 bl_0_127
* net 259 br_0_127
* net 260 bl_0_128
* net 261 br_0_128
* net 262 bl_0_129
* net 263 br_0_129
* net 264 bl_0_130
* net 265 br_0_130
* net 266 bl_0_131
* net 267 br_0_131
* net 268 bl_0_132
* net 269 br_0_132
* net 270 bl_0_133
* net 271 br_0_133
* net 272 bl_0_134
* net 273 br_0_134
* net 274 bl_0_135
* net 275 br_0_135
* net 276 bl_0_136
* net 277 br_0_136
* net 278 bl_0_137
* net 279 br_0_137
* net 280 bl_0_138
* net 281 br_0_138
* net 282 bl_0_139
* net 283 br_0_139
* net 284 bl_0_140
* net 285 br_0_140
* net 286 bl_0_141
* net 287 br_0_141
* net 288 bl_0_142
* net 289 br_0_142
* net 290 bl_0_143
* net 291 br_0_143
* net 292 bl_0_144
* net 293 br_0_144
* net 294 bl_0_145
* net 295 br_0_145
* net 296 bl_0_146
* net 297 br_0_146
* net 298 bl_0_147
* net 299 br_0_147
* net 300 bl_0_148
* net 301 br_0_148
* net 302 bl_0_149
* net 303 br_0_149
* net 304 bl_0_150
* net 305 br_0_150
* net 306 bl_0_151
* net 307 br_0_151
* net 308 bl_0_152
* net 309 br_0_152
* net 310 bl_0_153
* net 311 br_0_153
* net 312 bl_0_154
* net 313 br_0_154
* net 314 bl_0_155
* net 315 br_0_155
* net 316 bl_0_156
* net 317 br_0_156
* net 318 bl_0_157
* net 319 br_0_157
* net 320 bl_0_158
* net 321 br_0_158
* net 322 bl_0_159
* net 323 br_0_159
* net 324 bl_0_160
* net 325 br_0_160
* net 326 bl_0_161
* net 327 br_0_161
* net 328 bl_0_162
* net 329 br_0_162
* net 330 bl_0_163
* net 331 br_0_163
* net 332 bl_0_164
* net 333 br_0_164
* net 334 bl_0_165
* net 335 br_0_165
* net 336 bl_0_166
* net 337 br_0_166
* net 338 bl_0_167
* net 339 br_0_167
* net 340 bl_0_168
* net 341 br_0_168
* net 342 bl_0_169
* net 343 br_0_169
* net 344 bl_0_170
* net 345 br_0_170
* net 346 bl_0_171
* net 347 br_0_171
* net 348 bl_0_172
* net 349 br_0_172
* net 350 bl_0_173
* net 351 br_0_173
* net 352 bl_0_174
* net 353 br_0_174
* net 354 bl_0_175
* net 355 br_0_175
* net 356 bl_0_176
* net 357 br_0_176
* net 358 bl_0_177
* net 359 br_0_177
* net 360 bl_0_178
* net 361 br_0_178
* net 362 bl_0_179
* net 363 br_0_179
* net 364 bl_0_180
* net 365 br_0_180
* net 366 bl_0_181
* net 367 br_0_181
* net 368 bl_0_182
* net 369 br_0_182
* net 370 bl_0_183
* net 371 br_0_183
* net 372 bl_0_184
* net 373 br_0_184
* net 374 bl_0_185
* net 375 br_0_185
* net 376 bl_0_186
* net 377 br_0_186
* net 378 bl_0_187
* net 379 br_0_187
* net 380 bl_0_188
* net 381 br_0_188
* net 382 bl_0_189
* net 383 br_0_189
* net 384 bl_0_190
* net 385 br_0_190
* net 386 bl_0_191
* net 387 br_0_191
* net 388 bl_0_192
* net 389 br_0_192
* net 390 bl_0_193
* net 391 br_0_193
* net 392 bl_0_194
* net 393 br_0_194
* net 394 bl_0_195
* net 395 br_0_195
* net 396 bl_0_196
* net 397 br_0_196
* net 398 bl_0_197
* net 399 br_0_197
* net 400 bl_0_198
* net 401 br_0_198
* net 402 bl_0_199
* net 403 br_0_199
* net 404 bl_0_200
* net 405 br_0_200
* net 406 bl_0_201
* net 407 br_0_201
* net 408 bl_0_202
* net 409 br_0_202
* net 410 bl_0_203
* net 411 br_0_203
* net 412 bl_0_204
* net 413 br_0_204
* net 414 bl_0_205
* net 415 br_0_205
* net 416 bl_0_206
* net 417 br_0_206
* net 418 bl_0_207
* net 419 br_0_207
* net 420 bl_0_208
* net 421 br_0_208
* net 422 bl_0_209
* net 423 br_0_209
* net 424 bl_0_210
* net 425 br_0_210
* net 426 bl_0_211
* net 427 br_0_211
* net 428 bl_0_212
* net 429 br_0_212
* net 430 bl_0_213
* net 431 br_0_213
* net 432 bl_0_214
* net 433 br_0_214
* net 434 bl_0_215
* net 435 br_0_215
* net 436 bl_0_216
* net 437 br_0_216
* net 438 bl_0_217
* net 439 br_0_217
* net 440 bl_0_218
* net 441 br_0_218
* net 442 bl_0_219
* net 443 br_0_219
* net 444 bl_0_220
* net 445 br_0_220
* net 446 bl_0_221
* net 447 br_0_221
* net 448 bl_0_222
* net 449 br_0_222
* net 450 bl_0_223
* net 451 br_0_223
* net 452 bl_0_224
* net 453 br_0_224
* net 454 bl_0_225
* net 455 br_0_225
* net 456 bl_0_226
* net 457 br_0_226
* net 458 bl_0_227
* net 459 br_0_227
* net 460 bl_0_228
* net 461 br_0_228
* net 462 bl_0_229
* net 463 br_0_229
* net 464 bl_0_230
* net 465 br_0_230
* net 466 bl_0_231
* net 467 br_0_231
* net 468 bl_0_232
* net 469 br_0_232
* net 470 bl_0_233
* net 471 br_0_233
* net 472 bl_0_234
* net 473 br_0_234
* net 474 bl_0_235
* net 475 br_0_235
* net 476 bl_0_236
* net 477 br_0_236
* net 478 bl_0_237
* net 479 br_0_237
* net 480 bl_0_238
* net 481 br_0_238
* net 482 bl_0_239
* net 483 br_0_239
* net 484 bl_0_240
* net 485 br_0_240
* net 486 bl_0_241
* net 487 br_0_241
* net 488 bl_0_242
* net 489 br_0_242
* net 490 bl_0_243
* net 491 br_0_243
* net 492 bl_0_244
* net 493 br_0_244
* net 494 bl_0_245
* net 495 br_0_245
* net 496 bl_0_246
* net 497 br_0_246
* net 498 bl_0_247
* net 499 br_0_247
* net 500 bl_0_248
* net 501 br_0_248
* net 502 bl_0_249
* net 503 br_0_249
* net 504 bl_0_250
* net 505 br_0_250
* net 506 bl_0_251
* net 507 br_0_251
* net 508 bl_0_252
* net 509 br_0_252
* net 510 bl_0_253
* net 511 br_0_253
* net 512 bl_0_254
* net 513 br_0_254
* net 514 bl_0_255
* net 515 br_0_255
* net 516 bl_0_256
* net 517 br_0_256
* net 518 wl_0_0
* net 519 wl_0_1
* net 520 wl_0_2
* net 521 wl_0_3
* net 522 wl_0_4
* net 523 wl_0_5
* net 524 wl_0_6
* net 525 wl_0_7
* net 526 wl_0_8
* net 527 wl_0_9
* net 528 wl_0_10
* net 529 wl_0_11
* net 530 wl_0_12
* net 531 wl_0_13
* net 532 wl_0_14
* net 533 wl_0_15
* net 534 wl_0_16
* net 535 wl_0_17
* net 536 wl_0_18
* net 537 wl_0_19
* net 538 wl_0_20
* net 539 wl_0_21
* net 540 wl_0_22
* net 541 wl_0_23
* net 542 wl_0_24
* net 543 wl_0_25
* net 544 wl_0_26
* net 545 wl_0_27
* net 546 wl_0_28
* net 547 wl_0_29
* net 548 wl_0_30
* net 549 wl_0_31
* net 550 wl_0_32
* net 551 wl_0_33
* net 552 wl_0_34
* net 553 wl_0_35
* net 554 wl_0_36
* net 555 wl_0_37
* net 556 wl_0_38
* net 557 wl_0_39
* net 558 wl_0_40
* net 559 wl_0_41
* net 560 wl_0_42
* net 561 wl_0_43
* net 562 wl_0_44
* net 563 wl_0_45
* net 564 wl_0_46
* net 565 wl_0_47
* net 566 wl_0_48
* net 567 wl_0_49
* net 568 wl_0_50
* net 569 wl_0_51
* net 570 wl_0_52
* net 571 wl_0_53
* net 572 wl_0_54
* net 573 wl_0_55
* net 574 wl_0_56
* net 575 wl_0_57
* net 576 wl_0_58
* net 577 wl_0_59
* net 578 wl_0_60
* net 579 wl_0_61
* net 580 wl_0_62
* net 581 wl_0_63
* net 582 wl_0_64
* net 583 wl_0_65
* net 584 wl_0_66
* net 585 wl_0_67
* net 586 wl_0_68
* net 587 wl_0_69
* net 588 wl_0_70
* net 589 wl_0_71
* net 590 wl_0_72
* net 591 wl_0_73
* net 592 wl_0_74
* net 593 wl_0_75
* net 594 wl_0_76
* net 595 wl_0_77
* net 596 wl_0_78
* net 597 wl_0_79
* net 598 wl_0_80
* net 599 wl_0_81
* net 600 wl_0_82
* net 601 wl_0_83
* net 602 wl_0_84
* net 603 wl_0_85
* net 604 wl_0_86
* net 605 wl_0_87
* net 606 wl_0_88
* net 607 wl_0_89
* net 608 wl_0_90
* net 609 wl_0_91
* net 610 wl_0_92
* net 611 wl_0_93
* net 612 wl_0_94
* net 613 wl_0_95
* net 614 wl_0_96
* net 615 wl_0_97
* net 616 wl_0_98
* net 617 wl_0_99
* net 618 wl_0_100
* net 619 wl_0_101
* net 620 wl_0_102
* net 621 wl_0_103
* net 622 wl_0_104
* net 623 wl_0_105
* net 624 wl_0_106
* net 625 wl_0_107
* net 626 wl_0_108
* net 627 wl_0_109
* net 628 wl_0_110
* net 629 wl_0_111
* net 630 wl_0_112
* net 631 wl_0_113
* net 632 wl_0_114
* net 633 wl_0_115
* net 634 wl_0_116
* net 635 wl_0_117
* net 636 wl_0_118
* net 637 wl_0_119
* net 638 wl_0_120
* net 639 wl_0_121
* net 640 wl_0_122
* net 641 wl_0_123
* net 642 wl_0_124
* net 643 wl_0_125
* net 644 wl_0_126
* net 645 wl_0_127
* net 646 wl_0_128
* net 647 vdd
* net 648 gnd
* cell instance $1 r0 *1 0,0
X$1 1 518 519 520 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535
+ 536 537 538 539 540 541 542 543 544 545 546 547 548 549 550 551 552 553 554
+ 555 556 557 558 559 560 561 562 563 564 565 566 567 568 569 570 571 572 573
+ 574 575 576 577 578 579 580 2 581 3 582 583 584 585 586 587 588 589 590 591
+ 592 593 594 595 596 597 598 599 600 601 602 603 604 605 606 607 608 609 610
+ 611 612 613 614 615 616 617 618 619 620 621 622 623 624 625 626 627 628 629
+ 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644 645 646 647 648
+ freepdk45_sram_4kbytes_1rw_32x1024_8_replica_column
* cell instance $2 m0 *1 0.705,1.365
X$2 1 647 648 freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array
* cell instance $3 r0 *1 0.705,1.365
X$3 518 519 521 520 522 523 524 525 527 526 528 529 530 531 532 533 534 535 536
+ 537 538 539 540 541 543 542 544 545 546 547 548 549 550 551 552 553 554 555
+ 557 556 559 558 561 560 562 563 564 565 566 567 568 569 570 571 572 573 574
+ 575 576 577 578 579 580 581 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44 45 46 47
+ 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66 67 68 69 70 71 72 73
+ 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99
+ 100 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118
+ 119 120 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137
+ 138 139 140 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156
+ 157 158 159 160 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175
+ 176 177 178 179 180 181 182 183 184 185 186 187 188 189 190 191 192 193 194
+ 195 196 197 198 199 200 201 202 203 204 205 206 207 208 209 210 211 212 213
+ 214 215 216 217 218 219 220 221 222 223 224 225 226 227 228 229 230 231 232
+ 233 234 235 236 237 238 239 240 241 242 243 244 245 246 247 248 249 250 251
+ 252 253 254 255 256 257 258 259 260 582 261 262 263 264 265 266 267 268 269
+ 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284 285 286 287 288
+ 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304 305 306 307
+ 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324 325 326
+ 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344 345
+ 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364
+ 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383
+ 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459
+ 460 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478
+ 479 480 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497
+ 498 499 500 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516
+ 517 584 583 586 585 587 588 589 590 591 592 593 594 596 595 597 598 600 599
+ 601 602 603 604 605 606 607 608 609 610 612 611 613 614 615 616 618 617 620
+ 619 621 622 623 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638
+ 640 639 642 641 643 644 645 646 647 648
+ freepdk45_sram_4kbytes_1rw_32x1024_8_bitcell_array
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_replica_bitcell_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_5
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_5 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.36U AS=0.0432P AD=0.0432P PS=1.02U PD=1.02U
* device instance $3 r0 *1 0.2325,2.075 PMOS_VTG
M$3 3 1 2 3 PMOS_VTG L=0.05U W=1.08U AS=0.1296P AD=0.1296P PS=2.1U PD=2.1U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_5

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_4
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_4 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,2.075 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_4

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_6
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_6 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.26 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=1.08U AS=0.12555P AD=0.12555P PS=2.28U PD=2.28U
* device instance $5 r0 *1 0.2325,1.94 PMOS_VTG
M$5 3 1 2 3 PMOS_VTG L=0.05U W=3.24U AS=0.37665P AD=0.37665P PS=4.98U PD=4.98U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_6

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_16
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_16 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.2735 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=2.975U AS=0.33915P AD=0.33915P PS=5.5525U
+ PD=5.5525U
* device instance $11 r0 *1 0.2325,1.9 PMOS_VTG
M$11 3 1 2 3 PMOS_VTG L=0.05U W=8.9U AS=1.0146P AD=1.0146P PS=12.07U PD=12.07U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_16

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_15
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_15 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.275 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=3.6U AS=0.4095P AD=0.4095P PS=6.63U PD=6.63U
* device instance $13 r0 *1 0.2325,1.895 PMOS_VTG
M$13 3 1 2 3 PMOS_VTG L=0.05U W=10.8U AS=1.2285P AD=1.2285P PS=14.43U PD=14.43U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_15

* cell dff
* pin Q
* pin D
* pin clk
* pin vdd
* pin gnd
.SUBCKT dff 2 5 7 16 17
* net 2 Q
* net 5 D
* net 7 clk
* net 16 vdd
* net 17 gnd
* device instance $1 r0 *1 0.2925,1.5425 PMOS_VTG
M$1 16 5 13 16 PMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.035P PS=1.21U PD=0.64U
* device instance $2 r0 *1 0.4825,1.5425 PMOS_VTG
M$2 13 7 4 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $3 r0 *1 0.6725,1.5425 PMOS_VTG
M$3 4 1 14 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.035P PS=0.64U PD=0.64U
* device instance $4 r0 *1 0.8625,1.5425 PMOS_VTG
M$4 14 6 16 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.0851P PS=0.64U PD=1.275U
* device instance $5 r0 *1 1.1575,1.5425 PMOS_VTG
M$5 16 4 6 16 PMOS_VTG L=0.05U W=0.5U AS=0.0851P AD=0.0525P PS=1.275U PD=1.21U
* device instance $6 r0 *1 2.2325,1.4525 PMOS_VTG
M$6 8 7 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.038125P AD=0.0375P PS=0.7U PD=0.8U
* device instance $7 r0 *1 1.7925,1.5775 PMOS_VTG
M$7 16 6 15 16 PMOS_VTG L=0.05U W=0.5U AS=0.0875P AD=0.035P PS=1.245U PD=0.64U
* device instance $8 r0 *1 1.9825,1.5775 PMOS_VTG
M$8 15 1 8 16 PMOS_VTG L=0.05U W=0.5U AS=0.035P AD=0.038125P PS=0.64U PD=0.7U
* device instance $9 r0 *1 1.4975,1.65 PMOS_VTG
M$9 1 7 16 16 PMOS_VTG L=0.05U W=1U AS=0.105P AD=0.0875P PS=2.21U PD=1.245U
* device instance $10 r0 *1 2.3225,2.0175 PMOS_VTG
M$10 16 2 12 16 PMOS_VTG L=0.05U W=0.25U AS=0.055125P AD=0.02625P PS=1.21U
+ PD=0.71U
* device instance $11 r0 *1 2.5825,1.7925 PMOS_VTG
M$11 16 8 2 16 PMOS_VTG L=0.05U W=1U AS=0.055125P AD=0.105P PS=1.21U PD=2.21U
* device instance $12 r0 *1 2.0475,0.3475 NMOS_VTG
M$12 17 2 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.02625P PS=0.71U
+ PD=0.71U
* device instance $13 r0 *1 2.5825,0.7125 NMOS_VTG
M$13 17 8 2 17 NMOS_VTG L=0.05U W=0.5U AS=0.0775P AD=0.0525P PS=1.31U PD=1.21U
* device instance $14 r0 *1 0.2925,0.725 NMOS_VTG
M$14 17 5 9 17 NMOS_VTG L=0.05U W=0.25U AS=0.02625P AD=0.0175P PS=0.71U PD=0.39U
* device instance $15 r0 *1 0.4825,0.725 NMOS_VTG
M$15 9 1 4 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $16 r0 *1 0.6725,0.725 NMOS_VTG
M$16 4 7 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $17 r0 *1 0.8625,0.725 NMOS_VTG
M$17 17 6 10 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.0175P PS=0.93U PD=0.39U
* device instance $18 r0 *1 1.1575,0.725 NMOS_VTG
M$18 17 4 6 17 NMOS_VTG L=0.05U W=0.25U AS=0.0502P AD=0.02625P PS=0.93U PD=0.71U
* device instance $19 r0 *1 1.4975,0.6575 NMOS_VTG
M$19 1 7 17 17 NMOS_VTG L=0.05U W=0.5U AS=0.0525P AD=0.04375P PS=1.21U PD=0.745U
* device instance $20 r0 *1 1.7925,0.7825 NMOS_VTG
M$20 17 6 11 17 NMOS_VTG L=0.05U W=0.25U AS=0.04375P AD=0.0175P PS=0.745U
+ PD=0.39U
* device instance $21 r0 *1 1.9825,0.7825 NMOS_VTG
M$21 11 7 8 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0175P PS=0.39U PD=0.39U
* device instance $22 r0 *1 2.1725,0.7825 NMOS_VTG
M$22 8 1 3 17 NMOS_VTG L=0.05U W=0.25U AS=0.0175P AD=0.0275P PS=0.39U PD=0.72U
.ENDS dff

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pand3
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pand3 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 5 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0
* cell instance $2 r0 *1 0.965,0
X$2 2 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_0
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pand3

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_3

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0.9025,0
X$1 1 2 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_0
* cell instance $2 r0 *1 0,0
X$2 3 4 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_wordline_driver

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode2x4
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin out_2
* pin out_3
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode2x4 1 2 5 6
+ 7 8 9 10
* net 1 in_0
* net 2 in_1
* net 5 out_0
* net 6 out_1
* net 7 out_2
* net 8 out_3
* net 9 vdd
* net 10 gnd
* cell instance $1 m0 *1 2.0875,2.73
X$1 6 1 4 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec
* cell instance $2 m0 *1 2.0875,5.46
X$2 8 1 2 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec
* cell instance $8 r0 *1 0.56,0
X$8 1 3 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
* cell instance $9 r0 *1 2.0875,2.73
X$9 7 3 2 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec
* cell instance $15 m0 *1 0.56,2.73
X$15 2 4 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
* cell instance $16 r0 *1 2.0875,0
X$16 5 3 4 9 10 freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode2x4

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8
* pin in_0
* pin in_1
* pin out_0
* pin out_1
* pin in_2
* pin out_2
* pin out_3
* pin out_4
* pin out_5
* pin out_6
* pin out_7
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8 1 4 6 7
+ 8 9 10 11 12 13 14 15 16
* net 1 in_0
* net 4 in_1
* net 6 out_0
* net 7 out_1
* net 8 in_2
* net 9 out_2
* net 10 out_3
* net 11 out_4
* net 12 out_5
* net 13 out_6
* net 14 out_7
* net 15 vdd
* net 16 gnd
* cell instance $1 m0 *1 2.5075,2.73
X$1 7 1 3 5 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $2 m0 *1 2.5075,10.92
X$2 14 1 4 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $3 m0 *1 2.5075,5.46
X$3 10 1 4 5 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $4 m0 *1 2.5075,8.19
X$4 12 1 3 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $12 r0 *1 0.7,0
X$12 1 2 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
* cell instance $13 r0 *1 2.5075,0
X$13 6 2 3 5 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $14 r0 *1 2.5075,5.46
X$14 11 2 3 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $15 r0 *1 2.5075,2.73
X$15 9 2 4 5 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $16 r0 *1 2.5075,8.19
X$16 13 2 4 8 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* cell instance $27 m0 *1 0.7,2.73
X$27 4 3 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
* cell instance $40 r0 *1 0.7,2.73
X$40 8 5 15 16 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_hierarchical_predecode3x8

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux
* pin sel
* pin bl
* pin br_out
* pin bl_out
* pin br
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux 1 2 3 4 5 6
* net 1 sel
* net 2 bl
* net 3 br_out
* net 4 bl_out
* net 5 br
* net 6 gnd
* device instance $1 r0 *1 0.3525,0.44 NMOS_VTG
M$1 3 1 5 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
* device instance $2 r0 *1 0.3525,1.3 NMOS_VTG
M$2 4 1 2 6 NMOS_VTG L=0.05U W=0.72U AS=0.0918P AD=0.0918P PS=1.695U PD=1.695U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_column_mux

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pand2
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pand2 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_0
* cell instance $2 r0 *1 0.75,0
X$2 2 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pand2

* cell write_driver
* pin din
* pin en
* pin br
* pin bl
* pin vdd
* pin gnd
.SUBCKT write_driver 1 2 5 9 11 12
* net 1 din
* net 2 en
* net 5 br
* net 9 bl
* net 11 vdd
* net 12 gnd
* device instance $1 r0 *1 0.17,3.0725 PMOS_VTG
M$1 11 3 8 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $2 r0 *1 0.36,3.0725 PMOS_VTG
M$2 8 4 9 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $3 r0 *1 0.17,2.46 PMOS_VTG
M$3 11 1 7 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0252P PS=0.93U PD=0.5U
* device instance $4 r0 *1 0.36,2.46 PMOS_VTG
M$4 7 4 5 11 PMOS_VTG L=0.05U W=0.36U AS=0.0252P AD=0.0378P PS=0.5U PD=0.93U
* device instance $5 r0 *1 0.51,0.885 PMOS_VTG
M$5 4 2 11 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $6 r0 *1 0.17,0.885 PMOS_VTG
M$6 11 1 3 11 PMOS_VTG L=0.05U W=0.36U AS=0.0378P AD=0.0378P PS=0.93U PD=0.93U
* device instance $7 r0 *1 0.17,3.6775 NMOS_VTG
M$7 12 3 10 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $8 r0 *1 0.36,3.6775 NMOS_VTG
M$8 10 2 9 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $9 r0 *1 0.17,1.855 NMOS_VTG
M$9 12 1 6 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0126P PS=0.57U PD=0.32U
* device instance $10 r0 *1 0.36,1.855 NMOS_VTG
M$10 6 2 5 12 NMOS_VTG L=0.05U W=0.18U AS=0.0126P AD=0.0189P PS=0.32U PD=0.57U
* device instance $11 r0 *1 0.51,1.49 NMOS_VTG
M$11 4 2 12 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
* device instance $12 r0 *1 0.17,1.49 NMOS_VTG
M$12 12 1 3 12 NMOS_VTG L=0.05U W=0.18U AS=0.0189P AD=0.0189P PS=0.57U PD=0.57U
.ENDS write_driver

* cell sense_amp
* pin br
* pin bl
* pin dout
* pin en
* pin vdd
* pin gnd
.SUBCKT sense_amp 1 2 3 4 7 8
* net 1 br
* net 2 bl
* net 3 dout
* net 4 en
* net 7 vdd
* net 8 gnd
* device instance $1 r0 *1 0.2575,2.9725 PMOS_VTG
M$1 3 5 7 7 PMOS_VTG L=0.05U W=0.54U AS=0.0567P AD=0.0378P PS=1.29U PD=0.68U
* device instance $2 r0 *1 0.4475,2.9725 PMOS_VTG
M$2 7 3 5 7 PMOS_VTG L=0.05U W=0.54U AS=0.0378P AD=0.0567P PS=0.68U PD=1.29U
* device instance $3 r0 *1 0.4475,2.025 PMOS_VTG
M$3 5 4 1 7 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $4 r0 *1 0.2575,1.055 PMOS_VTG
M$4 2 4 3 7 PMOS_VTG L=0.05U W=0.72U AS=0.0756P AD=0.0756P PS=1.65U PD=1.65U
* device instance $5 r0 *1 0.3575,4.32 NMOS_VTG
M$5 6 4 8 8 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.02835P PS=0.75U PD=0.75U
* device instance $6 r0 *1 0.2575,3.8625 NMOS_VTG
M$6 3 5 6 8 NMOS_VTG L=0.05U W=0.27U AS=0.02835P AD=0.0189P PS=0.75U PD=0.41U
* device instance $7 r0 *1 0.4475,3.8625 NMOS_VTG
M$7 6 3 5 8 NMOS_VTG L=0.05U W=0.27U AS=0.0189P AD=0.02835P PS=0.41U PD=0.75U
.ENDS sense_amp

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0
* pin en_bar
* pin bl
* pin br
* pin vdd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0 1 2 3 4
* net 1 en_bar
* net 2 bl
* net 3 br
* net 4 vdd
* device instance $1 r0 *1 0.265,0.905 PMOS_VTG
M$1 2 1 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.48,0.905 PMOS_VTG
M$2 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.265,0.355 PMOS_VTG
M$3 2 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_precharge_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array
* pin wl_0_0
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array 1 2 3
* net 1 wl_0_0
* net 2 vdd
* net 3 gnd
* cell instance $1 r0 *1 0,0
X$1 1 2 3 dummy_cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 1 2 3 dummy_cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 1 2 3 dummy_cell_1rw
* cell instance $4 r0 *1 2.115,0
X$4 1 2 3 dummy_cell_1rw
* cell instance $5 r0 *1 2.82,0
X$5 1 2 3 dummy_cell_1rw
* cell instance $6 r0 *1 3.525,0
X$6 1 2 3 dummy_cell_1rw
* cell instance $7 r0 *1 4.23,0
X$7 1 2 3 dummy_cell_1rw
* cell instance $8 r0 *1 4.935,0
X$8 1 2 3 dummy_cell_1rw
* cell instance $9 r0 *1 5.64,0
X$9 1 2 3 dummy_cell_1rw
* cell instance $10 r0 *1 6.345,0
X$10 1 2 3 dummy_cell_1rw
* cell instance $11 r0 *1 7.05,0
X$11 1 2 3 dummy_cell_1rw
* cell instance $12 r0 *1 7.755,0
X$12 1 2 3 dummy_cell_1rw
* cell instance $13 r0 *1 8.46,0
X$13 1 2 3 dummy_cell_1rw
* cell instance $14 r0 *1 9.165,0
X$14 1 2 3 dummy_cell_1rw
* cell instance $15 r0 *1 9.87,0
X$15 1 2 3 dummy_cell_1rw
* cell instance $16 r0 *1 10.575,0
X$16 1 2 3 dummy_cell_1rw
* cell instance $17 r0 *1 11.28,0
X$17 1 2 3 dummy_cell_1rw
* cell instance $18 r0 *1 11.985,0
X$18 1 2 3 dummy_cell_1rw
* cell instance $19 r0 *1 12.69,0
X$19 1 2 3 dummy_cell_1rw
* cell instance $20 r0 *1 13.395,0
X$20 1 2 3 dummy_cell_1rw
* cell instance $21 r0 *1 14.1,0
X$21 1 2 3 dummy_cell_1rw
* cell instance $22 r0 *1 14.805,0
X$22 1 2 3 dummy_cell_1rw
* cell instance $23 r0 *1 15.51,0
X$23 1 2 3 dummy_cell_1rw
* cell instance $24 r0 *1 16.215,0
X$24 1 2 3 dummy_cell_1rw
* cell instance $25 r0 *1 16.92,0
X$25 1 2 3 dummy_cell_1rw
* cell instance $26 r0 *1 17.625,0
X$26 1 2 3 dummy_cell_1rw
* cell instance $27 r0 *1 18.33,0
X$27 1 2 3 dummy_cell_1rw
* cell instance $28 r0 *1 19.035,0
X$28 1 2 3 dummy_cell_1rw
* cell instance $29 r0 *1 19.74,0
X$29 1 2 3 dummy_cell_1rw
* cell instance $30 r0 *1 20.445,0
X$30 1 2 3 dummy_cell_1rw
* cell instance $31 r0 *1 21.15,0
X$31 1 2 3 dummy_cell_1rw
* cell instance $32 r0 *1 21.855,0
X$32 1 2 3 dummy_cell_1rw
* cell instance $33 r0 *1 22.56,0
X$33 1 2 3 dummy_cell_1rw
* cell instance $34 r0 *1 23.265,0
X$34 1 2 3 dummy_cell_1rw
* cell instance $35 r0 *1 23.97,0
X$35 1 2 3 dummy_cell_1rw
* cell instance $36 r0 *1 24.675,0
X$36 1 2 3 dummy_cell_1rw
* cell instance $37 r0 *1 25.38,0
X$37 1 2 3 dummy_cell_1rw
* cell instance $38 r0 *1 26.085,0
X$38 1 2 3 dummy_cell_1rw
* cell instance $39 r0 *1 26.79,0
X$39 1 2 3 dummy_cell_1rw
* cell instance $40 r0 *1 27.495,0
X$40 1 2 3 dummy_cell_1rw
* cell instance $41 r0 *1 28.2,0
X$41 1 2 3 dummy_cell_1rw
* cell instance $42 r0 *1 28.905,0
X$42 1 2 3 dummy_cell_1rw
* cell instance $43 r0 *1 29.61,0
X$43 1 2 3 dummy_cell_1rw
* cell instance $44 r0 *1 30.315,0
X$44 1 2 3 dummy_cell_1rw
* cell instance $45 r0 *1 31.02,0
X$45 1 2 3 dummy_cell_1rw
* cell instance $46 r0 *1 31.725,0
X$46 1 2 3 dummy_cell_1rw
* cell instance $47 r0 *1 32.43,0
X$47 1 2 3 dummy_cell_1rw
* cell instance $48 r0 *1 33.135,0
X$48 1 2 3 dummy_cell_1rw
* cell instance $49 r0 *1 33.84,0
X$49 1 2 3 dummy_cell_1rw
* cell instance $50 r0 *1 34.545,0
X$50 1 2 3 dummy_cell_1rw
* cell instance $51 r0 *1 35.25,0
X$51 1 2 3 dummy_cell_1rw
* cell instance $52 r0 *1 35.955,0
X$52 1 2 3 dummy_cell_1rw
* cell instance $53 r0 *1 36.66,0
X$53 1 2 3 dummy_cell_1rw
* cell instance $54 r0 *1 37.365,0
X$54 1 2 3 dummy_cell_1rw
* cell instance $55 r0 *1 38.07,0
X$55 1 2 3 dummy_cell_1rw
* cell instance $56 r0 *1 38.775,0
X$56 1 2 3 dummy_cell_1rw
* cell instance $57 r0 *1 39.48,0
X$57 1 2 3 dummy_cell_1rw
* cell instance $58 r0 *1 40.185,0
X$58 1 2 3 dummy_cell_1rw
* cell instance $59 r0 *1 40.89,0
X$59 1 2 3 dummy_cell_1rw
* cell instance $60 r0 *1 41.595,0
X$60 1 2 3 dummy_cell_1rw
* cell instance $61 r0 *1 42.3,0
X$61 1 2 3 dummy_cell_1rw
* cell instance $62 r0 *1 43.005,0
X$62 1 2 3 dummy_cell_1rw
* cell instance $63 r0 *1 43.71,0
X$63 1 2 3 dummy_cell_1rw
* cell instance $64 r0 *1 44.415,0
X$64 1 2 3 dummy_cell_1rw
* cell instance $65 r0 *1 45.12,0
X$65 1 2 3 dummy_cell_1rw
* cell instance $66 r0 *1 45.825,0
X$66 1 2 3 dummy_cell_1rw
* cell instance $67 r0 *1 46.53,0
X$67 1 2 3 dummy_cell_1rw
* cell instance $68 r0 *1 47.235,0
X$68 1 2 3 dummy_cell_1rw
* cell instance $69 r0 *1 47.94,0
X$69 1 2 3 dummy_cell_1rw
* cell instance $70 r0 *1 48.645,0
X$70 1 2 3 dummy_cell_1rw
* cell instance $71 r0 *1 49.35,0
X$71 1 2 3 dummy_cell_1rw
* cell instance $72 r0 *1 50.055,0
X$72 1 2 3 dummy_cell_1rw
* cell instance $73 r0 *1 50.76,0
X$73 1 2 3 dummy_cell_1rw
* cell instance $74 r0 *1 51.465,0
X$74 1 2 3 dummy_cell_1rw
* cell instance $75 r0 *1 52.17,0
X$75 1 2 3 dummy_cell_1rw
* cell instance $76 r0 *1 52.875,0
X$76 1 2 3 dummy_cell_1rw
* cell instance $77 r0 *1 53.58,0
X$77 1 2 3 dummy_cell_1rw
* cell instance $78 r0 *1 54.285,0
X$78 1 2 3 dummy_cell_1rw
* cell instance $79 r0 *1 54.99,0
X$79 1 2 3 dummy_cell_1rw
* cell instance $80 r0 *1 55.695,0
X$80 1 2 3 dummy_cell_1rw
* cell instance $81 r0 *1 56.4,0
X$81 1 2 3 dummy_cell_1rw
* cell instance $82 r0 *1 57.105,0
X$82 1 2 3 dummy_cell_1rw
* cell instance $83 r0 *1 57.81,0
X$83 1 2 3 dummy_cell_1rw
* cell instance $84 r0 *1 58.515,0
X$84 1 2 3 dummy_cell_1rw
* cell instance $85 r0 *1 59.22,0
X$85 1 2 3 dummy_cell_1rw
* cell instance $86 r0 *1 59.925,0
X$86 1 2 3 dummy_cell_1rw
* cell instance $87 r0 *1 60.63,0
X$87 1 2 3 dummy_cell_1rw
* cell instance $88 r0 *1 61.335,0
X$88 1 2 3 dummy_cell_1rw
* cell instance $89 r0 *1 62.04,0
X$89 1 2 3 dummy_cell_1rw
* cell instance $90 r0 *1 62.745,0
X$90 1 2 3 dummy_cell_1rw
* cell instance $91 r0 *1 63.45,0
X$91 1 2 3 dummy_cell_1rw
* cell instance $92 r0 *1 64.155,0
X$92 1 2 3 dummy_cell_1rw
* cell instance $93 r0 *1 64.86,0
X$93 1 2 3 dummy_cell_1rw
* cell instance $94 r0 *1 65.565,0
X$94 1 2 3 dummy_cell_1rw
* cell instance $95 r0 *1 66.27,0
X$95 1 2 3 dummy_cell_1rw
* cell instance $96 r0 *1 66.975,0
X$96 1 2 3 dummy_cell_1rw
* cell instance $97 r0 *1 67.68,0
X$97 1 2 3 dummy_cell_1rw
* cell instance $98 r0 *1 68.385,0
X$98 1 2 3 dummy_cell_1rw
* cell instance $99 r0 *1 69.09,0
X$99 1 2 3 dummy_cell_1rw
* cell instance $100 r0 *1 69.795,0
X$100 1 2 3 dummy_cell_1rw
* cell instance $101 r0 *1 70.5,0
X$101 1 2 3 dummy_cell_1rw
* cell instance $102 r0 *1 71.205,0
X$102 1 2 3 dummy_cell_1rw
* cell instance $103 r0 *1 71.91,0
X$103 1 2 3 dummy_cell_1rw
* cell instance $104 r0 *1 72.615,0
X$104 1 2 3 dummy_cell_1rw
* cell instance $105 r0 *1 73.32,0
X$105 1 2 3 dummy_cell_1rw
* cell instance $106 r0 *1 74.025,0
X$106 1 2 3 dummy_cell_1rw
* cell instance $107 r0 *1 74.73,0
X$107 1 2 3 dummy_cell_1rw
* cell instance $108 r0 *1 75.435,0
X$108 1 2 3 dummy_cell_1rw
* cell instance $109 r0 *1 76.14,0
X$109 1 2 3 dummy_cell_1rw
* cell instance $110 r0 *1 76.845,0
X$110 1 2 3 dummy_cell_1rw
* cell instance $111 r0 *1 77.55,0
X$111 1 2 3 dummy_cell_1rw
* cell instance $112 r0 *1 78.255,0
X$112 1 2 3 dummy_cell_1rw
* cell instance $113 r0 *1 78.96,0
X$113 1 2 3 dummy_cell_1rw
* cell instance $114 r0 *1 79.665,0
X$114 1 2 3 dummy_cell_1rw
* cell instance $115 r0 *1 80.37,0
X$115 1 2 3 dummy_cell_1rw
* cell instance $116 r0 *1 81.075,0
X$116 1 2 3 dummy_cell_1rw
* cell instance $117 r0 *1 81.78,0
X$117 1 2 3 dummy_cell_1rw
* cell instance $118 r0 *1 82.485,0
X$118 1 2 3 dummy_cell_1rw
* cell instance $119 r0 *1 83.19,0
X$119 1 2 3 dummy_cell_1rw
* cell instance $120 r0 *1 83.895,0
X$120 1 2 3 dummy_cell_1rw
* cell instance $121 r0 *1 84.6,0
X$121 1 2 3 dummy_cell_1rw
* cell instance $122 r0 *1 85.305,0
X$122 1 2 3 dummy_cell_1rw
* cell instance $123 r0 *1 86.01,0
X$123 1 2 3 dummy_cell_1rw
* cell instance $124 r0 *1 86.715,0
X$124 1 2 3 dummy_cell_1rw
* cell instance $125 r0 *1 87.42,0
X$125 1 2 3 dummy_cell_1rw
* cell instance $126 r0 *1 88.125,0
X$126 1 2 3 dummy_cell_1rw
* cell instance $127 r0 *1 88.83,0
X$127 1 2 3 dummy_cell_1rw
* cell instance $128 r0 *1 89.535,0
X$128 1 2 3 dummy_cell_1rw
* cell instance $129 r0 *1 90.24,0
X$129 1 2 3 dummy_cell_1rw
* cell instance $130 r0 *1 90.945,0
X$130 1 2 3 dummy_cell_1rw
* cell instance $131 r0 *1 91.65,0
X$131 1 2 3 dummy_cell_1rw
* cell instance $132 r0 *1 92.355,0
X$132 1 2 3 dummy_cell_1rw
* cell instance $133 r0 *1 93.06,0
X$133 1 2 3 dummy_cell_1rw
* cell instance $134 r0 *1 93.765,0
X$134 1 2 3 dummy_cell_1rw
* cell instance $135 r0 *1 94.47,0
X$135 1 2 3 dummy_cell_1rw
* cell instance $136 r0 *1 95.175,0
X$136 1 2 3 dummy_cell_1rw
* cell instance $137 r0 *1 95.88,0
X$137 1 2 3 dummy_cell_1rw
* cell instance $138 r0 *1 96.585,0
X$138 1 2 3 dummy_cell_1rw
* cell instance $139 r0 *1 97.29,0
X$139 1 2 3 dummy_cell_1rw
* cell instance $140 r0 *1 97.995,0
X$140 1 2 3 dummy_cell_1rw
* cell instance $141 r0 *1 98.7,0
X$141 1 2 3 dummy_cell_1rw
* cell instance $142 r0 *1 99.405,0
X$142 1 2 3 dummy_cell_1rw
* cell instance $143 r0 *1 100.11,0
X$143 1 2 3 dummy_cell_1rw
* cell instance $144 r0 *1 100.815,0
X$144 1 2 3 dummy_cell_1rw
* cell instance $145 r0 *1 101.52,0
X$145 1 2 3 dummy_cell_1rw
* cell instance $146 r0 *1 102.225,0
X$146 1 2 3 dummy_cell_1rw
* cell instance $147 r0 *1 102.93,0
X$147 1 2 3 dummy_cell_1rw
* cell instance $148 r0 *1 103.635,0
X$148 1 2 3 dummy_cell_1rw
* cell instance $149 r0 *1 104.34,0
X$149 1 2 3 dummy_cell_1rw
* cell instance $150 r0 *1 105.045,0
X$150 1 2 3 dummy_cell_1rw
* cell instance $151 r0 *1 105.75,0
X$151 1 2 3 dummy_cell_1rw
* cell instance $152 r0 *1 106.455,0
X$152 1 2 3 dummy_cell_1rw
* cell instance $153 r0 *1 107.16,0
X$153 1 2 3 dummy_cell_1rw
* cell instance $154 r0 *1 107.865,0
X$154 1 2 3 dummy_cell_1rw
* cell instance $155 r0 *1 108.57,0
X$155 1 2 3 dummy_cell_1rw
* cell instance $156 r0 *1 109.275,0
X$156 1 2 3 dummy_cell_1rw
* cell instance $157 r0 *1 109.98,0
X$157 1 2 3 dummy_cell_1rw
* cell instance $158 r0 *1 110.685,0
X$158 1 2 3 dummy_cell_1rw
* cell instance $159 r0 *1 111.39,0
X$159 1 2 3 dummy_cell_1rw
* cell instance $160 r0 *1 112.095,0
X$160 1 2 3 dummy_cell_1rw
* cell instance $161 r0 *1 112.8,0
X$161 1 2 3 dummy_cell_1rw
* cell instance $162 r0 *1 113.505,0
X$162 1 2 3 dummy_cell_1rw
* cell instance $163 r0 *1 114.21,0
X$163 1 2 3 dummy_cell_1rw
* cell instance $164 r0 *1 114.915,0
X$164 1 2 3 dummy_cell_1rw
* cell instance $165 r0 *1 115.62,0
X$165 1 2 3 dummy_cell_1rw
* cell instance $166 r0 *1 116.325,0
X$166 1 2 3 dummy_cell_1rw
* cell instance $167 r0 *1 117.03,0
X$167 1 2 3 dummy_cell_1rw
* cell instance $168 r0 *1 117.735,0
X$168 1 2 3 dummy_cell_1rw
* cell instance $169 r0 *1 118.44,0
X$169 1 2 3 dummy_cell_1rw
* cell instance $170 r0 *1 119.145,0
X$170 1 2 3 dummy_cell_1rw
* cell instance $171 r0 *1 119.85,0
X$171 1 2 3 dummy_cell_1rw
* cell instance $172 r0 *1 120.555,0
X$172 1 2 3 dummy_cell_1rw
* cell instance $173 r0 *1 121.26,0
X$173 1 2 3 dummy_cell_1rw
* cell instance $174 r0 *1 121.965,0
X$174 1 2 3 dummy_cell_1rw
* cell instance $175 r0 *1 122.67,0
X$175 1 2 3 dummy_cell_1rw
* cell instance $176 r0 *1 123.375,0
X$176 1 2 3 dummy_cell_1rw
* cell instance $177 r0 *1 124.08,0
X$177 1 2 3 dummy_cell_1rw
* cell instance $178 r0 *1 124.785,0
X$178 1 2 3 dummy_cell_1rw
* cell instance $179 r0 *1 125.49,0
X$179 1 2 3 dummy_cell_1rw
* cell instance $180 r0 *1 126.195,0
X$180 1 2 3 dummy_cell_1rw
* cell instance $181 r0 *1 126.9,0
X$181 1 2 3 dummy_cell_1rw
* cell instance $182 r0 *1 127.605,0
X$182 1 2 3 dummy_cell_1rw
* cell instance $183 r0 *1 128.31,0
X$183 1 2 3 dummy_cell_1rw
* cell instance $184 r0 *1 129.015,0
X$184 1 2 3 dummy_cell_1rw
* cell instance $185 r0 *1 129.72,0
X$185 1 2 3 dummy_cell_1rw
* cell instance $186 r0 *1 130.425,0
X$186 1 2 3 dummy_cell_1rw
* cell instance $187 r0 *1 131.13,0
X$187 1 2 3 dummy_cell_1rw
* cell instance $188 r0 *1 131.835,0
X$188 1 2 3 dummy_cell_1rw
* cell instance $189 r0 *1 132.54,0
X$189 1 2 3 dummy_cell_1rw
* cell instance $190 r0 *1 133.245,0
X$190 1 2 3 dummy_cell_1rw
* cell instance $191 r0 *1 133.95,0
X$191 1 2 3 dummy_cell_1rw
* cell instance $192 r0 *1 134.655,0
X$192 1 2 3 dummy_cell_1rw
* cell instance $193 r0 *1 135.36,0
X$193 1 2 3 dummy_cell_1rw
* cell instance $194 r0 *1 136.065,0
X$194 1 2 3 dummy_cell_1rw
* cell instance $195 r0 *1 136.77,0
X$195 1 2 3 dummy_cell_1rw
* cell instance $196 r0 *1 137.475,0
X$196 1 2 3 dummy_cell_1rw
* cell instance $197 r0 *1 138.18,0
X$197 1 2 3 dummy_cell_1rw
* cell instance $198 r0 *1 138.885,0
X$198 1 2 3 dummy_cell_1rw
* cell instance $199 r0 *1 139.59,0
X$199 1 2 3 dummy_cell_1rw
* cell instance $200 r0 *1 140.295,0
X$200 1 2 3 dummy_cell_1rw
* cell instance $201 r0 *1 141,0
X$201 1 2 3 dummy_cell_1rw
* cell instance $202 r0 *1 141.705,0
X$202 1 2 3 dummy_cell_1rw
* cell instance $203 r0 *1 142.41,0
X$203 1 2 3 dummy_cell_1rw
* cell instance $204 r0 *1 143.115,0
X$204 1 2 3 dummy_cell_1rw
* cell instance $205 r0 *1 143.82,0
X$205 1 2 3 dummy_cell_1rw
* cell instance $206 r0 *1 144.525,0
X$206 1 2 3 dummy_cell_1rw
* cell instance $207 r0 *1 145.23,0
X$207 1 2 3 dummy_cell_1rw
* cell instance $208 r0 *1 145.935,0
X$208 1 2 3 dummy_cell_1rw
* cell instance $209 r0 *1 146.64,0
X$209 1 2 3 dummy_cell_1rw
* cell instance $210 r0 *1 147.345,0
X$210 1 2 3 dummy_cell_1rw
* cell instance $211 r0 *1 148.05,0
X$211 1 2 3 dummy_cell_1rw
* cell instance $212 r0 *1 148.755,0
X$212 1 2 3 dummy_cell_1rw
* cell instance $213 r0 *1 149.46,0
X$213 1 2 3 dummy_cell_1rw
* cell instance $214 r0 *1 150.165,0
X$214 1 2 3 dummy_cell_1rw
* cell instance $215 r0 *1 150.87,0
X$215 1 2 3 dummy_cell_1rw
* cell instance $216 r0 *1 151.575,0
X$216 1 2 3 dummy_cell_1rw
* cell instance $217 r0 *1 152.28,0
X$217 1 2 3 dummy_cell_1rw
* cell instance $218 r0 *1 152.985,0
X$218 1 2 3 dummy_cell_1rw
* cell instance $219 r0 *1 153.69,0
X$219 1 2 3 dummy_cell_1rw
* cell instance $220 r0 *1 154.395,0
X$220 1 2 3 dummy_cell_1rw
* cell instance $221 r0 *1 155.1,0
X$221 1 2 3 dummy_cell_1rw
* cell instance $222 r0 *1 155.805,0
X$222 1 2 3 dummy_cell_1rw
* cell instance $223 r0 *1 156.51,0
X$223 1 2 3 dummy_cell_1rw
* cell instance $224 r0 *1 157.215,0
X$224 1 2 3 dummy_cell_1rw
* cell instance $225 r0 *1 157.92,0
X$225 1 2 3 dummy_cell_1rw
* cell instance $226 r0 *1 158.625,0
X$226 1 2 3 dummy_cell_1rw
* cell instance $227 r0 *1 159.33,0
X$227 1 2 3 dummy_cell_1rw
* cell instance $228 r0 *1 160.035,0
X$228 1 2 3 dummy_cell_1rw
* cell instance $229 r0 *1 160.74,0
X$229 1 2 3 dummy_cell_1rw
* cell instance $230 r0 *1 161.445,0
X$230 1 2 3 dummy_cell_1rw
* cell instance $231 r0 *1 162.15,0
X$231 1 2 3 dummy_cell_1rw
* cell instance $232 r0 *1 162.855,0
X$232 1 2 3 dummy_cell_1rw
* cell instance $233 r0 *1 163.56,0
X$233 1 2 3 dummy_cell_1rw
* cell instance $234 r0 *1 164.265,0
X$234 1 2 3 dummy_cell_1rw
* cell instance $235 r0 *1 164.97,0
X$235 1 2 3 dummy_cell_1rw
* cell instance $236 r0 *1 165.675,0
X$236 1 2 3 dummy_cell_1rw
* cell instance $237 r0 *1 166.38,0
X$237 1 2 3 dummy_cell_1rw
* cell instance $238 r0 *1 167.085,0
X$238 1 2 3 dummy_cell_1rw
* cell instance $239 r0 *1 167.79,0
X$239 1 2 3 dummy_cell_1rw
* cell instance $240 r0 *1 168.495,0
X$240 1 2 3 dummy_cell_1rw
* cell instance $241 r0 *1 169.2,0
X$241 1 2 3 dummy_cell_1rw
* cell instance $242 r0 *1 169.905,0
X$242 1 2 3 dummy_cell_1rw
* cell instance $243 r0 *1 170.61,0
X$243 1 2 3 dummy_cell_1rw
* cell instance $244 r0 *1 171.315,0
X$244 1 2 3 dummy_cell_1rw
* cell instance $245 r0 *1 172.02,0
X$245 1 2 3 dummy_cell_1rw
* cell instance $246 r0 *1 172.725,0
X$246 1 2 3 dummy_cell_1rw
* cell instance $247 r0 *1 173.43,0
X$247 1 2 3 dummy_cell_1rw
* cell instance $248 r0 *1 174.135,0
X$248 1 2 3 dummy_cell_1rw
* cell instance $249 r0 *1 174.84,0
X$249 1 2 3 dummy_cell_1rw
* cell instance $250 r0 *1 175.545,0
X$250 1 2 3 dummy_cell_1rw
* cell instance $251 r0 *1 176.25,0
X$251 1 2 3 dummy_cell_1rw
* cell instance $252 r0 *1 176.955,0
X$252 1 2 3 dummy_cell_1rw
* cell instance $253 r0 *1 177.66,0
X$253 1 2 3 dummy_cell_1rw
* cell instance $254 r0 *1 178.365,0
X$254 1 2 3 dummy_cell_1rw
* cell instance $255 r0 *1 179.07,0
X$255 1 2 3 dummy_cell_1rw
* cell instance $256 r0 *1 179.775,0
X$256 1 2 3 dummy_cell_1rw
* cell instance $257 r0 *1 180.48,0
X$257 1 2 3 dummy_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_dummy_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_replica_column
* pin wl_0_0
* pin wl_0_1
* pin wl_0_2
* pin wl_0_3
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_8
* pin wl_0_9
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_24
* pin wl_0_25
* pin wl_0_26
* pin wl_0_27
* pin wl_0_28
* pin wl_0_29
* pin wl_0_30
* pin wl_0_31
* pin wl_0_32
* pin wl_0_33
* pin wl_0_34
* pin wl_0_35
* pin wl_0_36
* pin wl_0_37
* pin wl_0_38
* pin wl_0_39
* pin wl_0_40
* pin wl_0_41
* pin wl_0_42
* pin wl_0_43
* pin wl_0_44
* pin wl_0_45
* pin wl_0_46
* pin wl_0_47
* pin wl_0_48
* pin wl_0_49
* pin wl_0_50
* pin wl_0_51
* pin wl_0_52
* pin wl_0_53
* pin wl_0_54
* pin wl_0_55
* pin wl_0_56
* pin wl_0_57
* pin wl_0_58
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_62
* pin wl_0_63
* pin bl_0_0
* pin wl_0_64
* pin br_0_0
* pin wl_0_65
* pin wl_0_66
* pin wl_0_67
* pin wl_0_68
* pin wl_0_69
* pin wl_0_70
* pin wl_0_71
* pin wl_0_72
* pin wl_0_73
* pin wl_0_74
* pin wl_0_75
* pin wl_0_76
* pin wl_0_77
* pin wl_0_78
* pin wl_0_79
* pin wl_0_80
* pin wl_0_81
* pin wl_0_82
* pin wl_0_83
* pin wl_0_84
* pin wl_0_85
* pin wl_0_86
* pin wl_0_87
* pin wl_0_88
* pin wl_0_89
* pin wl_0_90
* pin wl_0_91
* pin wl_0_92
* pin wl_0_93
* pin wl_0_94
* pin wl_0_95
* pin wl_0_96
* pin wl_0_97
* pin wl_0_98
* pin wl_0_99
* pin wl_0_100
* pin wl_0_101
* pin wl_0_102
* pin wl_0_103
* pin wl_0_104
* pin wl_0_105
* pin wl_0_106
* pin wl_0_107
* pin wl_0_108
* pin wl_0_109
* pin wl_0_110
* pin wl_0_111
* pin wl_0_112
* pin wl_0_113
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_117
* pin wl_0_118
* pin wl_0_119
* pin wl_0_120
* pin wl_0_121
* pin wl_0_122
* pin wl_0_123
* pin wl_0_124
* pin wl_0_125
* pin wl_0_126
* pin wl_0_127
* pin wl_0_128
* pin wl_0_129
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_replica_column 1 2 3 4 5 6 7 8 9
+ 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35
+ 36 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87
+ 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109
+ 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128
+ 129 130 131 132 133 134
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_2
* net 4 wl_0_3
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_8
* net 10 wl_0_9
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 wl_0_19
* net 21 wl_0_20
* net 22 wl_0_21
* net 23 wl_0_22
* net 24 wl_0_23
* net 25 wl_0_24
* net 26 wl_0_25
* net 27 wl_0_26
* net 28 wl_0_27
* net 29 wl_0_28
* net 30 wl_0_29
* net 31 wl_0_30
* net 32 wl_0_31
* net 33 wl_0_32
* net 34 wl_0_33
* net 35 wl_0_34
* net 36 wl_0_35
* net 37 wl_0_36
* net 38 wl_0_37
* net 39 wl_0_38
* net 40 wl_0_39
* net 41 wl_0_40
* net 42 wl_0_41
* net 43 wl_0_42
* net 44 wl_0_43
* net 45 wl_0_44
* net 46 wl_0_45
* net 47 wl_0_46
* net 48 wl_0_47
* net 49 wl_0_48
* net 50 wl_0_49
* net 51 wl_0_50
* net 52 wl_0_51
* net 53 wl_0_52
* net 54 wl_0_53
* net 55 wl_0_54
* net 56 wl_0_55
* net 57 wl_0_56
* net 58 wl_0_57
* net 59 wl_0_58
* net 60 wl_0_59
* net 61 wl_0_60
* net 62 wl_0_61
* net 63 wl_0_62
* net 64 wl_0_63
* net 65 bl_0_0
* net 66 wl_0_64
* net 67 br_0_0
* net 68 wl_0_65
* net 69 wl_0_66
* net 70 wl_0_67
* net 71 wl_0_68
* net 72 wl_0_69
* net 73 wl_0_70
* net 74 wl_0_71
* net 75 wl_0_72
* net 76 wl_0_73
* net 77 wl_0_74
* net 78 wl_0_75
* net 79 wl_0_76
* net 80 wl_0_77
* net 81 wl_0_78
* net 82 wl_0_79
* net 83 wl_0_80
* net 84 wl_0_81
* net 85 wl_0_82
* net 86 wl_0_83
* net 87 wl_0_84
* net 88 wl_0_85
* net 89 wl_0_86
* net 90 wl_0_87
* net 91 wl_0_88
* net 92 wl_0_89
* net 93 wl_0_90
* net 94 wl_0_91
* net 95 wl_0_92
* net 96 wl_0_93
* net 97 wl_0_94
* net 98 wl_0_95
* net 99 wl_0_96
* net 100 wl_0_97
* net 101 wl_0_98
* net 102 wl_0_99
* net 103 wl_0_100
* net 104 wl_0_101
* net 105 wl_0_102
* net 106 wl_0_103
* net 107 wl_0_104
* net 108 wl_0_105
* net 109 wl_0_106
* net 110 wl_0_107
* net 111 wl_0_108
* net 112 wl_0_109
* net 113 wl_0_110
* net 114 wl_0_111
* net 115 wl_0_112
* net 116 wl_0_113
* net 117 wl_0_114
* net 118 wl_0_115
* net 119 wl_0_116
* net 120 wl_0_117
* net 121 wl_0_118
* net 122 wl_0_119
* net 123 wl_0_120
* net 124 wl_0_121
* net 125 wl_0_122
* net 126 wl_0_123
* net 127 wl_0_124
* net 128 wl_0_125
* net 129 wl_0_126
* net 130 wl_0_127
* net 131 wl_0_128
* net 132 wl_0_129
* net 133 vdd
* net 134 gnd
* cell instance $1 m0 *1 0,1.365
X$1 65 1 67 133 134 replica_cell_1rw
* cell instance $2 r0 *1 0,1.365
X$2 65 2 67 133 134 replica_cell_1rw
* cell instance $3 m0 *1 0,4.095
X$3 65 3 67 133 134 replica_cell_1rw
* cell instance $4 r0 *1 0,4.095
X$4 65 4 67 133 134 replica_cell_1rw
* cell instance $5 m0 *1 0,6.825
X$5 65 5 67 133 134 replica_cell_1rw
* cell instance $6 r0 *1 0,6.825
X$6 65 6 67 133 134 replica_cell_1rw
* cell instance $7 m0 *1 0,9.555
X$7 65 7 67 133 134 replica_cell_1rw
* cell instance $8 r0 *1 0,9.555
X$8 65 8 67 133 134 replica_cell_1rw
* cell instance $9 m0 *1 0,12.285
X$9 65 9 67 133 134 replica_cell_1rw
* cell instance $10 r0 *1 0,12.285
X$10 65 10 67 133 134 replica_cell_1rw
* cell instance $11 m0 *1 0,15.015
X$11 65 11 67 133 134 replica_cell_1rw
* cell instance $12 r0 *1 0,15.015
X$12 65 12 67 133 134 replica_cell_1rw
* cell instance $13 m0 *1 0,17.745
X$13 65 13 67 133 134 replica_cell_1rw
* cell instance $14 r0 *1 0,17.745
X$14 65 14 67 133 134 replica_cell_1rw
* cell instance $15 m0 *1 0,20.475
X$15 65 15 67 133 134 replica_cell_1rw
* cell instance $16 r0 *1 0,20.475
X$16 65 16 67 133 134 replica_cell_1rw
* cell instance $17 m0 *1 0,23.205
X$17 65 17 67 133 134 replica_cell_1rw
* cell instance $18 r0 *1 0,23.205
X$18 65 18 67 133 134 replica_cell_1rw
* cell instance $19 m0 *1 0,25.935
X$19 65 19 67 133 134 replica_cell_1rw
* cell instance $20 r0 *1 0,25.935
X$20 65 20 67 133 134 replica_cell_1rw
* cell instance $21 m0 *1 0,28.665
X$21 65 21 67 133 134 replica_cell_1rw
* cell instance $22 r0 *1 0,28.665
X$22 65 22 67 133 134 replica_cell_1rw
* cell instance $23 m0 *1 0,31.395
X$23 65 23 67 133 134 replica_cell_1rw
* cell instance $24 r0 *1 0,31.395
X$24 65 24 67 133 134 replica_cell_1rw
* cell instance $25 m0 *1 0,34.125
X$25 65 25 67 133 134 replica_cell_1rw
* cell instance $26 r0 *1 0,34.125
X$26 65 26 67 133 134 replica_cell_1rw
* cell instance $27 m0 *1 0,36.855
X$27 65 27 67 133 134 replica_cell_1rw
* cell instance $28 r0 *1 0,36.855
X$28 65 28 67 133 134 replica_cell_1rw
* cell instance $29 m0 *1 0,39.585
X$29 65 29 67 133 134 replica_cell_1rw
* cell instance $30 r0 *1 0,39.585
X$30 65 30 67 133 134 replica_cell_1rw
* cell instance $31 m0 *1 0,42.315
X$31 65 31 67 133 134 replica_cell_1rw
* cell instance $32 r0 *1 0,42.315
X$32 65 32 67 133 134 replica_cell_1rw
* cell instance $33 m0 *1 0,45.045
X$33 65 33 67 133 134 replica_cell_1rw
* cell instance $34 r0 *1 0,45.045
X$34 65 34 67 133 134 replica_cell_1rw
* cell instance $35 m0 *1 0,47.775
X$35 65 35 67 133 134 replica_cell_1rw
* cell instance $36 r0 *1 0,47.775
X$36 65 36 67 133 134 replica_cell_1rw
* cell instance $37 m0 *1 0,50.505
X$37 65 37 67 133 134 replica_cell_1rw
* cell instance $38 r0 *1 0,50.505
X$38 65 38 67 133 134 replica_cell_1rw
* cell instance $39 m0 *1 0,53.235
X$39 65 39 67 133 134 replica_cell_1rw
* cell instance $40 r0 *1 0,53.235
X$40 65 40 67 133 134 replica_cell_1rw
* cell instance $41 m0 *1 0,55.965
X$41 65 41 67 133 134 replica_cell_1rw
* cell instance $42 r0 *1 0,55.965
X$42 65 42 67 133 134 replica_cell_1rw
* cell instance $43 m0 *1 0,58.695
X$43 65 43 67 133 134 replica_cell_1rw
* cell instance $44 r0 *1 0,58.695
X$44 65 44 67 133 134 replica_cell_1rw
* cell instance $45 m0 *1 0,61.425
X$45 65 45 67 133 134 replica_cell_1rw
* cell instance $46 r0 *1 0,61.425
X$46 65 46 67 133 134 replica_cell_1rw
* cell instance $47 m0 *1 0,64.155
X$47 65 47 67 133 134 replica_cell_1rw
* cell instance $48 r0 *1 0,64.155
X$48 65 48 67 133 134 replica_cell_1rw
* cell instance $49 m0 *1 0,66.885
X$49 65 49 67 133 134 replica_cell_1rw
* cell instance $50 r0 *1 0,66.885
X$50 65 50 67 133 134 replica_cell_1rw
* cell instance $51 m0 *1 0,69.615
X$51 65 51 67 133 134 replica_cell_1rw
* cell instance $52 r0 *1 0,69.615
X$52 65 52 67 133 134 replica_cell_1rw
* cell instance $53 m0 *1 0,72.345
X$53 65 53 67 133 134 replica_cell_1rw
* cell instance $54 r0 *1 0,72.345
X$54 65 54 67 133 134 replica_cell_1rw
* cell instance $55 m0 *1 0,75.075
X$55 65 55 67 133 134 replica_cell_1rw
* cell instance $56 r0 *1 0,75.075
X$56 65 56 67 133 134 replica_cell_1rw
* cell instance $57 m0 *1 0,77.805
X$57 65 57 67 133 134 replica_cell_1rw
* cell instance $58 r0 *1 0,77.805
X$58 65 58 67 133 134 replica_cell_1rw
* cell instance $59 m0 *1 0,80.535
X$59 65 59 67 133 134 replica_cell_1rw
* cell instance $60 r0 *1 0,80.535
X$60 65 60 67 133 134 replica_cell_1rw
* cell instance $61 m0 *1 0,83.265
X$61 65 61 67 133 134 replica_cell_1rw
* cell instance $62 r0 *1 0,83.265
X$62 65 62 67 133 134 replica_cell_1rw
* cell instance $63 m0 *1 0,85.995
X$63 65 63 67 133 134 replica_cell_1rw
* cell instance $64 r0 *1 0,85.995
X$64 65 64 67 133 134 replica_cell_1rw
* cell instance $65 m0 *1 0,88.725
X$65 65 66 67 133 134 replica_cell_1rw
* cell instance $66 r0 *1 0,88.725
X$66 65 68 67 133 134 replica_cell_1rw
* cell instance $67 m0 *1 0,91.455
X$67 65 69 67 133 134 replica_cell_1rw
* cell instance $68 r0 *1 0,91.455
X$68 65 70 67 133 134 replica_cell_1rw
* cell instance $69 m0 *1 0,94.185
X$69 65 71 67 133 134 replica_cell_1rw
* cell instance $70 r0 *1 0,94.185
X$70 65 72 67 133 134 replica_cell_1rw
* cell instance $71 m0 *1 0,96.915
X$71 65 73 67 133 134 replica_cell_1rw
* cell instance $72 r0 *1 0,96.915
X$72 65 74 67 133 134 replica_cell_1rw
* cell instance $73 m0 *1 0,99.645
X$73 65 75 67 133 134 replica_cell_1rw
* cell instance $74 r0 *1 0,99.645
X$74 65 76 67 133 134 replica_cell_1rw
* cell instance $75 m0 *1 0,102.375
X$75 65 77 67 133 134 replica_cell_1rw
* cell instance $76 r0 *1 0,102.375
X$76 65 78 67 133 134 replica_cell_1rw
* cell instance $77 m0 *1 0,105.105
X$77 65 79 67 133 134 replica_cell_1rw
* cell instance $78 r0 *1 0,105.105
X$78 65 80 67 133 134 replica_cell_1rw
* cell instance $79 m0 *1 0,107.835
X$79 65 81 67 133 134 replica_cell_1rw
* cell instance $80 r0 *1 0,107.835
X$80 65 82 67 133 134 replica_cell_1rw
* cell instance $81 m0 *1 0,110.565
X$81 65 83 67 133 134 replica_cell_1rw
* cell instance $82 r0 *1 0,110.565
X$82 65 84 67 133 134 replica_cell_1rw
* cell instance $83 m0 *1 0,113.295
X$83 65 85 67 133 134 replica_cell_1rw
* cell instance $84 r0 *1 0,113.295
X$84 65 86 67 133 134 replica_cell_1rw
* cell instance $85 m0 *1 0,116.025
X$85 65 87 67 133 134 replica_cell_1rw
* cell instance $86 r0 *1 0,116.025
X$86 65 88 67 133 134 replica_cell_1rw
* cell instance $87 m0 *1 0,118.755
X$87 65 89 67 133 134 replica_cell_1rw
* cell instance $88 r0 *1 0,118.755
X$88 65 90 67 133 134 replica_cell_1rw
* cell instance $89 m0 *1 0,121.485
X$89 65 91 67 133 134 replica_cell_1rw
* cell instance $90 r0 *1 0,121.485
X$90 65 92 67 133 134 replica_cell_1rw
* cell instance $91 m0 *1 0,124.215
X$91 65 93 67 133 134 replica_cell_1rw
* cell instance $92 r0 *1 0,124.215
X$92 65 94 67 133 134 replica_cell_1rw
* cell instance $93 m0 *1 0,126.945
X$93 65 95 67 133 134 replica_cell_1rw
* cell instance $94 r0 *1 0,126.945
X$94 65 96 67 133 134 replica_cell_1rw
* cell instance $95 m0 *1 0,129.675
X$95 65 97 67 133 134 replica_cell_1rw
* cell instance $96 r0 *1 0,129.675
X$96 65 98 67 133 134 replica_cell_1rw
* cell instance $97 m0 *1 0,132.405
X$97 65 99 67 133 134 replica_cell_1rw
* cell instance $98 r0 *1 0,132.405
X$98 65 100 67 133 134 replica_cell_1rw
* cell instance $99 m0 *1 0,135.135
X$99 65 101 67 133 134 replica_cell_1rw
* cell instance $100 r0 *1 0,135.135
X$100 65 102 67 133 134 replica_cell_1rw
* cell instance $101 m0 *1 0,137.865
X$101 65 103 67 133 134 replica_cell_1rw
* cell instance $102 r0 *1 0,137.865
X$102 65 104 67 133 134 replica_cell_1rw
* cell instance $103 m0 *1 0,140.595
X$103 65 105 67 133 134 replica_cell_1rw
* cell instance $104 r0 *1 0,140.595
X$104 65 106 67 133 134 replica_cell_1rw
* cell instance $105 m0 *1 0,143.325
X$105 65 107 67 133 134 replica_cell_1rw
* cell instance $106 r0 *1 0,143.325
X$106 65 108 67 133 134 replica_cell_1rw
* cell instance $107 m0 *1 0,146.055
X$107 65 109 67 133 134 replica_cell_1rw
* cell instance $108 r0 *1 0,146.055
X$108 65 110 67 133 134 replica_cell_1rw
* cell instance $109 m0 *1 0,148.785
X$109 65 111 67 133 134 replica_cell_1rw
* cell instance $110 r0 *1 0,148.785
X$110 65 112 67 133 134 replica_cell_1rw
* cell instance $111 m0 *1 0,151.515
X$111 65 113 67 133 134 replica_cell_1rw
* cell instance $112 r0 *1 0,151.515
X$112 65 114 67 133 134 replica_cell_1rw
* cell instance $113 m0 *1 0,154.245
X$113 65 115 67 133 134 replica_cell_1rw
* cell instance $114 r0 *1 0,154.245
X$114 65 116 67 133 134 replica_cell_1rw
* cell instance $115 m0 *1 0,156.975
X$115 65 117 67 133 134 replica_cell_1rw
* cell instance $116 r0 *1 0,156.975
X$116 65 118 67 133 134 replica_cell_1rw
* cell instance $117 m0 *1 0,159.705
X$117 65 119 67 133 134 replica_cell_1rw
* cell instance $118 r0 *1 0,159.705
X$118 65 120 67 133 134 replica_cell_1rw
* cell instance $119 m0 *1 0,162.435
X$119 65 121 67 133 134 replica_cell_1rw
* cell instance $120 r0 *1 0,162.435
X$120 65 122 67 133 134 replica_cell_1rw
* cell instance $121 m0 *1 0,165.165
X$121 65 123 67 133 134 replica_cell_1rw
* cell instance $122 r0 *1 0,165.165
X$122 65 124 67 133 134 replica_cell_1rw
* cell instance $123 m0 *1 0,167.895
X$123 65 125 67 133 134 replica_cell_1rw
* cell instance $124 r0 *1 0,167.895
X$124 65 126 67 133 134 replica_cell_1rw
* cell instance $125 m0 *1 0,170.625
X$125 65 127 67 133 134 replica_cell_1rw
* cell instance $126 r0 *1 0,170.625
X$126 65 128 67 133 134 replica_cell_1rw
* cell instance $127 m0 *1 0,173.355
X$127 65 129 67 133 134 replica_cell_1rw
* cell instance $128 r0 *1 0,173.355
X$128 65 130 67 133 134 replica_cell_1rw
* cell instance $129 m0 *1 0,176.085
X$129 65 131 67 133 134 replica_cell_1rw
* cell instance $130 r0 *1 0,176.085
X$130 65 132 67 133 134 replica_cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_replica_column

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_bitcell_array
* pin wl_0_0
* pin wl_0_1
* pin wl_0_3
* pin wl_0_2
* pin wl_0_4
* pin wl_0_5
* pin wl_0_6
* pin wl_0_7
* pin wl_0_9
* pin wl_0_8
* pin wl_0_10
* pin wl_0_11
* pin wl_0_12
* pin wl_0_13
* pin wl_0_14
* pin wl_0_15
* pin wl_0_16
* pin wl_0_17
* pin wl_0_18
* pin wl_0_19
* pin wl_0_20
* pin wl_0_21
* pin wl_0_22
* pin wl_0_23
* pin wl_0_25
* pin wl_0_24
* pin wl_0_26
* pin wl_0_27
* pin wl_0_28
* pin wl_0_29
* pin wl_0_30
* pin wl_0_31
* pin wl_0_32
* pin wl_0_33
* pin wl_0_34
* pin wl_0_35
* pin wl_0_36
* pin wl_0_37
* pin wl_0_39
* pin wl_0_38
* pin wl_0_41
* pin wl_0_40
* pin wl_0_43
* pin wl_0_42
* pin wl_0_44
* pin wl_0_45
* pin wl_0_46
* pin wl_0_47
* pin wl_0_48
* pin wl_0_49
* pin wl_0_50
* pin wl_0_51
* pin wl_0_52
* pin wl_0_53
* pin wl_0_54
* pin wl_0_55
* pin wl_0_56
* pin wl_0_57
* pin wl_0_58
* pin wl_0_59
* pin wl_0_60
* pin wl_0_61
* pin wl_0_62
* pin wl_0_63
* pin bl_0_0
* pin br_0_0
* pin bl_0_1
* pin br_0_1
* pin bl_0_2
* pin br_0_2
* pin bl_0_3
* pin br_0_3
* pin bl_0_4
* pin br_0_4
* pin bl_0_5
* pin br_0_5
* pin bl_0_6
* pin br_0_6
* pin bl_0_7
* pin br_0_7
* pin bl_0_8
* pin br_0_8
* pin bl_0_9
* pin br_0_9
* pin bl_0_10
* pin br_0_10
* pin bl_0_11
* pin br_0_11
* pin bl_0_12
* pin br_0_12
* pin bl_0_13
* pin br_0_13
* pin bl_0_14
* pin br_0_14
* pin bl_0_15
* pin br_0_15
* pin bl_0_16
* pin br_0_16
* pin bl_0_17
* pin br_0_17
* pin bl_0_18
* pin br_0_18
* pin bl_0_19
* pin br_0_19
* pin bl_0_20
* pin br_0_20
* pin bl_0_21
* pin br_0_21
* pin bl_0_22
* pin br_0_22
* pin bl_0_23
* pin br_0_23
* pin bl_0_24
* pin br_0_24
* pin bl_0_25
* pin br_0_25
* pin bl_0_26
* pin br_0_26
* pin bl_0_27
* pin br_0_27
* pin bl_0_28
* pin br_0_28
* pin bl_0_29
* pin br_0_29
* pin bl_0_30
* pin br_0_30
* pin bl_0_31
* pin br_0_31
* pin bl_0_32
* pin br_0_32
* pin bl_0_33
* pin br_0_33
* pin bl_0_34
* pin br_0_34
* pin bl_0_35
* pin br_0_35
* pin bl_0_36
* pin br_0_36
* pin bl_0_37
* pin br_0_37
* pin bl_0_38
* pin br_0_38
* pin bl_0_39
* pin br_0_39
* pin bl_0_40
* pin br_0_40
* pin bl_0_41
* pin br_0_41
* pin bl_0_42
* pin br_0_42
* pin bl_0_43
* pin br_0_43
* pin bl_0_44
* pin br_0_44
* pin bl_0_45
* pin br_0_45
* pin bl_0_46
* pin br_0_46
* pin bl_0_47
* pin br_0_47
* pin bl_0_48
* pin br_0_48
* pin bl_0_49
* pin br_0_49
* pin bl_0_50
* pin br_0_50
* pin bl_0_51
* pin br_0_51
* pin bl_0_52
* pin br_0_52
* pin bl_0_53
* pin br_0_53
* pin bl_0_54
* pin br_0_54
* pin bl_0_55
* pin br_0_55
* pin bl_0_56
* pin br_0_56
* pin bl_0_57
* pin br_0_57
* pin bl_0_58
* pin br_0_58
* pin bl_0_59
* pin br_0_59
* pin bl_0_60
* pin br_0_60
* pin bl_0_61
* pin br_0_61
* pin bl_0_62
* pin br_0_62
* pin bl_0_63
* pin br_0_63
* pin bl_0_64
* pin br_0_64
* pin bl_0_65
* pin br_0_65
* pin bl_0_66
* pin br_0_66
* pin bl_0_67
* pin br_0_67
* pin bl_0_68
* pin br_0_68
* pin bl_0_69
* pin br_0_69
* pin bl_0_70
* pin br_0_70
* pin bl_0_71
* pin br_0_71
* pin bl_0_72
* pin br_0_72
* pin bl_0_73
* pin br_0_73
* pin bl_0_74
* pin br_0_74
* pin bl_0_75
* pin br_0_75
* pin bl_0_76
* pin br_0_76
* pin bl_0_77
* pin br_0_77
* pin bl_0_78
* pin br_0_78
* pin bl_0_79
* pin br_0_79
* pin bl_0_80
* pin br_0_80
* pin bl_0_81
* pin br_0_81
* pin bl_0_82
* pin br_0_82
* pin bl_0_83
* pin br_0_83
* pin bl_0_84
* pin br_0_84
* pin bl_0_85
* pin br_0_85
* pin bl_0_86
* pin br_0_86
* pin bl_0_87
* pin br_0_87
* pin bl_0_88
* pin br_0_88
* pin bl_0_89
* pin br_0_89
* pin bl_0_90
* pin br_0_90
* pin bl_0_91
* pin br_0_91
* pin bl_0_92
* pin br_0_92
* pin bl_0_93
* pin br_0_93
* pin bl_0_94
* pin br_0_94
* pin bl_0_95
* pin br_0_95
* pin bl_0_96
* pin br_0_96
* pin bl_0_97
* pin br_0_97
* pin bl_0_98
* pin br_0_98
* pin bl_0_99
* pin br_0_99
* pin bl_0_100
* pin br_0_100
* pin bl_0_101
* pin br_0_101
* pin bl_0_102
* pin br_0_102
* pin bl_0_103
* pin br_0_103
* pin bl_0_104
* pin br_0_104
* pin bl_0_105
* pin br_0_105
* pin bl_0_106
* pin br_0_106
* pin bl_0_107
* pin br_0_107
* pin bl_0_108
* pin br_0_108
* pin bl_0_109
* pin br_0_109
* pin bl_0_110
* pin br_0_110
* pin bl_0_111
* pin br_0_111
* pin bl_0_112
* pin br_0_112
* pin bl_0_113
* pin br_0_113
* pin bl_0_114
* pin br_0_114
* pin bl_0_115
* pin br_0_115
* pin bl_0_116
* pin br_0_116
* pin bl_0_117
* pin br_0_117
* pin bl_0_118
* pin br_0_118
* pin bl_0_119
* pin br_0_119
* pin bl_0_120
* pin br_0_120
* pin bl_0_121
* pin br_0_121
* pin bl_0_122
* pin br_0_122
* pin bl_0_123
* pin br_0_123
* pin bl_0_124
* pin br_0_124
* pin bl_0_125
* pin br_0_125
* pin bl_0_126
* pin br_0_126
* pin bl_0_127
* pin br_0_127
* pin bl_0_128
* pin wl_0_64
* pin br_0_128
* pin bl_0_129
* pin br_0_129
* pin bl_0_130
* pin br_0_130
* pin bl_0_131
* pin br_0_131
* pin bl_0_132
* pin br_0_132
* pin bl_0_133
* pin br_0_133
* pin bl_0_134
* pin br_0_134
* pin bl_0_135
* pin br_0_135
* pin bl_0_136
* pin br_0_136
* pin bl_0_137
* pin br_0_137
* pin bl_0_138
* pin br_0_138
* pin bl_0_139
* pin br_0_139
* pin bl_0_140
* pin br_0_140
* pin bl_0_141
* pin br_0_141
* pin bl_0_142
* pin br_0_142
* pin bl_0_143
* pin br_0_143
* pin bl_0_144
* pin br_0_144
* pin bl_0_145
* pin br_0_145
* pin bl_0_146
* pin br_0_146
* pin bl_0_147
* pin br_0_147
* pin bl_0_148
* pin br_0_148
* pin bl_0_149
* pin br_0_149
* pin bl_0_150
* pin br_0_150
* pin bl_0_151
* pin br_0_151
* pin bl_0_152
* pin br_0_152
* pin bl_0_153
* pin br_0_153
* pin bl_0_154
* pin br_0_154
* pin bl_0_155
* pin br_0_155
* pin bl_0_156
* pin br_0_156
* pin bl_0_157
* pin br_0_157
* pin bl_0_158
* pin br_0_158
* pin bl_0_159
* pin br_0_159
* pin bl_0_160
* pin br_0_160
* pin bl_0_161
* pin br_0_161
* pin bl_0_162
* pin br_0_162
* pin bl_0_163
* pin br_0_163
* pin bl_0_164
* pin br_0_164
* pin bl_0_165
* pin br_0_165
* pin bl_0_166
* pin br_0_166
* pin bl_0_167
* pin br_0_167
* pin bl_0_168
* pin br_0_168
* pin bl_0_169
* pin br_0_169
* pin bl_0_170
* pin br_0_170
* pin bl_0_171
* pin br_0_171
* pin bl_0_172
* pin br_0_172
* pin bl_0_173
* pin br_0_173
* pin bl_0_174
* pin br_0_174
* pin bl_0_175
* pin br_0_175
* pin bl_0_176
* pin br_0_176
* pin bl_0_177
* pin br_0_177
* pin bl_0_178
* pin br_0_178
* pin bl_0_179
* pin br_0_179
* pin bl_0_180
* pin br_0_180
* pin bl_0_181
* pin br_0_181
* pin bl_0_182
* pin br_0_182
* pin bl_0_183
* pin br_0_183
* pin bl_0_184
* pin br_0_184
* pin bl_0_185
* pin br_0_185
* pin bl_0_186
* pin br_0_186
* pin bl_0_187
* pin br_0_187
* pin bl_0_188
* pin br_0_188
* pin bl_0_189
* pin br_0_189
* pin bl_0_190
* pin br_0_190
* pin bl_0_191
* pin br_0_191
* pin bl_0_192
* pin br_0_192
* pin bl_0_193
* pin br_0_193
* pin bl_0_194
* pin br_0_194
* pin bl_0_195
* pin br_0_195
* pin bl_0_196
* pin br_0_196
* pin bl_0_197
* pin br_0_197
* pin bl_0_198
* pin br_0_198
* pin bl_0_199
* pin br_0_199
* pin bl_0_200
* pin br_0_200
* pin bl_0_201
* pin br_0_201
* pin bl_0_202
* pin br_0_202
* pin bl_0_203
* pin br_0_203
* pin bl_0_204
* pin br_0_204
* pin bl_0_205
* pin br_0_205
* pin bl_0_206
* pin br_0_206
* pin bl_0_207
* pin br_0_207
* pin bl_0_208
* pin br_0_208
* pin bl_0_209
* pin br_0_209
* pin bl_0_210
* pin br_0_210
* pin bl_0_211
* pin br_0_211
* pin bl_0_212
* pin br_0_212
* pin bl_0_213
* pin br_0_213
* pin bl_0_214
* pin br_0_214
* pin bl_0_215
* pin br_0_215
* pin bl_0_216
* pin br_0_216
* pin bl_0_217
* pin br_0_217
* pin bl_0_218
* pin br_0_218
* pin bl_0_219
* pin br_0_219
* pin bl_0_220
* pin br_0_220
* pin bl_0_221
* pin br_0_221
* pin bl_0_222
* pin br_0_222
* pin bl_0_223
* pin br_0_223
* pin bl_0_224
* pin br_0_224
* pin bl_0_225
* pin br_0_225
* pin bl_0_226
* pin br_0_226
* pin bl_0_227
* pin br_0_227
* pin bl_0_228
* pin br_0_228
* pin bl_0_229
* pin br_0_229
* pin bl_0_230
* pin br_0_230
* pin bl_0_231
* pin br_0_231
* pin bl_0_232
* pin br_0_232
* pin bl_0_233
* pin br_0_233
* pin bl_0_234
* pin br_0_234
* pin bl_0_235
* pin br_0_235
* pin bl_0_236
* pin br_0_236
* pin bl_0_237
* pin br_0_237
* pin bl_0_238
* pin br_0_238
* pin bl_0_239
* pin br_0_239
* pin bl_0_240
* pin br_0_240
* pin bl_0_241
* pin br_0_241
* pin bl_0_242
* pin br_0_242
* pin bl_0_243
* pin br_0_243
* pin bl_0_244
* pin br_0_244
* pin bl_0_245
* pin br_0_245
* pin bl_0_246
* pin br_0_246
* pin bl_0_247
* pin br_0_247
* pin bl_0_248
* pin br_0_248
* pin bl_0_249
* pin br_0_249
* pin bl_0_250
* pin br_0_250
* pin bl_0_251
* pin br_0_251
* pin bl_0_252
* pin br_0_252
* pin bl_0_253
* pin br_0_253
* pin bl_0_254
* pin br_0_254
* pin bl_0_255
* pin br_0_255
* pin bl_0_256
* pin br_0_256
* pin wl_0_66
* pin wl_0_65
* pin wl_0_68
* pin wl_0_67
* pin wl_0_69
* pin wl_0_70
* pin wl_0_71
* pin wl_0_72
* pin wl_0_73
* pin wl_0_74
* pin wl_0_75
* pin wl_0_76
* pin wl_0_78
* pin wl_0_77
* pin wl_0_79
* pin wl_0_80
* pin wl_0_82
* pin wl_0_81
* pin wl_0_83
* pin wl_0_84
* pin wl_0_85
* pin wl_0_86
* pin wl_0_87
* pin wl_0_88
* pin wl_0_89
* pin wl_0_90
* pin wl_0_91
* pin wl_0_92
* pin wl_0_94
* pin wl_0_93
* pin wl_0_95
* pin wl_0_96
* pin wl_0_97
* pin wl_0_98
* pin wl_0_100
* pin wl_0_99
* pin wl_0_102
* pin wl_0_101
* pin wl_0_103
* pin wl_0_104
* pin wl_0_105
* pin wl_0_106
* pin wl_0_107
* pin wl_0_108
* pin wl_0_109
* pin wl_0_110
* pin wl_0_111
* pin wl_0_112
* pin wl_0_113
* pin wl_0_114
* pin wl_0_115
* pin wl_0_116
* pin wl_0_117
* pin wl_0_118
* pin wl_0_119
* pin wl_0_120
* pin wl_0_122
* pin wl_0_121
* pin wl_0_124
* pin wl_0_123
* pin wl_0_125
* pin wl_0_126
* pin wl_0_127
* pin wl_0_128
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_bitcell_array 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36
+ 37 38 39 40 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84 85 86 87 88
+ 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120 121 122 123 124 125 126 127 128 129
+ 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144 145 146 147 148
+ 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164 165 166 167
+ 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184 185 186
+ 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204 205
+ 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243
+ 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262
+ 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319
+ 320 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338
+ 339 340 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357
+ 358 359 360 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376
+ 377 378 379 380 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395
+ 396 397 398 399 400 401 402 403 404 405 406 407 408 409 410 411 412 413 414
+ 415 416 417 418 419 420 421 422 423 424 425 426 427 428 429 430 431 432 433
+ 434 435 436 437 438 439 440 441 442 443 444 445 446 447 448 449 450 451 452
+ 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468 469 470 471
+ 472 473 474 475 476 477 478 479 480 481 482 483 484 485 486 487 488 489 490
+ 491 492 493 494 495 496 497 498 499 500 501 502 503 504 505 506 507 508 509
+ 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524 525 526 527 528
+ 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544 545 546 547
+ 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564 565 566
+ 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584 585
+ 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604
+ 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623
+ 624 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642
+ 643 644 645
* net 1 wl_0_0
* net 2 wl_0_1
* net 3 wl_0_3
* net 4 wl_0_2
* net 5 wl_0_4
* net 6 wl_0_5
* net 7 wl_0_6
* net 8 wl_0_7
* net 9 wl_0_9
* net 10 wl_0_8
* net 11 wl_0_10
* net 12 wl_0_11
* net 13 wl_0_12
* net 14 wl_0_13
* net 15 wl_0_14
* net 16 wl_0_15
* net 17 wl_0_16
* net 18 wl_0_17
* net 19 wl_0_18
* net 20 wl_0_19
* net 21 wl_0_20
* net 22 wl_0_21
* net 23 wl_0_22
* net 24 wl_0_23
* net 25 wl_0_25
* net 26 wl_0_24
* net 27 wl_0_26
* net 28 wl_0_27
* net 29 wl_0_28
* net 30 wl_0_29
* net 31 wl_0_30
* net 32 wl_0_31
* net 33 wl_0_32
* net 34 wl_0_33
* net 35 wl_0_34
* net 36 wl_0_35
* net 37 wl_0_36
* net 38 wl_0_37
* net 39 wl_0_39
* net 40 wl_0_38
* net 41 wl_0_41
* net 42 wl_0_40
* net 43 wl_0_43
* net 44 wl_0_42
* net 45 wl_0_44
* net 46 wl_0_45
* net 47 wl_0_46
* net 48 wl_0_47
* net 49 wl_0_48
* net 50 wl_0_49
* net 51 wl_0_50
* net 52 wl_0_51
* net 53 wl_0_52
* net 54 wl_0_53
* net 55 wl_0_54
* net 56 wl_0_55
* net 57 wl_0_56
* net 58 wl_0_57
* net 59 wl_0_58
* net 60 wl_0_59
* net 61 wl_0_60
* net 62 wl_0_61
* net 63 wl_0_62
* net 64 wl_0_63
* net 65 bl_0_0
* net 66 br_0_0
* net 67 bl_0_1
* net 68 br_0_1
* net 69 bl_0_2
* net 70 br_0_2
* net 71 bl_0_3
* net 72 br_0_3
* net 73 bl_0_4
* net 74 br_0_4
* net 75 bl_0_5
* net 76 br_0_5
* net 77 bl_0_6
* net 78 br_0_6
* net 79 bl_0_7
* net 80 br_0_7
* net 81 bl_0_8
* net 82 br_0_8
* net 83 bl_0_9
* net 84 br_0_9
* net 85 bl_0_10
* net 86 br_0_10
* net 87 bl_0_11
* net 88 br_0_11
* net 89 bl_0_12
* net 90 br_0_12
* net 91 bl_0_13
* net 92 br_0_13
* net 93 bl_0_14
* net 94 br_0_14
* net 95 bl_0_15
* net 96 br_0_15
* net 97 bl_0_16
* net 98 br_0_16
* net 99 bl_0_17
* net 100 br_0_17
* net 101 bl_0_18
* net 102 br_0_18
* net 103 bl_0_19
* net 104 br_0_19
* net 105 bl_0_20
* net 106 br_0_20
* net 107 bl_0_21
* net 108 br_0_21
* net 109 bl_0_22
* net 110 br_0_22
* net 111 bl_0_23
* net 112 br_0_23
* net 113 bl_0_24
* net 114 br_0_24
* net 115 bl_0_25
* net 116 br_0_25
* net 117 bl_0_26
* net 118 br_0_26
* net 119 bl_0_27
* net 120 br_0_27
* net 121 bl_0_28
* net 122 br_0_28
* net 123 bl_0_29
* net 124 br_0_29
* net 125 bl_0_30
* net 126 br_0_30
* net 127 bl_0_31
* net 128 br_0_31
* net 129 bl_0_32
* net 130 br_0_32
* net 131 bl_0_33
* net 132 br_0_33
* net 133 bl_0_34
* net 134 br_0_34
* net 135 bl_0_35
* net 136 br_0_35
* net 137 bl_0_36
* net 138 br_0_36
* net 139 bl_0_37
* net 140 br_0_37
* net 141 bl_0_38
* net 142 br_0_38
* net 143 bl_0_39
* net 144 br_0_39
* net 145 bl_0_40
* net 146 br_0_40
* net 147 bl_0_41
* net 148 br_0_41
* net 149 bl_0_42
* net 150 br_0_42
* net 151 bl_0_43
* net 152 br_0_43
* net 153 bl_0_44
* net 154 br_0_44
* net 155 bl_0_45
* net 156 br_0_45
* net 157 bl_0_46
* net 158 br_0_46
* net 159 bl_0_47
* net 160 br_0_47
* net 161 bl_0_48
* net 162 br_0_48
* net 163 bl_0_49
* net 164 br_0_49
* net 165 bl_0_50
* net 166 br_0_50
* net 167 bl_0_51
* net 168 br_0_51
* net 169 bl_0_52
* net 170 br_0_52
* net 171 bl_0_53
* net 172 br_0_53
* net 173 bl_0_54
* net 174 br_0_54
* net 175 bl_0_55
* net 176 br_0_55
* net 177 bl_0_56
* net 178 br_0_56
* net 179 bl_0_57
* net 180 br_0_57
* net 181 bl_0_58
* net 182 br_0_58
* net 183 bl_0_59
* net 184 br_0_59
* net 185 bl_0_60
* net 186 br_0_60
* net 187 bl_0_61
* net 188 br_0_61
* net 189 bl_0_62
* net 190 br_0_62
* net 191 bl_0_63
* net 192 br_0_63
* net 193 bl_0_64
* net 194 br_0_64
* net 195 bl_0_65
* net 196 br_0_65
* net 197 bl_0_66
* net 198 br_0_66
* net 199 bl_0_67
* net 200 br_0_67
* net 201 bl_0_68
* net 202 br_0_68
* net 203 bl_0_69
* net 204 br_0_69
* net 205 bl_0_70
* net 206 br_0_70
* net 207 bl_0_71
* net 208 br_0_71
* net 209 bl_0_72
* net 210 br_0_72
* net 211 bl_0_73
* net 212 br_0_73
* net 213 bl_0_74
* net 214 br_0_74
* net 215 bl_0_75
* net 216 br_0_75
* net 217 bl_0_76
* net 218 br_0_76
* net 219 bl_0_77
* net 220 br_0_77
* net 221 bl_0_78
* net 222 br_0_78
* net 223 bl_0_79
* net 224 br_0_79
* net 225 bl_0_80
* net 226 br_0_80
* net 227 bl_0_81
* net 228 br_0_81
* net 229 bl_0_82
* net 230 br_0_82
* net 231 bl_0_83
* net 232 br_0_83
* net 233 bl_0_84
* net 234 br_0_84
* net 235 bl_0_85
* net 236 br_0_85
* net 237 bl_0_86
* net 238 br_0_86
* net 239 bl_0_87
* net 240 br_0_87
* net 241 bl_0_88
* net 242 br_0_88
* net 243 bl_0_89
* net 244 br_0_89
* net 245 bl_0_90
* net 246 br_0_90
* net 247 bl_0_91
* net 248 br_0_91
* net 249 bl_0_92
* net 250 br_0_92
* net 251 bl_0_93
* net 252 br_0_93
* net 253 bl_0_94
* net 254 br_0_94
* net 255 bl_0_95
* net 256 br_0_95
* net 257 bl_0_96
* net 258 br_0_96
* net 259 bl_0_97
* net 260 br_0_97
* net 261 bl_0_98
* net 262 br_0_98
* net 263 bl_0_99
* net 264 br_0_99
* net 265 bl_0_100
* net 266 br_0_100
* net 267 bl_0_101
* net 268 br_0_101
* net 269 bl_0_102
* net 270 br_0_102
* net 271 bl_0_103
* net 272 br_0_103
* net 273 bl_0_104
* net 274 br_0_104
* net 275 bl_0_105
* net 276 br_0_105
* net 277 bl_0_106
* net 278 br_0_106
* net 279 bl_0_107
* net 280 br_0_107
* net 281 bl_0_108
* net 282 br_0_108
* net 283 bl_0_109
* net 284 br_0_109
* net 285 bl_0_110
* net 286 br_0_110
* net 287 bl_0_111
* net 288 br_0_111
* net 289 bl_0_112
* net 290 br_0_112
* net 291 bl_0_113
* net 292 br_0_113
* net 293 bl_0_114
* net 294 br_0_114
* net 295 bl_0_115
* net 296 br_0_115
* net 297 bl_0_116
* net 298 br_0_116
* net 299 bl_0_117
* net 300 br_0_117
* net 301 bl_0_118
* net 302 br_0_118
* net 303 bl_0_119
* net 304 br_0_119
* net 305 bl_0_120
* net 306 br_0_120
* net 307 bl_0_121
* net 308 br_0_121
* net 309 bl_0_122
* net 310 br_0_122
* net 311 bl_0_123
* net 312 br_0_123
* net 313 bl_0_124
* net 314 br_0_124
* net 315 bl_0_125
* net 316 br_0_125
* net 317 bl_0_126
* net 318 br_0_126
* net 319 bl_0_127
* net 320 br_0_127
* net 321 bl_0_128
* net 322 wl_0_64
* net 323 br_0_128
* net 324 bl_0_129
* net 325 br_0_129
* net 326 bl_0_130
* net 327 br_0_130
* net 328 bl_0_131
* net 329 br_0_131
* net 330 bl_0_132
* net 331 br_0_132
* net 332 bl_0_133
* net 333 br_0_133
* net 334 bl_0_134
* net 335 br_0_134
* net 336 bl_0_135
* net 337 br_0_135
* net 338 bl_0_136
* net 339 br_0_136
* net 340 bl_0_137
* net 341 br_0_137
* net 342 bl_0_138
* net 343 br_0_138
* net 344 bl_0_139
* net 345 br_0_139
* net 346 bl_0_140
* net 347 br_0_140
* net 348 bl_0_141
* net 349 br_0_141
* net 350 bl_0_142
* net 351 br_0_142
* net 352 bl_0_143
* net 353 br_0_143
* net 354 bl_0_144
* net 355 br_0_144
* net 356 bl_0_145
* net 357 br_0_145
* net 358 bl_0_146
* net 359 br_0_146
* net 360 bl_0_147
* net 361 br_0_147
* net 362 bl_0_148
* net 363 br_0_148
* net 364 bl_0_149
* net 365 br_0_149
* net 366 bl_0_150
* net 367 br_0_150
* net 368 bl_0_151
* net 369 br_0_151
* net 370 bl_0_152
* net 371 br_0_152
* net 372 bl_0_153
* net 373 br_0_153
* net 374 bl_0_154
* net 375 br_0_154
* net 376 bl_0_155
* net 377 br_0_155
* net 378 bl_0_156
* net 379 br_0_156
* net 380 bl_0_157
* net 381 br_0_157
* net 382 bl_0_158
* net 383 br_0_158
* net 384 bl_0_159
* net 385 br_0_159
* net 386 bl_0_160
* net 387 br_0_160
* net 388 bl_0_161
* net 389 br_0_161
* net 390 bl_0_162
* net 391 br_0_162
* net 392 bl_0_163
* net 393 br_0_163
* net 394 bl_0_164
* net 395 br_0_164
* net 396 bl_0_165
* net 397 br_0_165
* net 398 bl_0_166
* net 399 br_0_166
* net 400 bl_0_167
* net 401 br_0_167
* net 402 bl_0_168
* net 403 br_0_168
* net 404 bl_0_169
* net 405 br_0_169
* net 406 bl_0_170
* net 407 br_0_170
* net 408 bl_0_171
* net 409 br_0_171
* net 410 bl_0_172
* net 411 br_0_172
* net 412 bl_0_173
* net 413 br_0_173
* net 414 bl_0_174
* net 415 br_0_174
* net 416 bl_0_175
* net 417 br_0_175
* net 418 bl_0_176
* net 419 br_0_176
* net 420 bl_0_177
* net 421 br_0_177
* net 422 bl_0_178
* net 423 br_0_178
* net 424 bl_0_179
* net 425 br_0_179
* net 426 bl_0_180
* net 427 br_0_180
* net 428 bl_0_181
* net 429 br_0_181
* net 430 bl_0_182
* net 431 br_0_182
* net 432 bl_0_183
* net 433 br_0_183
* net 434 bl_0_184
* net 435 br_0_184
* net 436 bl_0_185
* net 437 br_0_185
* net 438 bl_0_186
* net 439 br_0_186
* net 440 bl_0_187
* net 441 br_0_187
* net 442 bl_0_188
* net 443 br_0_188
* net 444 bl_0_189
* net 445 br_0_189
* net 446 bl_0_190
* net 447 br_0_190
* net 448 bl_0_191
* net 449 br_0_191
* net 450 bl_0_192
* net 451 br_0_192
* net 452 bl_0_193
* net 453 br_0_193
* net 454 bl_0_194
* net 455 br_0_194
* net 456 bl_0_195
* net 457 br_0_195
* net 458 bl_0_196
* net 459 br_0_196
* net 460 bl_0_197
* net 461 br_0_197
* net 462 bl_0_198
* net 463 br_0_198
* net 464 bl_0_199
* net 465 br_0_199
* net 466 bl_0_200
* net 467 br_0_200
* net 468 bl_0_201
* net 469 br_0_201
* net 470 bl_0_202
* net 471 br_0_202
* net 472 bl_0_203
* net 473 br_0_203
* net 474 bl_0_204
* net 475 br_0_204
* net 476 bl_0_205
* net 477 br_0_205
* net 478 bl_0_206
* net 479 br_0_206
* net 480 bl_0_207
* net 481 br_0_207
* net 482 bl_0_208
* net 483 br_0_208
* net 484 bl_0_209
* net 485 br_0_209
* net 486 bl_0_210
* net 487 br_0_210
* net 488 bl_0_211
* net 489 br_0_211
* net 490 bl_0_212
* net 491 br_0_212
* net 492 bl_0_213
* net 493 br_0_213
* net 494 bl_0_214
* net 495 br_0_214
* net 496 bl_0_215
* net 497 br_0_215
* net 498 bl_0_216
* net 499 br_0_216
* net 500 bl_0_217
* net 501 br_0_217
* net 502 bl_0_218
* net 503 br_0_218
* net 504 bl_0_219
* net 505 br_0_219
* net 506 bl_0_220
* net 507 br_0_220
* net 508 bl_0_221
* net 509 br_0_221
* net 510 bl_0_222
* net 511 br_0_222
* net 512 bl_0_223
* net 513 br_0_223
* net 514 bl_0_224
* net 515 br_0_224
* net 516 bl_0_225
* net 517 br_0_225
* net 518 bl_0_226
* net 519 br_0_226
* net 520 bl_0_227
* net 521 br_0_227
* net 522 bl_0_228
* net 523 br_0_228
* net 524 bl_0_229
* net 525 br_0_229
* net 526 bl_0_230
* net 527 br_0_230
* net 528 bl_0_231
* net 529 br_0_231
* net 530 bl_0_232
* net 531 br_0_232
* net 532 bl_0_233
* net 533 br_0_233
* net 534 bl_0_234
* net 535 br_0_234
* net 536 bl_0_235
* net 537 br_0_235
* net 538 bl_0_236
* net 539 br_0_236
* net 540 bl_0_237
* net 541 br_0_237
* net 542 bl_0_238
* net 543 br_0_238
* net 544 bl_0_239
* net 545 br_0_239
* net 546 bl_0_240
* net 547 br_0_240
* net 548 bl_0_241
* net 549 br_0_241
* net 550 bl_0_242
* net 551 br_0_242
* net 552 bl_0_243
* net 553 br_0_243
* net 554 bl_0_244
* net 555 br_0_244
* net 556 bl_0_245
* net 557 br_0_245
* net 558 bl_0_246
* net 559 br_0_246
* net 560 bl_0_247
* net 561 br_0_247
* net 562 bl_0_248
* net 563 br_0_248
* net 564 bl_0_249
* net 565 br_0_249
* net 566 bl_0_250
* net 567 br_0_250
* net 568 bl_0_251
* net 569 br_0_251
* net 570 bl_0_252
* net 571 br_0_252
* net 572 bl_0_253
* net 573 br_0_253
* net 574 bl_0_254
* net 575 br_0_254
* net 576 bl_0_255
* net 577 br_0_255
* net 578 bl_0_256
* net 579 br_0_256
* net 580 wl_0_66
* net 581 wl_0_65
* net 582 wl_0_68
* net 583 wl_0_67
* net 584 wl_0_69
* net 585 wl_0_70
* net 586 wl_0_71
* net 587 wl_0_72
* net 588 wl_0_73
* net 589 wl_0_74
* net 590 wl_0_75
* net 591 wl_0_76
* net 592 wl_0_78
* net 593 wl_0_77
* net 594 wl_0_79
* net 595 wl_0_80
* net 596 wl_0_82
* net 597 wl_0_81
* net 598 wl_0_83
* net 599 wl_0_84
* net 600 wl_0_85
* net 601 wl_0_86
* net 602 wl_0_87
* net 603 wl_0_88
* net 604 wl_0_89
* net 605 wl_0_90
* net 606 wl_0_91
* net 607 wl_0_92
* net 608 wl_0_94
* net 609 wl_0_93
* net 610 wl_0_95
* net 611 wl_0_96
* net 612 wl_0_97
* net 613 wl_0_98
* net 614 wl_0_100
* net 615 wl_0_99
* net 616 wl_0_102
* net 617 wl_0_101
* net 618 wl_0_103
* net 619 wl_0_104
* net 620 wl_0_105
* net 621 wl_0_106
* net 622 wl_0_107
* net 623 wl_0_108
* net 624 wl_0_109
* net 625 wl_0_110
* net 626 wl_0_111
* net 627 wl_0_112
* net 628 wl_0_113
* net 629 wl_0_114
* net 630 wl_0_115
* net 631 wl_0_116
* net 632 wl_0_117
* net 633 wl_0_118
* net 634 wl_0_119
* net 635 wl_0_120
* net 636 wl_0_122
* net 637 wl_0_121
* net 638 wl_0_124
* net 639 wl_0_123
* net 640 wl_0_125
* net 641 wl_0_126
* net 642 wl_0_127
* net 643 wl_0_128
* net 644 vdd
* net 645 gnd
* cell instance $1 r0 *1 0,0
X$1 65 1 66 644 645 cell_1rw
* cell instance $2 r0 *1 0.705,0
X$2 67 1 68 644 645 cell_1rw
* cell instance $3 r0 *1 1.41,0
X$3 69 1 70 644 645 cell_1rw
* cell instance $4 r0 *1 2.115,0
X$4 71 1 72 644 645 cell_1rw
* cell instance $5 r0 *1 2.82,0
X$5 73 1 74 644 645 cell_1rw
* cell instance $6 r0 *1 3.525,0
X$6 75 1 76 644 645 cell_1rw
* cell instance $7 r0 *1 4.23,0
X$7 77 1 78 644 645 cell_1rw
* cell instance $8 r0 *1 4.935,0
X$8 79 1 80 644 645 cell_1rw
* cell instance $9 r0 *1 5.64,0
X$9 81 1 82 644 645 cell_1rw
* cell instance $10 r0 *1 6.345,0
X$10 83 1 84 644 645 cell_1rw
* cell instance $11 r0 *1 7.05,0
X$11 85 1 86 644 645 cell_1rw
* cell instance $12 r0 *1 7.755,0
X$12 87 1 88 644 645 cell_1rw
* cell instance $13 r0 *1 8.46,0
X$13 89 1 90 644 645 cell_1rw
* cell instance $14 r0 *1 9.165,0
X$14 91 1 92 644 645 cell_1rw
* cell instance $15 r0 *1 9.87,0
X$15 93 1 94 644 645 cell_1rw
* cell instance $16 r0 *1 10.575,0
X$16 95 1 96 644 645 cell_1rw
* cell instance $17 r0 *1 11.28,0
X$17 97 1 98 644 645 cell_1rw
* cell instance $18 r0 *1 11.985,0
X$18 99 1 100 644 645 cell_1rw
* cell instance $19 r0 *1 12.69,0
X$19 101 1 102 644 645 cell_1rw
* cell instance $20 r0 *1 13.395,0
X$20 103 1 104 644 645 cell_1rw
* cell instance $21 r0 *1 14.1,0
X$21 105 1 106 644 645 cell_1rw
* cell instance $22 r0 *1 14.805,0
X$22 107 1 108 644 645 cell_1rw
* cell instance $23 r0 *1 15.51,0
X$23 109 1 110 644 645 cell_1rw
* cell instance $24 r0 *1 16.215,0
X$24 111 1 112 644 645 cell_1rw
* cell instance $25 r0 *1 16.92,0
X$25 113 1 114 644 645 cell_1rw
* cell instance $26 r0 *1 17.625,0
X$26 115 1 116 644 645 cell_1rw
* cell instance $27 r0 *1 18.33,0
X$27 117 1 118 644 645 cell_1rw
* cell instance $28 r0 *1 19.035,0
X$28 119 1 120 644 645 cell_1rw
* cell instance $29 r0 *1 19.74,0
X$29 121 1 122 644 645 cell_1rw
* cell instance $30 r0 *1 20.445,0
X$30 123 1 124 644 645 cell_1rw
* cell instance $31 r0 *1 21.15,0
X$31 125 1 126 644 645 cell_1rw
* cell instance $32 r0 *1 21.855,0
X$32 127 1 128 644 645 cell_1rw
* cell instance $33 r0 *1 22.56,0
X$33 129 1 130 644 645 cell_1rw
* cell instance $34 r0 *1 23.265,0
X$34 131 1 132 644 645 cell_1rw
* cell instance $35 r0 *1 23.97,0
X$35 133 1 134 644 645 cell_1rw
* cell instance $36 r0 *1 24.675,0
X$36 135 1 136 644 645 cell_1rw
* cell instance $37 r0 *1 25.38,0
X$37 137 1 138 644 645 cell_1rw
* cell instance $38 r0 *1 26.085,0
X$38 139 1 140 644 645 cell_1rw
* cell instance $39 r0 *1 26.79,0
X$39 141 1 142 644 645 cell_1rw
* cell instance $40 r0 *1 27.495,0
X$40 143 1 144 644 645 cell_1rw
* cell instance $41 r0 *1 28.2,0
X$41 145 1 146 644 645 cell_1rw
* cell instance $42 r0 *1 28.905,0
X$42 147 1 148 644 645 cell_1rw
* cell instance $43 r0 *1 29.61,0
X$43 149 1 150 644 645 cell_1rw
* cell instance $44 r0 *1 30.315,0
X$44 151 1 152 644 645 cell_1rw
* cell instance $45 r0 *1 31.02,0
X$45 153 1 154 644 645 cell_1rw
* cell instance $46 r0 *1 31.725,0
X$46 155 1 156 644 645 cell_1rw
* cell instance $47 r0 *1 32.43,0
X$47 157 1 158 644 645 cell_1rw
* cell instance $48 r0 *1 33.135,0
X$48 159 1 160 644 645 cell_1rw
* cell instance $49 r0 *1 33.84,0
X$49 161 1 162 644 645 cell_1rw
* cell instance $50 r0 *1 34.545,0
X$50 163 1 164 644 645 cell_1rw
* cell instance $51 r0 *1 35.25,0
X$51 165 1 166 644 645 cell_1rw
* cell instance $52 r0 *1 35.955,0
X$52 167 1 168 644 645 cell_1rw
* cell instance $53 r0 *1 36.66,0
X$53 169 1 170 644 645 cell_1rw
* cell instance $54 r0 *1 37.365,0
X$54 171 1 172 644 645 cell_1rw
* cell instance $55 r0 *1 38.07,0
X$55 173 1 174 644 645 cell_1rw
* cell instance $56 r0 *1 38.775,0
X$56 175 1 176 644 645 cell_1rw
* cell instance $57 r0 *1 39.48,0
X$57 177 1 178 644 645 cell_1rw
* cell instance $58 r0 *1 40.185,0
X$58 179 1 180 644 645 cell_1rw
* cell instance $59 r0 *1 40.89,0
X$59 181 1 182 644 645 cell_1rw
* cell instance $60 r0 *1 41.595,0
X$60 183 1 184 644 645 cell_1rw
* cell instance $61 r0 *1 42.3,0
X$61 185 1 186 644 645 cell_1rw
* cell instance $62 r0 *1 43.005,0
X$62 187 1 188 644 645 cell_1rw
* cell instance $63 r0 *1 43.71,0
X$63 189 1 190 644 645 cell_1rw
* cell instance $64 r0 *1 44.415,0
X$64 191 1 192 644 645 cell_1rw
* cell instance $65 r0 *1 45.12,0
X$65 193 1 194 644 645 cell_1rw
* cell instance $66 r0 *1 45.825,0
X$66 195 1 196 644 645 cell_1rw
* cell instance $67 r0 *1 46.53,0
X$67 197 1 198 644 645 cell_1rw
* cell instance $68 r0 *1 47.235,0
X$68 199 1 200 644 645 cell_1rw
* cell instance $69 r0 *1 47.94,0
X$69 201 1 202 644 645 cell_1rw
* cell instance $70 r0 *1 48.645,0
X$70 203 1 204 644 645 cell_1rw
* cell instance $71 r0 *1 49.35,0
X$71 205 1 206 644 645 cell_1rw
* cell instance $72 r0 *1 50.055,0
X$72 207 1 208 644 645 cell_1rw
* cell instance $73 r0 *1 50.76,0
X$73 209 1 210 644 645 cell_1rw
* cell instance $74 r0 *1 51.465,0
X$74 211 1 212 644 645 cell_1rw
* cell instance $75 r0 *1 52.17,0
X$75 213 1 214 644 645 cell_1rw
* cell instance $76 r0 *1 52.875,0
X$76 215 1 216 644 645 cell_1rw
* cell instance $77 r0 *1 53.58,0
X$77 217 1 218 644 645 cell_1rw
* cell instance $78 r0 *1 54.285,0
X$78 219 1 220 644 645 cell_1rw
* cell instance $79 r0 *1 54.99,0
X$79 221 1 222 644 645 cell_1rw
* cell instance $80 r0 *1 55.695,0
X$80 223 1 224 644 645 cell_1rw
* cell instance $81 r0 *1 56.4,0
X$81 225 1 226 644 645 cell_1rw
* cell instance $82 r0 *1 57.105,0
X$82 227 1 228 644 645 cell_1rw
* cell instance $83 r0 *1 57.81,0
X$83 229 1 230 644 645 cell_1rw
* cell instance $84 r0 *1 58.515,0
X$84 231 1 232 644 645 cell_1rw
* cell instance $85 r0 *1 59.22,0
X$85 233 1 234 644 645 cell_1rw
* cell instance $86 r0 *1 59.925,0
X$86 235 1 236 644 645 cell_1rw
* cell instance $87 r0 *1 60.63,0
X$87 237 1 238 644 645 cell_1rw
* cell instance $88 r0 *1 61.335,0
X$88 239 1 240 644 645 cell_1rw
* cell instance $89 r0 *1 62.04,0
X$89 241 1 242 644 645 cell_1rw
* cell instance $90 r0 *1 62.745,0
X$90 243 1 244 644 645 cell_1rw
* cell instance $91 r0 *1 63.45,0
X$91 245 1 246 644 645 cell_1rw
* cell instance $92 r0 *1 64.155,0
X$92 247 1 248 644 645 cell_1rw
* cell instance $93 r0 *1 64.86,0
X$93 249 1 250 644 645 cell_1rw
* cell instance $94 r0 *1 65.565,0
X$94 251 1 252 644 645 cell_1rw
* cell instance $95 r0 *1 66.27,0
X$95 253 1 254 644 645 cell_1rw
* cell instance $96 r0 *1 66.975,0
X$96 255 1 256 644 645 cell_1rw
* cell instance $97 r0 *1 67.68,0
X$97 257 1 258 644 645 cell_1rw
* cell instance $98 r0 *1 68.385,0
X$98 259 1 260 644 645 cell_1rw
* cell instance $99 r0 *1 69.09,0
X$99 261 1 262 644 645 cell_1rw
* cell instance $100 r0 *1 69.795,0
X$100 263 1 264 644 645 cell_1rw
* cell instance $101 r0 *1 70.5,0
X$101 265 1 266 644 645 cell_1rw
* cell instance $102 r0 *1 71.205,0
X$102 267 1 268 644 645 cell_1rw
* cell instance $103 r0 *1 71.91,0
X$103 269 1 270 644 645 cell_1rw
* cell instance $104 r0 *1 72.615,0
X$104 271 1 272 644 645 cell_1rw
* cell instance $105 r0 *1 73.32,0
X$105 273 1 274 644 645 cell_1rw
* cell instance $106 r0 *1 74.025,0
X$106 275 1 276 644 645 cell_1rw
* cell instance $107 r0 *1 74.73,0
X$107 277 1 278 644 645 cell_1rw
* cell instance $108 r0 *1 75.435,0
X$108 279 1 280 644 645 cell_1rw
* cell instance $109 r0 *1 76.14,0
X$109 281 1 282 644 645 cell_1rw
* cell instance $110 r0 *1 76.845,0
X$110 283 1 284 644 645 cell_1rw
* cell instance $111 r0 *1 77.55,0
X$111 285 1 286 644 645 cell_1rw
* cell instance $112 r0 *1 78.255,0
X$112 287 1 288 644 645 cell_1rw
* cell instance $113 r0 *1 78.96,0
X$113 289 1 290 644 645 cell_1rw
* cell instance $114 r0 *1 79.665,0
X$114 291 1 292 644 645 cell_1rw
* cell instance $115 r0 *1 80.37,0
X$115 293 1 294 644 645 cell_1rw
* cell instance $116 r0 *1 81.075,0
X$116 295 1 296 644 645 cell_1rw
* cell instance $117 r0 *1 81.78,0
X$117 297 1 298 644 645 cell_1rw
* cell instance $118 r0 *1 82.485,0
X$118 299 1 300 644 645 cell_1rw
* cell instance $119 r0 *1 83.19,0
X$119 301 1 302 644 645 cell_1rw
* cell instance $120 r0 *1 83.895,0
X$120 303 1 304 644 645 cell_1rw
* cell instance $121 r0 *1 84.6,0
X$121 305 1 306 644 645 cell_1rw
* cell instance $122 r0 *1 85.305,0
X$122 307 1 308 644 645 cell_1rw
* cell instance $123 r0 *1 86.01,0
X$123 309 1 310 644 645 cell_1rw
* cell instance $124 r0 *1 86.715,0
X$124 311 1 312 644 645 cell_1rw
* cell instance $125 r0 *1 87.42,0
X$125 313 1 314 644 645 cell_1rw
* cell instance $126 r0 *1 88.125,0
X$126 315 1 316 644 645 cell_1rw
* cell instance $127 r0 *1 88.83,0
X$127 317 1 318 644 645 cell_1rw
* cell instance $128 r0 *1 89.535,0
X$128 319 1 320 644 645 cell_1rw
* cell instance $129 r0 *1 90.24,0
X$129 321 1 323 644 645 cell_1rw
* cell instance $130 r0 *1 90.945,0
X$130 324 1 325 644 645 cell_1rw
* cell instance $131 r0 *1 91.65,0
X$131 326 1 327 644 645 cell_1rw
* cell instance $132 r0 *1 92.355,0
X$132 328 1 329 644 645 cell_1rw
* cell instance $133 r0 *1 93.06,0
X$133 330 1 331 644 645 cell_1rw
* cell instance $134 r0 *1 93.765,0
X$134 332 1 333 644 645 cell_1rw
* cell instance $135 r0 *1 94.47,0
X$135 334 1 335 644 645 cell_1rw
* cell instance $136 r0 *1 95.175,0
X$136 336 1 337 644 645 cell_1rw
* cell instance $137 r0 *1 95.88,0
X$137 338 1 339 644 645 cell_1rw
* cell instance $138 r0 *1 96.585,0
X$138 340 1 341 644 645 cell_1rw
* cell instance $139 r0 *1 97.29,0
X$139 342 1 343 644 645 cell_1rw
* cell instance $140 r0 *1 97.995,0
X$140 344 1 345 644 645 cell_1rw
* cell instance $141 r0 *1 98.7,0
X$141 346 1 347 644 645 cell_1rw
* cell instance $142 r0 *1 99.405,0
X$142 348 1 349 644 645 cell_1rw
* cell instance $143 r0 *1 100.11,0
X$143 350 1 351 644 645 cell_1rw
* cell instance $144 r0 *1 100.815,0
X$144 352 1 353 644 645 cell_1rw
* cell instance $145 r0 *1 101.52,0
X$145 354 1 355 644 645 cell_1rw
* cell instance $146 r0 *1 102.225,0
X$146 356 1 357 644 645 cell_1rw
* cell instance $147 r0 *1 102.93,0
X$147 358 1 359 644 645 cell_1rw
* cell instance $148 r0 *1 103.635,0
X$148 360 1 361 644 645 cell_1rw
* cell instance $149 r0 *1 104.34,0
X$149 362 1 363 644 645 cell_1rw
* cell instance $150 r0 *1 105.045,0
X$150 364 1 365 644 645 cell_1rw
* cell instance $151 r0 *1 105.75,0
X$151 366 1 367 644 645 cell_1rw
* cell instance $152 r0 *1 106.455,0
X$152 368 1 369 644 645 cell_1rw
* cell instance $153 r0 *1 107.16,0
X$153 370 1 371 644 645 cell_1rw
* cell instance $154 r0 *1 107.865,0
X$154 372 1 373 644 645 cell_1rw
* cell instance $155 r0 *1 108.57,0
X$155 374 1 375 644 645 cell_1rw
* cell instance $156 r0 *1 109.275,0
X$156 376 1 377 644 645 cell_1rw
* cell instance $157 r0 *1 109.98,0
X$157 378 1 379 644 645 cell_1rw
* cell instance $158 r0 *1 110.685,0
X$158 380 1 381 644 645 cell_1rw
* cell instance $159 r0 *1 111.39,0
X$159 382 1 383 644 645 cell_1rw
* cell instance $160 r0 *1 112.095,0
X$160 384 1 385 644 645 cell_1rw
* cell instance $161 r0 *1 112.8,0
X$161 386 1 387 644 645 cell_1rw
* cell instance $162 r0 *1 113.505,0
X$162 388 1 389 644 645 cell_1rw
* cell instance $163 r0 *1 114.21,0
X$163 390 1 391 644 645 cell_1rw
* cell instance $164 r0 *1 114.915,0
X$164 392 1 393 644 645 cell_1rw
* cell instance $165 r0 *1 115.62,0
X$165 394 1 395 644 645 cell_1rw
* cell instance $166 r0 *1 116.325,0
X$166 396 1 397 644 645 cell_1rw
* cell instance $167 r0 *1 117.03,0
X$167 398 1 399 644 645 cell_1rw
* cell instance $168 r0 *1 117.735,0
X$168 400 1 401 644 645 cell_1rw
* cell instance $169 r0 *1 118.44,0
X$169 402 1 403 644 645 cell_1rw
* cell instance $170 r0 *1 119.145,0
X$170 404 1 405 644 645 cell_1rw
* cell instance $171 r0 *1 119.85,0
X$171 406 1 407 644 645 cell_1rw
* cell instance $172 r0 *1 120.555,0
X$172 408 1 409 644 645 cell_1rw
* cell instance $173 r0 *1 121.26,0
X$173 410 1 411 644 645 cell_1rw
* cell instance $174 r0 *1 121.965,0
X$174 412 1 413 644 645 cell_1rw
* cell instance $175 r0 *1 122.67,0
X$175 414 1 415 644 645 cell_1rw
* cell instance $176 r0 *1 123.375,0
X$176 416 1 417 644 645 cell_1rw
* cell instance $177 r0 *1 124.08,0
X$177 418 1 419 644 645 cell_1rw
* cell instance $178 r0 *1 124.785,0
X$178 420 1 421 644 645 cell_1rw
* cell instance $179 r0 *1 125.49,0
X$179 422 1 423 644 645 cell_1rw
* cell instance $180 r0 *1 126.195,0
X$180 424 1 425 644 645 cell_1rw
* cell instance $181 r0 *1 126.9,0
X$181 426 1 427 644 645 cell_1rw
* cell instance $182 r0 *1 127.605,0
X$182 428 1 429 644 645 cell_1rw
* cell instance $183 r0 *1 128.31,0
X$183 430 1 431 644 645 cell_1rw
* cell instance $184 r0 *1 129.015,0
X$184 432 1 433 644 645 cell_1rw
* cell instance $185 r0 *1 129.72,0
X$185 434 1 435 644 645 cell_1rw
* cell instance $186 r0 *1 130.425,0
X$186 436 1 437 644 645 cell_1rw
* cell instance $187 r0 *1 131.13,0
X$187 438 1 439 644 645 cell_1rw
* cell instance $188 r0 *1 131.835,0
X$188 440 1 441 644 645 cell_1rw
* cell instance $189 r0 *1 132.54,0
X$189 442 1 443 644 645 cell_1rw
* cell instance $190 r0 *1 133.245,0
X$190 444 1 445 644 645 cell_1rw
* cell instance $191 r0 *1 133.95,0
X$191 446 1 447 644 645 cell_1rw
* cell instance $192 r0 *1 134.655,0
X$192 448 1 449 644 645 cell_1rw
* cell instance $193 r0 *1 135.36,0
X$193 450 1 451 644 645 cell_1rw
* cell instance $194 r0 *1 136.065,0
X$194 452 1 453 644 645 cell_1rw
* cell instance $195 r0 *1 136.77,0
X$195 454 1 455 644 645 cell_1rw
* cell instance $196 r0 *1 137.475,0
X$196 456 1 457 644 645 cell_1rw
* cell instance $197 r0 *1 138.18,0
X$197 458 1 459 644 645 cell_1rw
* cell instance $198 r0 *1 138.885,0
X$198 460 1 461 644 645 cell_1rw
* cell instance $199 r0 *1 139.59,0
X$199 462 1 463 644 645 cell_1rw
* cell instance $200 r0 *1 140.295,0
X$200 464 1 465 644 645 cell_1rw
* cell instance $201 r0 *1 141,0
X$201 466 1 467 644 645 cell_1rw
* cell instance $202 r0 *1 141.705,0
X$202 468 1 469 644 645 cell_1rw
* cell instance $203 r0 *1 142.41,0
X$203 470 1 471 644 645 cell_1rw
* cell instance $204 r0 *1 143.115,0
X$204 472 1 473 644 645 cell_1rw
* cell instance $205 r0 *1 143.82,0
X$205 474 1 475 644 645 cell_1rw
* cell instance $206 r0 *1 144.525,0
X$206 476 1 477 644 645 cell_1rw
* cell instance $207 r0 *1 145.23,0
X$207 478 1 479 644 645 cell_1rw
* cell instance $208 r0 *1 145.935,0
X$208 480 1 481 644 645 cell_1rw
* cell instance $209 r0 *1 146.64,0
X$209 482 1 483 644 645 cell_1rw
* cell instance $210 r0 *1 147.345,0
X$210 484 1 485 644 645 cell_1rw
* cell instance $211 r0 *1 148.05,0
X$211 486 1 487 644 645 cell_1rw
* cell instance $212 r0 *1 148.755,0
X$212 488 1 489 644 645 cell_1rw
* cell instance $213 r0 *1 149.46,0
X$213 490 1 491 644 645 cell_1rw
* cell instance $214 r0 *1 150.165,0
X$214 492 1 493 644 645 cell_1rw
* cell instance $215 r0 *1 150.87,0
X$215 494 1 495 644 645 cell_1rw
* cell instance $216 r0 *1 151.575,0
X$216 496 1 497 644 645 cell_1rw
* cell instance $217 r0 *1 152.28,0
X$217 498 1 499 644 645 cell_1rw
* cell instance $218 r0 *1 152.985,0
X$218 500 1 501 644 645 cell_1rw
* cell instance $219 r0 *1 153.69,0
X$219 502 1 503 644 645 cell_1rw
* cell instance $220 r0 *1 154.395,0
X$220 504 1 505 644 645 cell_1rw
* cell instance $221 r0 *1 155.1,0
X$221 506 1 507 644 645 cell_1rw
* cell instance $222 r0 *1 155.805,0
X$222 508 1 509 644 645 cell_1rw
* cell instance $223 r0 *1 156.51,0
X$223 510 1 511 644 645 cell_1rw
* cell instance $224 r0 *1 157.215,0
X$224 512 1 513 644 645 cell_1rw
* cell instance $225 r0 *1 157.92,0
X$225 514 1 515 644 645 cell_1rw
* cell instance $226 r0 *1 158.625,0
X$226 516 1 517 644 645 cell_1rw
* cell instance $227 r0 *1 159.33,0
X$227 518 1 519 644 645 cell_1rw
* cell instance $228 r0 *1 160.035,0
X$228 520 1 521 644 645 cell_1rw
* cell instance $229 r0 *1 160.74,0
X$229 522 1 523 644 645 cell_1rw
* cell instance $230 r0 *1 161.445,0
X$230 524 1 525 644 645 cell_1rw
* cell instance $231 r0 *1 162.15,0
X$231 526 1 527 644 645 cell_1rw
* cell instance $232 r0 *1 162.855,0
X$232 528 1 529 644 645 cell_1rw
* cell instance $233 r0 *1 163.56,0
X$233 530 1 531 644 645 cell_1rw
* cell instance $234 r0 *1 164.265,0
X$234 532 1 533 644 645 cell_1rw
* cell instance $235 r0 *1 164.97,0
X$235 534 1 535 644 645 cell_1rw
* cell instance $236 r0 *1 165.675,0
X$236 536 1 537 644 645 cell_1rw
* cell instance $237 r0 *1 166.38,0
X$237 538 1 539 644 645 cell_1rw
* cell instance $238 r0 *1 167.085,0
X$238 540 1 541 644 645 cell_1rw
* cell instance $239 r0 *1 167.79,0
X$239 542 1 543 644 645 cell_1rw
* cell instance $240 r0 *1 168.495,0
X$240 544 1 545 644 645 cell_1rw
* cell instance $241 r0 *1 169.2,0
X$241 546 1 547 644 645 cell_1rw
* cell instance $242 r0 *1 169.905,0
X$242 548 1 549 644 645 cell_1rw
* cell instance $243 r0 *1 170.61,0
X$243 550 1 551 644 645 cell_1rw
* cell instance $244 r0 *1 171.315,0
X$244 552 1 553 644 645 cell_1rw
* cell instance $245 r0 *1 172.02,0
X$245 554 1 555 644 645 cell_1rw
* cell instance $246 r0 *1 172.725,0
X$246 556 1 557 644 645 cell_1rw
* cell instance $247 r0 *1 173.43,0
X$247 558 1 559 644 645 cell_1rw
* cell instance $248 r0 *1 174.135,0
X$248 560 1 561 644 645 cell_1rw
* cell instance $249 r0 *1 174.84,0
X$249 562 1 563 644 645 cell_1rw
* cell instance $250 r0 *1 175.545,0
X$250 564 1 565 644 645 cell_1rw
* cell instance $251 r0 *1 176.25,0
X$251 566 1 567 644 645 cell_1rw
* cell instance $252 r0 *1 176.955,0
X$252 568 1 569 644 645 cell_1rw
* cell instance $253 r0 *1 177.66,0
X$253 570 1 571 644 645 cell_1rw
* cell instance $254 r0 *1 178.365,0
X$254 572 1 573 644 645 cell_1rw
* cell instance $255 r0 *1 179.07,0
X$255 574 1 575 644 645 cell_1rw
* cell instance $256 r0 *1 179.775,0
X$256 576 1 577 644 645 cell_1rw
* cell instance $257 r0 *1 180.48,0
X$257 578 1 579 644 645 cell_1rw
* cell instance $258 m0 *1 0.705,2.73
X$258 67 2 68 644 645 cell_1rw
* cell instance $259 m0 *1 0,2.73
X$259 65 2 66 644 645 cell_1rw
* cell instance $260 m0 *1 1.41,2.73
X$260 69 2 70 644 645 cell_1rw
* cell instance $261 m0 *1 2.115,2.73
X$261 71 2 72 644 645 cell_1rw
* cell instance $262 m0 *1 2.82,2.73
X$262 73 2 74 644 645 cell_1rw
* cell instance $263 m0 *1 3.525,2.73
X$263 75 2 76 644 645 cell_1rw
* cell instance $264 m0 *1 4.23,2.73
X$264 77 2 78 644 645 cell_1rw
* cell instance $265 m0 *1 4.935,2.73
X$265 79 2 80 644 645 cell_1rw
* cell instance $266 m0 *1 5.64,2.73
X$266 81 2 82 644 645 cell_1rw
* cell instance $267 m0 *1 6.345,2.73
X$267 83 2 84 644 645 cell_1rw
* cell instance $268 m0 *1 7.05,2.73
X$268 85 2 86 644 645 cell_1rw
* cell instance $269 m0 *1 7.755,2.73
X$269 87 2 88 644 645 cell_1rw
* cell instance $270 m0 *1 8.46,2.73
X$270 89 2 90 644 645 cell_1rw
* cell instance $271 m0 *1 9.165,2.73
X$271 91 2 92 644 645 cell_1rw
* cell instance $272 m0 *1 9.87,2.73
X$272 93 2 94 644 645 cell_1rw
* cell instance $273 m0 *1 10.575,2.73
X$273 95 2 96 644 645 cell_1rw
* cell instance $274 m0 *1 11.28,2.73
X$274 97 2 98 644 645 cell_1rw
* cell instance $275 m0 *1 11.985,2.73
X$275 99 2 100 644 645 cell_1rw
* cell instance $276 m0 *1 12.69,2.73
X$276 101 2 102 644 645 cell_1rw
* cell instance $277 m0 *1 13.395,2.73
X$277 103 2 104 644 645 cell_1rw
* cell instance $278 m0 *1 14.1,2.73
X$278 105 2 106 644 645 cell_1rw
* cell instance $279 m0 *1 14.805,2.73
X$279 107 2 108 644 645 cell_1rw
* cell instance $280 m0 *1 15.51,2.73
X$280 109 2 110 644 645 cell_1rw
* cell instance $281 m0 *1 16.215,2.73
X$281 111 2 112 644 645 cell_1rw
* cell instance $282 m0 *1 16.92,2.73
X$282 113 2 114 644 645 cell_1rw
* cell instance $283 m0 *1 17.625,2.73
X$283 115 2 116 644 645 cell_1rw
* cell instance $284 m0 *1 18.33,2.73
X$284 117 2 118 644 645 cell_1rw
* cell instance $285 m0 *1 19.035,2.73
X$285 119 2 120 644 645 cell_1rw
* cell instance $286 m0 *1 19.74,2.73
X$286 121 2 122 644 645 cell_1rw
* cell instance $287 m0 *1 20.445,2.73
X$287 123 2 124 644 645 cell_1rw
* cell instance $288 m0 *1 21.15,2.73
X$288 125 2 126 644 645 cell_1rw
* cell instance $289 m0 *1 21.855,2.73
X$289 127 2 128 644 645 cell_1rw
* cell instance $290 m0 *1 22.56,2.73
X$290 129 2 130 644 645 cell_1rw
* cell instance $291 m0 *1 23.265,2.73
X$291 131 2 132 644 645 cell_1rw
* cell instance $292 m0 *1 23.97,2.73
X$292 133 2 134 644 645 cell_1rw
* cell instance $293 m0 *1 24.675,2.73
X$293 135 2 136 644 645 cell_1rw
* cell instance $294 m0 *1 25.38,2.73
X$294 137 2 138 644 645 cell_1rw
* cell instance $295 m0 *1 26.085,2.73
X$295 139 2 140 644 645 cell_1rw
* cell instance $296 m0 *1 26.79,2.73
X$296 141 2 142 644 645 cell_1rw
* cell instance $297 m0 *1 27.495,2.73
X$297 143 2 144 644 645 cell_1rw
* cell instance $298 m0 *1 28.2,2.73
X$298 145 2 146 644 645 cell_1rw
* cell instance $299 m0 *1 28.905,2.73
X$299 147 2 148 644 645 cell_1rw
* cell instance $300 m0 *1 29.61,2.73
X$300 149 2 150 644 645 cell_1rw
* cell instance $301 m0 *1 30.315,2.73
X$301 151 2 152 644 645 cell_1rw
* cell instance $302 m0 *1 31.02,2.73
X$302 153 2 154 644 645 cell_1rw
* cell instance $303 m0 *1 31.725,2.73
X$303 155 2 156 644 645 cell_1rw
* cell instance $304 m0 *1 32.43,2.73
X$304 157 2 158 644 645 cell_1rw
* cell instance $305 m0 *1 33.135,2.73
X$305 159 2 160 644 645 cell_1rw
* cell instance $306 m0 *1 33.84,2.73
X$306 161 2 162 644 645 cell_1rw
* cell instance $307 m0 *1 34.545,2.73
X$307 163 2 164 644 645 cell_1rw
* cell instance $308 m0 *1 35.25,2.73
X$308 165 2 166 644 645 cell_1rw
* cell instance $309 m0 *1 35.955,2.73
X$309 167 2 168 644 645 cell_1rw
* cell instance $310 m0 *1 36.66,2.73
X$310 169 2 170 644 645 cell_1rw
* cell instance $311 m0 *1 37.365,2.73
X$311 171 2 172 644 645 cell_1rw
* cell instance $312 m0 *1 38.07,2.73
X$312 173 2 174 644 645 cell_1rw
* cell instance $313 m0 *1 38.775,2.73
X$313 175 2 176 644 645 cell_1rw
* cell instance $314 m0 *1 39.48,2.73
X$314 177 2 178 644 645 cell_1rw
* cell instance $315 m0 *1 40.185,2.73
X$315 179 2 180 644 645 cell_1rw
* cell instance $316 m0 *1 40.89,2.73
X$316 181 2 182 644 645 cell_1rw
* cell instance $317 m0 *1 41.595,2.73
X$317 183 2 184 644 645 cell_1rw
* cell instance $318 m0 *1 42.3,2.73
X$318 185 2 186 644 645 cell_1rw
* cell instance $319 m0 *1 43.005,2.73
X$319 187 2 188 644 645 cell_1rw
* cell instance $320 m0 *1 43.71,2.73
X$320 189 2 190 644 645 cell_1rw
* cell instance $321 m0 *1 44.415,2.73
X$321 191 2 192 644 645 cell_1rw
* cell instance $322 m0 *1 45.12,2.73
X$322 193 2 194 644 645 cell_1rw
* cell instance $323 m0 *1 45.825,2.73
X$323 195 2 196 644 645 cell_1rw
* cell instance $324 m0 *1 46.53,2.73
X$324 197 2 198 644 645 cell_1rw
* cell instance $325 m0 *1 47.235,2.73
X$325 199 2 200 644 645 cell_1rw
* cell instance $326 m0 *1 47.94,2.73
X$326 201 2 202 644 645 cell_1rw
* cell instance $327 m0 *1 48.645,2.73
X$327 203 2 204 644 645 cell_1rw
* cell instance $328 m0 *1 49.35,2.73
X$328 205 2 206 644 645 cell_1rw
* cell instance $329 m0 *1 50.055,2.73
X$329 207 2 208 644 645 cell_1rw
* cell instance $330 m0 *1 50.76,2.73
X$330 209 2 210 644 645 cell_1rw
* cell instance $331 m0 *1 51.465,2.73
X$331 211 2 212 644 645 cell_1rw
* cell instance $332 m0 *1 52.17,2.73
X$332 213 2 214 644 645 cell_1rw
* cell instance $333 m0 *1 52.875,2.73
X$333 215 2 216 644 645 cell_1rw
* cell instance $334 m0 *1 53.58,2.73
X$334 217 2 218 644 645 cell_1rw
* cell instance $335 m0 *1 54.285,2.73
X$335 219 2 220 644 645 cell_1rw
* cell instance $336 m0 *1 54.99,2.73
X$336 221 2 222 644 645 cell_1rw
* cell instance $337 m0 *1 55.695,2.73
X$337 223 2 224 644 645 cell_1rw
* cell instance $338 m0 *1 56.4,2.73
X$338 225 2 226 644 645 cell_1rw
* cell instance $339 m0 *1 57.105,2.73
X$339 227 2 228 644 645 cell_1rw
* cell instance $340 m0 *1 57.81,2.73
X$340 229 2 230 644 645 cell_1rw
* cell instance $341 m0 *1 58.515,2.73
X$341 231 2 232 644 645 cell_1rw
* cell instance $342 m0 *1 59.22,2.73
X$342 233 2 234 644 645 cell_1rw
* cell instance $343 m0 *1 59.925,2.73
X$343 235 2 236 644 645 cell_1rw
* cell instance $344 m0 *1 60.63,2.73
X$344 237 2 238 644 645 cell_1rw
* cell instance $345 m0 *1 61.335,2.73
X$345 239 2 240 644 645 cell_1rw
* cell instance $346 m0 *1 62.04,2.73
X$346 241 2 242 644 645 cell_1rw
* cell instance $347 m0 *1 62.745,2.73
X$347 243 2 244 644 645 cell_1rw
* cell instance $348 m0 *1 63.45,2.73
X$348 245 2 246 644 645 cell_1rw
* cell instance $349 m0 *1 64.155,2.73
X$349 247 2 248 644 645 cell_1rw
* cell instance $350 m0 *1 64.86,2.73
X$350 249 2 250 644 645 cell_1rw
* cell instance $351 m0 *1 65.565,2.73
X$351 251 2 252 644 645 cell_1rw
* cell instance $352 m0 *1 66.27,2.73
X$352 253 2 254 644 645 cell_1rw
* cell instance $353 m0 *1 66.975,2.73
X$353 255 2 256 644 645 cell_1rw
* cell instance $354 m0 *1 67.68,2.73
X$354 257 2 258 644 645 cell_1rw
* cell instance $355 m0 *1 68.385,2.73
X$355 259 2 260 644 645 cell_1rw
* cell instance $356 m0 *1 69.09,2.73
X$356 261 2 262 644 645 cell_1rw
* cell instance $357 m0 *1 69.795,2.73
X$357 263 2 264 644 645 cell_1rw
* cell instance $358 m0 *1 70.5,2.73
X$358 265 2 266 644 645 cell_1rw
* cell instance $359 m0 *1 71.205,2.73
X$359 267 2 268 644 645 cell_1rw
* cell instance $360 m0 *1 71.91,2.73
X$360 269 2 270 644 645 cell_1rw
* cell instance $361 m0 *1 72.615,2.73
X$361 271 2 272 644 645 cell_1rw
* cell instance $362 m0 *1 73.32,2.73
X$362 273 2 274 644 645 cell_1rw
* cell instance $363 m0 *1 74.025,2.73
X$363 275 2 276 644 645 cell_1rw
* cell instance $364 m0 *1 74.73,2.73
X$364 277 2 278 644 645 cell_1rw
* cell instance $365 m0 *1 75.435,2.73
X$365 279 2 280 644 645 cell_1rw
* cell instance $366 m0 *1 76.14,2.73
X$366 281 2 282 644 645 cell_1rw
* cell instance $367 m0 *1 76.845,2.73
X$367 283 2 284 644 645 cell_1rw
* cell instance $368 m0 *1 77.55,2.73
X$368 285 2 286 644 645 cell_1rw
* cell instance $369 m0 *1 78.255,2.73
X$369 287 2 288 644 645 cell_1rw
* cell instance $370 m0 *1 78.96,2.73
X$370 289 2 290 644 645 cell_1rw
* cell instance $371 m0 *1 79.665,2.73
X$371 291 2 292 644 645 cell_1rw
* cell instance $372 m0 *1 80.37,2.73
X$372 293 2 294 644 645 cell_1rw
* cell instance $373 m0 *1 81.075,2.73
X$373 295 2 296 644 645 cell_1rw
* cell instance $374 m0 *1 81.78,2.73
X$374 297 2 298 644 645 cell_1rw
* cell instance $375 m0 *1 82.485,2.73
X$375 299 2 300 644 645 cell_1rw
* cell instance $376 m0 *1 83.19,2.73
X$376 301 2 302 644 645 cell_1rw
* cell instance $377 m0 *1 83.895,2.73
X$377 303 2 304 644 645 cell_1rw
* cell instance $378 m0 *1 84.6,2.73
X$378 305 2 306 644 645 cell_1rw
* cell instance $379 m0 *1 85.305,2.73
X$379 307 2 308 644 645 cell_1rw
* cell instance $380 m0 *1 86.01,2.73
X$380 309 2 310 644 645 cell_1rw
* cell instance $381 m0 *1 86.715,2.73
X$381 311 2 312 644 645 cell_1rw
* cell instance $382 m0 *1 87.42,2.73
X$382 313 2 314 644 645 cell_1rw
* cell instance $383 m0 *1 88.125,2.73
X$383 315 2 316 644 645 cell_1rw
* cell instance $384 m0 *1 88.83,2.73
X$384 317 2 318 644 645 cell_1rw
* cell instance $385 m0 *1 89.535,2.73
X$385 319 2 320 644 645 cell_1rw
* cell instance $386 m0 *1 90.24,2.73
X$386 321 2 323 644 645 cell_1rw
* cell instance $387 m0 *1 90.945,2.73
X$387 324 2 325 644 645 cell_1rw
* cell instance $388 m0 *1 91.65,2.73
X$388 326 2 327 644 645 cell_1rw
* cell instance $389 m0 *1 92.355,2.73
X$389 328 2 329 644 645 cell_1rw
* cell instance $390 m0 *1 93.06,2.73
X$390 330 2 331 644 645 cell_1rw
* cell instance $391 m0 *1 93.765,2.73
X$391 332 2 333 644 645 cell_1rw
* cell instance $392 m0 *1 94.47,2.73
X$392 334 2 335 644 645 cell_1rw
* cell instance $393 m0 *1 95.175,2.73
X$393 336 2 337 644 645 cell_1rw
* cell instance $394 m0 *1 95.88,2.73
X$394 338 2 339 644 645 cell_1rw
* cell instance $395 m0 *1 96.585,2.73
X$395 340 2 341 644 645 cell_1rw
* cell instance $396 m0 *1 97.29,2.73
X$396 342 2 343 644 645 cell_1rw
* cell instance $397 m0 *1 97.995,2.73
X$397 344 2 345 644 645 cell_1rw
* cell instance $398 m0 *1 98.7,2.73
X$398 346 2 347 644 645 cell_1rw
* cell instance $399 m0 *1 99.405,2.73
X$399 348 2 349 644 645 cell_1rw
* cell instance $400 m0 *1 100.11,2.73
X$400 350 2 351 644 645 cell_1rw
* cell instance $401 m0 *1 100.815,2.73
X$401 352 2 353 644 645 cell_1rw
* cell instance $402 m0 *1 101.52,2.73
X$402 354 2 355 644 645 cell_1rw
* cell instance $403 m0 *1 102.225,2.73
X$403 356 2 357 644 645 cell_1rw
* cell instance $404 m0 *1 102.93,2.73
X$404 358 2 359 644 645 cell_1rw
* cell instance $405 m0 *1 103.635,2.73
X$405 360 2 361 644 645 cell_1rw
* cell instance $406 m0 *1 104.34,2.73
X$406 362 2 363 644 645 cell_1rw
* cell instance $407 m0 *1 105.045,2.73
X$407 364 2 365 644 645 cell_1rw
* cell instance $408 m0 *1 105.75,2.73
X$408 366 2 367 644 645 cell_1rw
* cell instance $409 m0 *1 106.455,2.73
X$409 368 2 369 644 645 cell_1rw
* cell instance $410 m0 *1 107.16,2.73
X$410 370 2 371 644 645 cell_1rw
* cell instance $411 m0 *1 107.865,2.73
X$411 372 2 373 644 645 cell_1rw
* cell instance $412 m0 *1 108.57,2.73
X$412 374 2 375 644 645 cell_1rw
* cell instance $413 m0 *1 109.275,2.73
X$413 376 2 377 644 645 cell_1rw
* cell instance $414 m0 *1 109.98,2.73
X$414 378 2 379 644 645 cell_1rw
* cell instance $415 m0 *1 110.685,2.73
X$415 380 2 381 644 645 cell_1rw
* cell instance $416 m0 *1 111.39,2.73
X$416 382 2 383 644 645 cell_1rw
* cell instance $417 m0 *1 112.095,2.73
X$417 384 2 385 644 645 cell_1rw
* cell instance $418 m0 *1 112.8,2.73
X$418 386 2 387 644 645 cell_1rw
* cell instance $419 m0 *1 113.505,2.73
X$419 388 2 389 644 645 cell_1rw
* cell instance $420 m0 *1 114.21,2.73
X$420 390 2 391 644 645 cell_1rw
* cell instance $421 m0 *1 114.915,2.73
X$421 392 2 393 644 645 cell_1rw
* cell instance $422 m0 *1 115.62,2.73
X$422 394 2 395 644 645 cell_1rw
* cell instance $423 m0 *1 116.325,2.73
X$423 396 2 397 644 645 cell_1rw
* cell instance $424 m0 *1 117.03,2.73
X$424 398 2 399 644 645 cell_1rw
* cell instance $425 m0 *1 117.735,2.73
X$425 400 2 401 644 645 cell_1rw
* cell instance $426 m0 *1 118.44,2.73
X$426 402 2 403 644 645 cell_1rw
* cell instance $427 m0 *1 119.145,2.73
X$427 404 2 405 644 645 cell_1rw
* cell instance $428 m0 *1 119.85,2.73
X$428 406 2 407 644 645 cell_1rw
* cell instance $429 m0 *1 120.555,2.73
X$429 408 2 409 644 645 cell_1rw
* cell instance $430 m0 *1 121.26,2.73
X$430 410 2 411 644 645 cell_1rw
* cell instance $431 m0 *1 121.965,2.73
X$431 412 2 413 644 645 cell_1rw
* cell instance $432 m0 *1 122.67,2.73
X$432 414 2 415 644 645 cell_1rw
* cell instance $433 m0 *1 123.375,2.73
X$433 416 2 417 644 645 cell_1rw
* cell instance $434 m0 *1 124.08,2.73
X$434 418 2 419 644 645 cell_1rw
* cell instance $435 m0 *1 124.785,2.73
X$435 420 2 421 644 645 cell_1rw
* cell instance $436 m0 *1 125.49,2.73
X$436 422 2 423 644 645 cell_1rw
* cell instance $437 m0 *1 126.195,2.73
X$437 424 2 425 644 645 cell_1rw
* cell instance $438 m0 *1 126.9,2.73
X$438 426 2 427 644 645 cell_1rw
* cell instance $439 m0 *1 127.605,2.73
X$439 428 2 429 644 645 cell_1rw
* cell instance $440 m0 *1 128.31,2.73
X$440 430 2 431 644 645 cell_1rw
* cell instance $441 m0 *1 129.015,2.73
X$441 432 2 433 644 645 cell_1rw
* cell instance $442 m0 *1 129.72,2.73
X$442 434 2 435 644 645 cell_1rw
* cell instance $443 m0 *1 130.425,2.73
X$443 436 2 437 644 645 cell_1rw
* cell instance $444 m0 *1 131.13,2.73
X$444 438 2 439 644 645 cell_1rw
* cell instance $445 m0 *1 131.835,2.73
X$445 440 2 441 644 645 cell_1rw
* cell instance $446 m0 *1 132.54,2.73
X$446 442 2 443 644 645 cell_1rw
* cell instance $447 m0 *1 133.245,2.73
X$447 444 2 445 644 645 cell_1rw
* cell instance $448 m0 *1 133.95,2.73
X$448 446 2 447 644 645 cell_1rw
* cell instance $449 m0 *1 134.655,2.73
X$449 448 2 449 644 645 cell_1rw
* cell instance $450 m0 *1 135.36,2.73
X$450 450 2 451 644 645 cell_1rw
* cell instance $451 m0 *1 136.065,2.73
X$451 452 2 453 644 645 cell_1rw
* cell instance $452 m0 *1 136.77,2.73
X$452 454 2 455 644 645 cell_1rw
* cell instance $453 m0 *1 137.475,2.73
X$453 456 2 457 644 645 cell_1rw
* cell instance $454 m0 *1 138.18,2.73
X$454 458 2 459 644 645 cell_1rw
* cell instance $455 m0 *1 138.885,2.73
X$455 460 2 461 644 645 cell_1rw
* cell instance $456 m0 *1 139.59,2.73
X$456 462 2 463 644 645 cell_1rw
* cell instance $457 m0 *1 140.295,2.73
X$457 464 2 465 644 645 cell_1rw
* cell instance $458 m0 *1 141,2.73
X$458 466 2 467 644 645 cell_1rw
* cell instance $459 m0 *1 141.705,2.73
X$459 468 2 469 644 645 cell_1rw
* cell instance $460 m0 *1 142.41,2.73
X$460 470 2 471 644 645 cell_1rw
* cell instance $461 m0 *1 143.115,2.73
X$461 472 2 473 644 645 cell_1rw
* cell instance $462 m0 *1 143.82,2.73
X$462 474 2 475 644 645 cell_1rw
* cell instance $463 m0 *1 144.525,2.73
X$463 476 2 477 644 645 cell_1rw
* cell instance $464 m0 *1 145.23,2.73
X$464 478 2 479 644 645 cell_1rw
* cell instance $465 m0 *1 145.935,2.73
X$465 480 2 481 644 645 cell_1rw
* cell instance $466 m0 *1 146.64,2.73
X$466 482 2 483 644 645 cell_1rw
* cell instance $467 m0 *1 147.345,2.73
X$467 484 2 485 644 645 cell_1rw
* cell instance $468 m0 *1 148.05,2.73
X$468 486 2 487 644 645 cell_1rw
* cell instance $469 m0 *1 148.755,2.73
X$469 488 2 489 644 645 cell_1rw
* cell instance $470 m0 *1 149.46,2.73
X$470 490 2 491 644 645 cell_1rw
* cell instance $471 m0 *1 150.165,2.73
X$471 492 2 493 644 645 cell_1rw
* cell instance $472 m0 *1 150.87,2.73
X$472 494 2 495 644 645 cell_1rw
* cell instance $473 m0 *1 151.575,2.73
X$473 496 2 497 644 645 cell_1rw
* cell instance $474 m0 *1 152.28,2.73
X$474 498 2 499 644 645 cell_1rw
* cell instance $475 m0 *1 152.985,2.73
X$475 500 2 501 644 645 cell_1rw
* cell instance $476 m0 *1 153.69,2.73
X$476 502 2 503 644 645 cell_1rw
* cell instance $477 m0 *1 154.395,2.73
X$477 504 2 505 644 645 cell_1rw
* cell instance $478 m0 *1 155.1,2.73
X$478 506 2 507 644 645 cell_1rw
* cell instance $479 m0 *1 155.805,2.73
X$479 508 2 509 644 645 cell_1rw
* cell instance $480 m0 *1 156.51,2.73
X$480 510 2 511 644 645 cell_1rw
* cell instance $481 m0 *1 157.215,2.73
X$481 512 2 513 644 645 cell_1rw
* cell instance $482 m0 *1 157.92,2.73
X$482 514 2 515 644 645 cell_1rw
* cell instance $483 m0 *1 158.625,2.73
X$483 516 2 517 644 645 cell_1rw
* cell instance $484 m0 *1 159.33,2.73
X$484 518 2 519 644 645 cell_1rw
* cell instance $485 m0 *1 160.035,2.73
X$485 520 2 521 644 645 cell_1rw
* cell instance $486 m0 *1 160.74,2.73
X$486 522 2 523 644 645 cell_1rw
* cell instance $487 m0 *1 161.445,2.73
X$487 524 2 525 644 645 cell_1rw
* cell instance $488 m0 *1 162.15,2.73
X$488 526 2 527 644 645 cell_1rw
* cell instance $489 m0 *1 162.855,2.73
X$489 528 2 529 644 645 cell_1rw
* cell instance $490 m0 *1 163.56,2.73
X$490 530 2 531 644 645 cell_1rw
* cell instance $491 m0 *1 164.265,2.73
X$491 532 2 533 644 645 cell_1rw
* cell instance $492 m0 *1 164.97,2.73
X$492 534 2 535 644 645 cell_1rw
* cell instance $493 m0 *1 165.675,2.73
X$493 536 2 537 644 645 cell_1rw
* cell instance $494 m0 *1 166.38,2.73
X$494 538 2 539 644 645 cell_1rw
* cell instance $495 m0 *1 167.085,2.73
X$495 540 2 541 644 645 cell_1rw
* cell instance $496 m0 *1 167.79,2.73
X$496 542 2 543 644 645 cell_1rw
* cell instance $497 m0 *1 168.495,2.73
X$497 544 2 545 644 645 cell_1rw
* cell instance $498 m0 *1 169.2,2.73
X$498 546 2 547 644 645 cell_1rw
* cell instance $499 m0 *1 169.905,2.73
X$499 548 2 549 644 645 cell_1rw
* cell instance $500 m0 *1 170.61,2.73
X$500 550 2 551 644 645 cell_1rw
* cell instance $501 m0 *1 171.315,2.73
X$501 552 2 553 644 645 cell_1rw
* cell instance $502 m0 *1 172.02,2.73
X$502 554 2 555 644 645 cell_1rw
* cell instance $503 m0 *1 172.725,2.73
X$503 556 2 557 644 645 cell_1rw
* cell instance $504 m0 *1 173.43,2.73
X$504 558 2 559 644 645 cell_1rw
* cell instance $505 m0 *1 174.135,2.73
X$505 560 2 561 644 645 cell_1rw
* cell instance $506 m0 *1 174.84,2.73
X$506 562 2 563 644 645 cell_1rw
* cell instance $507 m0 *1 175.545,2.73
X$507 564 2 565 644 645 cell_1rw
* cell instance $508 m0 *1 176.25,2.73
X$508 566 2 567 644 645 cell_1rw
* cell instance $509 m0 *1 176.955,2.73
X$509 568 2 569 644 645 cell_1rw
* cell instance $510 m0 *1 177.66,2.73
X$510 570 2 571 644 645 cell_1rw
* cell instance $511 m0 *1 178.365,2.73
X$511 572 2 573 644 645 cell_1rw
* cell instance $512 m0 *1 179.07,2.73
X$512 574 2 575 644 645 cell_1rw
* cell instance $513 m0 *1 179.775,2.73
X$513 576 2 577 644 645 cell_1rw
* cell instance $514 m0 *1 180.48,2.73
X$514 578 2 579 644 645 cell_1rw
* cell instance $515 m0 *1 0.705,5.46
X$515 67 3 68 644 645 cell_1rw
* cell instance $516 m0 *1 0,5.46
X$516 65 3 66 644 645 cell_1rw
* cell instance $517 m0 *1 1.41,5.46
X$517 69 3 70 644 645 cell_1rw
* cell instance $518 m0 *1 2.115,5.46
X$518 71 3 72 644 645 cell_1rw
* cell instance $519 m0 *1 2.82,5.46
X$519 73 3 74 644 645 cell_1rw
* cell instance $520 m0 *1 3.525,5.46
X$520 75 3 76 644 645 cell_1rw
* cell instance $521 m0 *1 4.23,5.46
X$521 77 3 78 644 645 cell_1rw
* cell instance $522 m0 *1 4.935,5.46
X$522 79 3 80 644 645 cell_1rw
* cell instance $523 m0 *1 5.64,5.46
X$523 81 3 82 644 645 cell_1rw
* cell instance $524 m0 *1 6.345,5.46
X$524 83 3 84 644 645 cell_1rw
* cell instance $525 m0 *1 7.05,5.46
X$525 85 3 86 644 645 cell_1rw
* cell instance $526 m0 *1 7.755,5.46
X$526 87 3 88 644 645 cell_1rw
* cell instance $527 m0 *1 8.46,5.46
X$527 89 3 90 644 645 cell_1rw
* cell instance $528 m0 *1 9.165,5.46
X$528 91 3 92 644 645 cell_1rw
* cell instance $529 m0 *1 9.87,5.46
X$529 93 3 94 644 645 cell_1rw
* cell instance $530 m0 *1 10.575,5.46
X$530 95 3 96 644 645 cell_1rw
* cell instance $531 m0 *1 11.28,5.46
X$531 97 3 98 644 645 cell_1rw
* cell instance $532 m0 *1 11.985,5.46
X$532 99 3 100 644 645 cell_1rw
* cell instance $533 m0 *1 12.69,5.46
X$533 101 3 102 644 645 cell_1rw
* cell instance $534 m0 *1 13.395,5.46
X$534 103 3 104 644 645 cell_1rw
* cell instance $535 m0 *1 14.1,5.46
X$535 105 3 106 644 645 cell_1rw
* cell instance $536 m0 *1 14.805,5.46
X$536 107 3 108 644 645 cell_1rw
* cell instance $537 m0 *1 15.51,5.46
X$537 109 3 110 644 645 cell_1rw
* cell instance $538 m0 *1 16.215,5.46
X$538 111 3 112 644 645 cell_1rw
* cell instance $539 m0 *1 16.92,5.46
X$539 113 3 114 644 645 cell_1rw
* cell instance $540 m0 *1 17.625,5.46
X$540 115 3 116 644 645 cell_1rw
* cell instance $541 m0 *1 18.33,5.46
X$541 117 3 118 644 645 cell_1rw
* cell instance $542 m0 *1 19.035,5.46
X$542 119 3 120 644 645 cell_1rw
* cell instance $543 m0 *1 19.74,5.46
X$543 121 3 122 644 645 cell_1rw
* cell instance $544 m0 *1 20.445,5.46
X$544 123 3 124 644 645 cell_1rw
* cell instance $545 m0 *1 21.15,5.46
X$545 125 3 126 644 645 cell_1rw
* cell instance $546 m0 *1 21.855,5.46
X$546 127 3 128 644 645 cell_1rw
* cell instance $547 m0 *1 22.56,5.46
X$547 129 3 130 644 645 cell_1rw
* cell instance $548 m0 *1 23.265,5.46
X$548 131 3 132 644 645 cell_1rw
* cell instance $549 m0 *1 23.97,5.46
X$549 133 3 134 644 645 cell_1rw
* cell instance $550 m0 *1 24.675,5.46
X$550 135 3 136 644 645 cell_1rw
* cell instance $551 m0 *1 25.38,5.46
X$551 137 3 138 644 645 cell_1rw
* cell instance $552 m0 *1 26.085,5.46
X$552 139 3 140 644 645 cell_1rw
* cell instance $553 m0 *1 26.79,5.46
X$553 141 3 142 644 645 cell_1rw
* cell instance $554 m0 *1 27.495,5.46
X$554 143 3 144 644 645 cell_1rw
* cell instance $555 m0 *1 28.2,5.46
X$555 145 3 146 644 645 cell_1rw
* cell instance $556 m0 *1 28.905,5.46
X$556 147 3 148 644 645 cell_1rw
* cell instance $557 m0 *1 29.61,5.46
X$557 149 3 150 644 645 cell_1rw
* cell instance $558 m0 *1 30.315,5.46
X$558 151 3 152 644 645 cell_1rw
* cell instance $559 m0 *1 31.02,5.46
X$559 153 3 154 644 645 cell_1rw
* cell instance $560 m0 *1 31.725,5.46
X$560 155 3 156 644 645 cell_1rw
* cell instance $561 m0 *1 32.43,5.46
X$561 157 3 158 644 645 cell_1rw
* cell instance $562 m0 *1 33.135,5.46
X$562 159 3 160 644 645 cell_1rw
* cell instance $563 m0 *1 33.84,5.46
X$563 161 3 162 644 645 cell_1rw
* cell instance $564 m0 *1 34.545,5.46
X$564 163 3 164 644 645 cell_1rw
* cell instance $565 m0 *1 35.25,5.46
X$565 165 3 166 644 645 cell_1rw
* cell instance $566 m0 *1 35.955,5.46
X$566 167 3 168 644 645 cell_1rw
* cell instance $567 m0 *1 36.66,5.46
X$567 169 3 170 644 645 cell_1rw
* cell instance $568 m0 *1 37.365,5.46
X$568 171 3 172 644 645 cell_1rw
* cell instance $569 m0 *1 38.07,5.46
X$569 173 3 174 644 645 cell_1rw
* cell instance $570 m0 *1 38.775,5.46
X$570 175 3 176 644 645 cell_1rw
* cell instance $571 m0 *1 39.48,5.46
X$571 177 3 178 644 645 cell_1rw
* cell instance $572 m0 *1 40.185,5.46
X$572 179 3 180 644 645 cell_1rw
* cell instance $573 m0 *1 40.89,5.46
X$573 181 3 182 644 645 cell_1rw
* cell instance $574 m0 *1 41.595,5.46
X$574 183 3 184 644 645 cell_1rw
* cell instance $575 m0 *1 42.3,5.46
X$575 185 3 186 644 645 cell_1rw
* cell instance $576 m0 *1 43.005,5.46
X$576 187 3 188 644 645 cell_1rw
* cell instance $577 m0 *1 43.71,5.46
X$577 189 3 190 644 645 cell_1rw
* cell instance $578 m0 *1 44.415,5.46
X$578 191 3 192 644 645 cell_1rw
* cell instance $579 m0 *1 45.12,5.46
X$579 193 3 194 644 645 cell_1rw
* cell instance $580 m0 *1 45.825,5.46
X$580 195 3 196 644 645 cell_1rw
* cell instance $581 m0 *1 46.53,5.46
X$581 197 3 198 644 645 cell_1rw
* cell instance $582 m0 *1 47.235,5.46
X$582 199 3 200 644 645 cell_1rw
* cell instance $583 m0 *1 47.94,5.46
X$583 201 3 202 644 645 cell_1rw
* cell instance $584 m0 *1 48.645,5.46
X$584 203 3 204 644 645 cell_1rw
* cell instance $585 m0 *1 49.35,5.46
X$585 205 3 206 644 645 cell_1rw
* cell instance $586 m0 *1 50.055,5.46
X$586 207 3 208 644 645 cell_1rw
* cell instance $587 m0 *1 50.76,5.46
X$587 209 3 210 644 645 cell_1rw
* cell instance $588 m0 *1 51.465,5.46
X$588 211 3 212 644 645 cell_1rw
* cell instance $589 m0 *1 52.17,5.46
X$589 213 3 214 644 645 cell_1rw
* cell instance $590 m0 *1 52.875,5.46
X$590 215 3 216 644 645 cell_1rw
* cell instance $591 m0 *1 53.58,5.46
X$591 217 3 218 644 645 cell_1rw
* cell instance $592 m0 *1 54.285,5.46
X$592 219 3 220 644 645 cell_1rw
* cell instance $593 m0 *1 54.99,5.46
X$593 221 3 222 644 645 cell_1rw
* cell instance $594 m0 *1 55.695,5.46
X$594 223 3 224 644 645 cell_1rw
* cell instance $595 m0 *1 56.4,5.46
X$595 225 3 226 644 645 cell_1rw
* cell instance $596 m0 *1 57.105,5.46
X$596 227 3 228 644 645 cell_1rw
* cell instance $597 m0 *1 57.81,5.46
X$597 229 3 230 644 645 cell_1rw
* cell instance $598 m0 *1 58.515,5.46
X$598 231 3 232 644 645 cell_1rw
* cell instance $599 m0 *1 59.22,5.46
X$599 233 3 234 644 645 cell_1rw
* cell instance $600 m0 *1 59.925,5.46
X$600 235 3 236 644 645 cell_1rw
* cell instance $601 m0 *1 60.63,5.46
X$601 237 3 238 644 645 cell_1rw
* cell instance $602 m0 *1 61.335,5.46
X$602 239 3 240 644 645 cell_1rw
* cell instance $603 m0 *1 62.04,5.46
X$603 241 3 242 644 645 cell_1rw
* cell instance $604 m0 *1 62.745,5.46
X$604 243 3 244 644 645 cell_1rw
* cell instance $605 m0 *1 63.45,5.46
X$605 245 3 246 644 645 cell_1rw
* cell instance $606 m0 *1 64.155,5.46
X$606 247 3 248 644 645 cell_1rw
* cell instance $607 m0 *1 64.86,5.46
X$607 249 3 250 644 645 cell_1rw
* cell instance $608 m0 *1 65.565,5.46
X$608 251 3 252 644 645 cell_1rw
* cell instance $609 m0 *1 66.27,5.46
X$609 253 3 254 644 645 cell_1rw
* cell instance $610 m0 *1 66.975,5.46
X$610 255 3 256 644 645 cell_1rw
* cell instance $611 m0 *1 67.68,5.46
X$611 257 3 258 644 645 cell_1rw
* cell instance $612 m0 *1 68.385,5.46
X$612 259 3 260 644 645 cell_1rw
* cell instance $613 m0 *1 69.09,5.46
X$613 261 3 262 644 645 cell_1rw
* cell instance $614 m0 *1 69.795,5.46
X$614 263 3 264 644 645 cell_1rw
* cell instance $615 m0 *1 70.5,5.46
X$615 265 3 266 644 645 cell_1rw
* cell instance $616 m0 *1 71.205,5.46
X$616 267 3 268 644 645 cell_1rw
* cell instance $617 m0 *1 71.91,5.46
X$617 269 3 270 644 645 cell_1rw
* cell instance $618 m0 *1 72.615,5.46
X$618 271 3 272 644 645 cell_1rw
* cell instance $619 m0 *1 73.32,5.46
X$619 273 3 274 644 645 cell_1rw
* cell instance $620 m0 *1 74.025,5.46
X$620 275 3 276 644 645 cell_1rw
* cell instance $621 m0 *1 74.73,5.46
X$621 277 3 278 644 645 cell_1rw
* cell instance $622 m0 *1 75.435,5.46
X$622 279 3 280 644 645 cell_1rw
* cell instance $623 m0 *1 76.14,5.46
X$623 281 3 282 644 645 cell_1rw
* cell instance $624 m0 *1 76.845,5.46
X$624 283 3 284 644 645 cell_1rw
* cell instance $625 m0 *1 77.55,5.46
X$625 285 3 286 644 645 cell_1rw
* cell instance $626 m0 *1 78.255,5.46
X$626 287 3 288 644 645 cell_1rw
* cell instance $627 m0 *1 78.96,5.46
X$627 289 3 290 644 645 cell_1rw
* cell instance $628 m0 *1 79.665,5.46
X$628 291 3 292 644 645 cell_1rw
* cell instance $629 m0 *1 80.37,5.46
X$629 293 3 294 644 645 cell_1rw
* cell instance $630 m0 *1 81.075,5.46
X$630 295 3 296 644 645 cell_1rw
* cell instance $631 m0 *1 81.78,5.46
X$631 297 3 298 644 645 cell_1rw
* cell instance $632 m0 *1 82.485,5.46
X$632 299 3 300 644 645 cell_1rw
* cell instance $633 m0 *1 83.19,5.46
X$633 301 3 302 644 645 cell_1rw
* cell instance $634 m0 *1 83.895,5.46
X$634 303 3 304 644 645 cell_1rw
* cell instance $635 m0 *1 84.6,5.46
X$635 305 3 306 644 645 cell_1rw
* cell instance $636 m0 *1 85.305,5.46
X$636 307 3 308 644 645 cell_1rw
* cell instance $637 m0 *1 86.01,5.46
X$637 309 3 310 644 645 cell_1rw
* cell instance $638 m0 *1 86.715,5.46
X$638 311 3 312 644 645 cell_1rw
* cell instance $639 m0 *1 87.42,5.46
X$639 313 3 314 644 645 cell_1rw
* cell instance $640 m0 *1 88.125,5.46
X$640 315 3 316 644 645 cell_1rw
* cell instance $641 m0 *1 88.83,5.46
X$641 317 3 318 644 645 cell_1rw
* cell instance $642 m0 *1 89.535,5.46
X$642 319 3 320 644 645 cell_1rw
* cell instance $643 m0 *1 90.24,5.46
X$643 321 3 323 644 645 cell_1rw
* cell instance $644 m0 *1 90.945,5.46
X$644 324 3 325 644 645 cell_1rw
* cell instance $645 m0 *1 91.65,5.46
X$645 326 3 327 644 645 cell_1rw
* cell instance $646 m0 *1 92.355,5.46
X$646 328 3 329 644 645 cell_1rw
* cell instance $647 m0 *1 93.06,5.46
X$647 330 3 331 644 645 cell_1rw
* cell instance $648 m0 *1 93.765,5.46
X$648 332 3 333 644 645 cell_1rw
* cell instance $649 m0 *1 94.47,5.46
X$649 334 3 335 644 645 cell_1rw
* cell instance $650 m0 *1 95.175,5.46
X$650 336 3 337 644 645 cell_1rw
* cell instance $651 m0 *1 95.88,5.46
X$651 338 3 339 644 645 cell_1rw
* cell instance $652 m0 *1 96.585,5.46
X$652 340 3 341 644 645 cell_1rw
* cell instance $653 m0 *1 97.29,5.46
X$653 342 3 343 644 645 cell_1rw
* cell instance $654 m0 *1 97.995,5.46
X$654 344 3 345 644 645 cell_1rw
* cell instance $655 m0 *1 98.7,5.46
X$655 346 3 347 644 645 cell_1rw
* cell instance $656 m0 *1 99.405,5.46
X$656 348 3 349 644 645 cell_1rw
* cell instance $657 m0 *1 100.11,5.46
X$657 350 3 351 644 645 cell_1rw
* cell instance $658 m0 *1 100.815,5.46
X$658 352 3 353 644 645 cell_1rw
* cell instance $659 m0 *1 101.52,5.46
X$659 354 3 355 644 645 cell_1rw
* cell instance $660 m0 *1 102.225,5.46
X$660 356 3 357 644 645 cell_1rw
* cell instance $661 m0 *1 102.93,5.46
X$661 358 3 359 644 645 cell_1rw
* cell instance $662 m0 *1 103.635,5.46
X$662 360 3 361 644 645 cell_1rw
* cell instance $663 m0 *1 104.34,5.46
X$663 362 3 363 644 645 cell_1rw
* cell instance $664 m0 *1 105.045,5.46
X$664 364 3 365 644 645 cell_1rw
* cell instance $665 m0 *1 105.75,5.46
X$665 366 3 367 644 645 cell_1rw
* cell instance $666 m0 *1 106.455,5.46
X$666 368 3 369 644 645 cell_1rw
* cell instance $667 m0 *1 107.16,5.46
X$667 370 3 371 644 645 cell_1rw
* cell instance $668 m0 *1 107.865,5.46
X$668 372 3 373 644 645 cell_1rw
* cell instance $669 m0 *1 108.57,5.46
X$669 374 3 375 644 645 cell_1rw
* cell instance $670 m0 *1 109.275,5.46
X$670 376 3 377 644 645 cell_1rw
* cell instance $671 m0 *1 109.98,5.46
X$671 378 3 379 644 645 cell_1rw
* cell instance $672 m0 *1 110.685,5.46
X$672 380 3 381 644 645 cell_1rw
* cell instance $673 m0 *1 111.39,5.46
X$673 382 3 383 644 645 cell_1rw
* cell instance $674 m0 *1 112.095,5.46
X$674 384 3 385 644 645 cell_1rw
* cell instance $675 m0 *1 112.8,5.46
X$675 386 3 387 644 645 cell_1rw
* cell instance $676 m0 *1 113.505,5.46
X$676 388 3 389 644 645 cell_1rw
* cell instance $677 m0 *1 114.21,5.46
X$677 390 3 391 644 645 cell_1rw
* cell instance $678 m0 *1 114.915,5.46
X$678 392 3 393 644 645 cell_1rw
* cell instance $679 m0 *1 115.62,5.46
X$679 394 3 395 644 645 cell_1rw
* cell instance $680 m0 *1 116.325,5.46
X$680 396 3 397 644 645 cell_1rw
* cell instance $681 m0 *1 117.03,5.46
X$681 398 3 399 644 645 cell_1rw
* cell instance $682 m0 *1 117.735,5.46
X$682 400 3 401 644 645 cell_1rw
* cell instance $683 m0 *1 118.44,5.46
X$683 402 3 403 644 645 cell_1rw
* cell instance $684 m0 *1 119.145,5.46
X$684 404 3 405 644 645 cell_1rw
* cell instance $685 m0 *1 119.85,5.46
X$685 406 3 407 644 645 cell_1rw
* cell instance $686 m0 *1 120.555,5.46
X$686 408 3 409 644 645 cell_1rw
* cell instance $687 m0 *1 121.26,5.46
X$687 410 3 411 644 645 cell_1rw
* cell instance $688 m0 *1 121.965,5.46
X$688 412 3 413 644 645 cell_1rw
* cell instance $689 m0 *1 122.67,5.46
X$689 414 3 415 644 645 cell_1rw
* cell instance $690 m0 *1 123.375,5.46
X$690 416 3 417 644 645 cell_1rw
* cell instance $691 m0 *1 124.08,5.46
X$691 418 3 419 644 645 cell_1rw
* cell instance $692 m0 *1 124.785,5.46
X$692 420 3 421 644 645 cell_1rw
* cell instance $693 m0 *1 125.49,5.46
X$693 422 3 423 644 645 cell_1rw
* cell instance $694 m0 *1 126.195,5.46
X$694 424 3 425 644 645 cell_1rw
* cell instance $695 m0 *1 126.9,5.46
X$695 426 3 427 644 645 cell_1rw
* cell instance $696 m0 *1 127.605,5.46
X$696 428 3 429 644 645 cell_1rw
* cell instance $697 m0 *1 128.31,5.46
X$697 430 3 431 644 645 cell_1rw
* cell instance $698 m0 *1 129.015,5.46
X$698 432 3 433 644 645 cell_1rw
* cell instance $699 m0 *1 129.72,5.46
X$699 434 3 435 644 645 cell_1rw
* cell instance $700 m0 *1 130.425,5.46
X$700 436 3 437 644 645 cell_1rw
* cell instance $701 m0 *1 131.13,5.46
X$701 438 3 439 644 645 cell_1rw
* cell instance $702 m0 *1 131.835,5.46
X$702 440 3 441 644 645 cell_1rw
* cell instance $703 m0 *1 132.54,5.46
X$703 442 3 443 644 645 cell_1rw
* cell instance $704 m0 *1 133.245,5.46
X$704 444 3 445 644 645 cell_1rw
* cell instance $705 m0 *1 133.95,5.46
X$705 446 3 447 644 645 cell_1rw
* cell instance $706 m0 *1 134.655,5.46
X$706 448 3 449 644 645 cell_1rw
* cell instance $707 m0 *1 135.36,5.46
X$707 450 3 451 644 645 cell_1rw
* cell instance $708 m0 *1 136.065,5.46
X$708 452 3 453 644 645 cell_1rw
* cell instance $709 m0 *1 136.77,5.46
X$709 454 3 455 644 645 cell_1rw
* cell instance $710 m0 *1 137.475,5.46
X$710 456 3 457 644 645 cell_1rw
* cell instance $711 m0 *1 138.18,5.46
X$711 458 3 459 644 645 cell_1rw
* cell instance $712 m0 *1 138.885,5.46
X$712 460 3 461 644 645 cell_1rw
* cell instance $713 m0 *1 139.59,5.46
X$713 462 3 463 644 645 cell_1rw
* cell instance $714 m0 *1 140.295,5.46
X$714 464 3 465 644 645 cell_1rw
* cell instance $715 m0 *1 141,5.46
X$715 466 3 467 644 645 cell_1rw
* cell instance $716 m0 *1 141.705,5.46
X$716 468 3 469 644 645 cell_1rw
* cell instance $717 m0 *1 142.41,5.46
X$717 470 3 471 644 645 cell_1rw
* cell instance $718 m0 *1 143.115,5.46
X$718 472 3 473 644 645 cell_1rw
* cell instance $719 m0 *1 143.82,5.46
X$719 474 3 475 644 645 cell_1rw
* cell instance $720 m0 *1 144.525,5.46
X$720 476 3 477 644 645 cell_1rw
* cell instance $721 m0 *1 145.23,5.46
X$721 478 3 479 644 645 cell_1rw
* cell instance $722 m0 *1 145.935,5.46
X$722 480 3 481 644 645 cell_1rw
* cell instance $723 m0 *1 146.64,5.46
X$723 482 3 483 644 645 cell_1rw
* cell instance $724 m0 *1 147.345,5.46
X$724 484 3 485 644 645 cell_1rw
* cell instance $725 m0 *1 148.05,5.46
X$725 486 3 487 644 645 cell_1rw
* cell instance $726 m0 *1 148.755,5.46
X$726 488 3 489 644 645 cell_1rw
* cell instance $727 m0 *1 149.46,5.46
X$727 490 3 491 644 645 cell_1rw
* cell instance $728 m0 *1 150.165,5.46
X$728 492 3 493 644 645 cell_1rw
* cell instance $729 m0 *1 150.87,5.46
X$729 494 3 495 644 645 cell_1rw
* cell instance $730 m0 *1 151.575,5.46
X$730 496 3 497 644 645 cell_1rw
* cell instance $731 m0 *1 152.28,5.46
X$731 498 3 499 644 645 cell_1rw
* cell instance $732 m0 *1 152.985,5.46
X$732 500 3 501 644 645 cell_1rw
* cell instance $733 m0 *1 153.69,5.46
X$733 502 3 503 644 645 cell_1rw
* cell instance $734 m0 *1 154.395,5.46
X$734 504 3 505 644 645 cell_1rw
* cell instance $735 m0 *1 155.1,5.46
X$735 506 3 507 644 645 cell_1rw
* cell instance $736 m0 *1 155.805,5.46
X$736 508 3 509 644 645 cell_1rw
* cell instance $737 m0 *1 156.51,5.46
X$737 510 3 511 644 645 cell_1rw
* cell instance $738 m0 *1 157.215,5.46
X$738 512 3 513 644 645 cell_1rw
* cell instance $739 m0 *1 157.92,5.46
X$739 514 3 515 644 645 cell_1rw
* cell instance $740 m0 *1 158.625,5.46
X$740 516 3 517 644 645 cell_1rw
* cell instance $741 m0 *1 159.33,5.46
X$741 518 3 519 644 645 cell_1rw
* cell instance $742 m0 *1 160.035,5.46
X$742 520 3 521 644 645 cell_1rw
* cell instance $743 m0 *1 160.74,5.46
X$743 522 3 523 644 645 cell_1rw
* cell instance $744 m0 *1 161.445,5.46
X$744 524 3 525 644 645 cell_1rw
* cell instance $745 m0 *1 162.15,5.46
X$745 526 3 527 644 645 cell_1rw
* cell instance $746 m0 *1 162.855,5.46
X$746 528 3 529 644 645 cell_1rw
* cell instance $747 m0 *1 163.56,5.46
X$747 530 3 531 644 645 cell_1rw
* cell instance $748 m0 *1 164.265,5.46
X$748 532 3 533 644 645 cell_1rw
* cell instance $749 m0 *1 164.97,5.46
X$749 534 3 535 644 645 cell_1rw
* cell instance $750 m0 *1 165.675,5.46
X$750 536 3 537 644 645 cell_1rw
* cell instance $751 m0 *1 166.38,5.46
X$751 538 3 539 644 645 cell_1rw
* cell instance $752 m0 *1 167.085,5.46
X$752 540 3 541 644 645 cell_1rw
* cell instance $753 m0 *1 167.79,5.46
X$753 542 3 543 644 645 cell_1rw
* cell instance $754 m0 *1 168.495,5.46
X$754 544 3 545 644 645 cell_1rw
* cell instance $755 m0 *1 169.2,5.46
X$755 546 3 547 644 645 cell_1rw
* cell instance $756 m0 *1 169.905,5.46
X$756 548 3 549 644 645 cell_1rw
* cell instance $757 m0 *1 170.61,5.46
X$757 550 3 551 644 645 cell_1rw
* cell instance $758 m0 *1 171.315,5.46
X$758 552 3 553 644 645 cell_1rw
* cell instance $759 m0 *1 172.02,5.46
X$759 554 3 555 644 645 cell_1rw
* cell instance $760 m0 *1 172.725,5.46
X$760 556 3 557 644 645 cell_1rw
* cell instance $761 m0 *1 173.43,5.46
X$761 558 3 559 644 645 cell_1rw
* cell instance $762 m0 *1 174.135,5.46
X$762 560 3 561 644 645 cell_1rw
* cell instance $763 m0 *1 174.84,5.46
X$763 562 3 563 644 645 cell_1rw
* cell instance $764 m0 *1 175.545,5.46
X$764 564 3 565 644 645 cell_1rw
* cell instance $765 m0 *1 176.25,5.46
X$765 566 3 567 644 645 cell_1rw
* cell instance $766 m0 *1 176.955,5.46
X$766 568 3 569 644 645 cell_1rw
* cell instance $767 m0 *1 177.66,5.46
X$767 570 3 571 644 645 cell_1rw
* cell instance $768 m0 *1 178.365,5.46
X$768 572 3 573 644 645 cell_1rw
* cell instance $769 m0 *1 179.07,5.46
X$769 574 3 575 644 645 cell_1rw
* cell instance $770 m0 *1 179.775,5.46
X$770 576 3 577 644 645 cell_1rw
* cell instance $771 m0 *1 180.48,5.46
X$771 578 3 579 644 645 cell_1rw
* cell instance $772 r0 *1 0.705,2.73
X$772 67 4 68 644 645 cell_1rw
* cell instance $773 r0 *1 0,2.73
X$773 65 4 66 644 645 cell_1rw
* cell instance $774 r0 *1 1.41,2.73
X$774 69 4 70 644 645 cell_1rw
* cell instance $775 r0 *1 2.115,2.73
X$775 71 4 72 644 645 cell_1rw
* cell instance $776 r0 *1 2.82,2.73
X$776 73 4 74 644 645 cell_1rw
* cell instance $777 r0 *1 3.525,2.73
X$777 75 4 76 644 645 cell_1rw
* cell instance $778 r0 *1 4.23,2.73
X$778 77 4 78 644 645 cell_1rw
* cell instance $779 r0 *1 4.935,2.73
X$779 79 4 80 644 645 cell_1rw
* cell instance $780 r0 *1 5.64,2.73
X$780 81 4 82 644 645 cell_1rw
* cell instance $781 r0 *1 6.345,2.73
X$781 83 4 84 644 645 cell_1rw
* cell instance $782 r0 *1 7.05,2.73
X$782 85 4 86 644 645 cell_1rw
* cell instance $783 r0 *1 7.755,2.73
X$783 87 4 88 644 645 cell_1rw
* cell instance $784 r0 *1 8.46,2.73
X$784 89 4 90 644 645 cell_1rw
* cell instance $785 r0 *1 9.165,2.73
X$785 91 4 92 644 645 cell_1rw
* cell instance $786 r0 *1 9.87,2.73
X$786 93 4 94 644 645 cell_1rw
* cell instance $787 r0 *1 10.575,2.73
X$787 95 4 96 644 645 cell_1rw
* cell instance $788 r0 *1 11.28,2.73
X$788 97 4 98 644 645 cell_1rw
* cell instance $789 r0 *1 11.985,2.73
X$789 99 4 100 644 645 cell_1rw
* cell instance $790 r0 *1 12.69,2.73
X$790 101 4 102 644 645 cell_1rw
* cell instance $791 r0 *1 13.395,2.73
X$791 103 4 104 644 645 cell_1rw
* cell instance $792 r0 *1 14.1,2.73
X$792 105 4 106 644 645 cell_1rw
* cell instance $793 r0 *1 14.805,2.73
X$793 107 4 108 644 645 cell_1rw
* cell instance $794 r0 *1 15.51,2.73
X$794 109 4 110 644 645 cell_1rw
* cell instance $795 r0 *1 16.215,2.73
X$795 111 4 112 644 645 cell_1rw
* cell instance $796 r0 *1 16.92,2.73
X$796 113 4 114 644 645 cell_1rw
* cell instance $797 r0 *1 17.625,2.73
X$797 115 4 116 644 645 cell_1rw
* cell instance $798 r0 *1 18.33,2.73
X$798 117 4 118 644 645 cell_1rw
* cell instance $799 r0 *1 19.035,2.73
X$799 119 4 120 644 645 cell_1rw
* cell instance $800 r0 *1 19.74,2.73
X$800 121 4 122 644 645 cell_1rw
* cell instance $801 r0 *1 20.445,2.73
X$801 123 4 124 644 645 cell_1rw
* cell instance $802 r0 *1 21.15,2.73
X$802 125 4 126 644 645 cell_1rw
* cell instance $803 r0 *1 21.855,2.73
X$803 127 4 128 644 645 cell_1rw
* cell instance $804 r0 *1 22.56,2.73
X$804 129 4 130 644 645 cell_1rw
* cell instance $805 r0 *1 23.265,2.73
X$805 131 4 132 644 645 cell_1rw
* cell instance $806 r0 *1 23.97,2.73
X$806 133 4 134 644 645 cell_1rw
* cell instance $807 r0 *1 24.675,2.73
X$807 135 4 136 644 645 cell_1rw
* cell instance $808 r0 *1 25.38,2.73
X$808 137 4 138 644 645 cell_1rw
* cell instance $809 r0 *1 26.085,2.73
X$809 139 4 140 644 645 cell_1rw
* cell instance $810 r0 *1 26.79,2.73
X$810 141 4 142 644 645 cell_1rw
* cell instance $811 r0 *1 27.495,2.73
X$811 143 4 144 644 645 cell_1rw
* cell instance $812 r0 *1 28.2,2.73
X$812 145 4 146 644 645 cell_1rw
* cell instance $813 r0 *1 28.905,2.73
X$813 147 4 148 644 645 cell_1rw
* cell instance $814 r0 *1 29.61,2.73
X$814 149 4 150 644 645 cell_1rw
* cell instance $815 r0 *1 30.315,2.73
X$815 151 4 152 644 645 cell_1rw
* cell instance $816 r0 *1 31.02,2.73
X$816 153 4 154 644 645 cell_1rw
* cell instance $817 r0 *1 31.725,2.73
X$817 155 4 156 644 645 cell_1rw
* cell instance $818 r0 *1 32.43,2.73
X$818 157 4 158 644 645 cell_1rw
* cell instance $819 r0 *1 33.135,2.73
X$819 159 4 160 644 645 cell_1rw
* cell instance $820 r0 *1 33.84,2.73
X$820 161 4 162 644 645 cell_1rw
* cell instance $821 r0 *1 34.545,2.73
X$821 163 4 164 644 645 cell_1rw
* cell instance $822 r0 *1 35.25,2.73
X$822 165 4 166 644 645 cell_1rw
* cell instance $823 r0 *1 35.955,2.73
X$823 167 4 168 644 645 cell_1rw
* cell instance $824 r0 *1 36.66,2.73
X$824 169 4 170 644 645 cell_1rw
* cell instance $825 r0 *1 37.365,2.73
X$825 171 4 172 644 645 cell_1rw
* cell instance $826 r0 *1 38.07,2.73
X$826 173 4 174 644 645 cell_1rw
* cell instance $827 r0 *1 38.775,2.73
X$827 175 4 176 644 645 cell_1rw
* cell instance $828 r0 *1 39.48,2.73
X$828 177 4 178 644 645 cell_1rw
* cell instance $829 r0 *1 40.185,2.73
X$829 179 4 180 644 645 cell_1rw
* cell instance $830 r0 *1 40.89,2.73
X$830 181 4 182 644 645 cell_1rw
* cell instance $831 r0 *1 41.595,2.73
X$831 183 4 184 644 645 cell_1rw
* cell instance $832 r0 *1 42.3,2.73
X$832 185 4 186 644 645 cell_1rw
* cell instance $833 r0 *1 43.005,2.73
X$833 187 4 188 644 645 cell_1rw
* cell instance $834 r0 *1 43.71,2.73
X$834 189 4 190 644 645 cell_1rw
* cell instance $835 r0 *1 44.415,2.73
X$835 191 4 192 644 645 cell_1rw
* cell instance $836 r0 *1 45.12,2.73
X$836 193 4 194 644 645 cell_1rw
* cell instance $837 r0 *1 45.825,2.73
X$837 195 4 196 644 645 cell_1rw
* cell instance $838 r0 *1 46.53,2.73
X$838 197 4 198 644 645 cell_1rw
* cell instance $839 r0 *1 47.235,2.73
X$839 199 4 200 644 645 cell_1rw
* cell instance $840 r0 *1 47.94,2.73
X$840 201 4 202 644 645 cell_1rw
* cell instance $841 r0 *1 48.645,2.73
X$841 203 4 204 644 645 cell_1rw
* cell instance $842 r0 *1 49.35,2.73
X$842 205 4 206 644 645 cell_1rw
* cell instance $843 r0 *1 50.055,2.73
X$843 207 4 208 644 645 cell_1rw
* cell instance $844 r0 *1 50.76,2.73
X$844 209 4 210 644 645 cell_1rw
* cell instance $845 r0 *1 51.465,2.73
X$845 211 4 212 644 645 cell_1rw
* cell instance $846 r0 *1 52.17,2.73
X$846 213 4 214 644 645 cell_1rw
* cell instance $847 r0 *1 52.875,2.73
X$847 215 4 216 644 645 cell_1rw
* cell instance $848 r0 *1 53.58,2.73
X$848 217 4 218 644 645 cell_1rw
* cell instance $849 r0 *1 54.285,2.73
X$849 219 4 220 644 645 cell_1rw
* cell instance $850 r0 *1 54.99,2.73
X$850 221 4 222 644 645 cell_1rw
* cell instance $851 r0 *1 55.695,2.73
X$851 223 4 224 644 645 cell_1rw
* cell instance $852 r0 *1 56.4,2.73
X$852 225 4 226 644 645 cell_1rw
* cell instance $853 r0 *1 57.105,2.73
X$853 227 4 228 644 645 cell_1rw
* cell instance $854 r0 *1 57.81,2.73
X$854 229 4 230 644 645 cell_1rw
* cell instance $855 r0 *1 58.515,2.73
X$855 231 4 232 644 645 cell_1rw
* cell instance $856 r0 *1 59.22,2.73
X$856 233 4 234 644 645 cell_1rw
* cell instance $857 r0 *1 59.925,2.73
X$857 235 4 236 644 645 cell_1rw
* cell instance $858 r0 *1 60.63,2.73
X$858 237 4 238 644 645 cell_1rw
* cell instance $859 r0 *1 61.335,2.73
X$859 239 4 240 644 645 cell_1rw
* cell instance $860 r0 *1 62.04,2.73
X$860 241 4 242 644 645 cell_1rw
* cell instance $861 r0 *1 62.745,2.73
X$861 243 4 244 644 645 cell_1rw
* cell instance $862 r0 *1 63.45,2.73
X$862 245 4 246 644 645 cell_1rw
* cell instance $863 r0 *1 64.155,2.73
X$863 247 4 248 644 645 cell_1rw
* cell instance $864 r0 *1 64.86,2.73
X$864 249 4 250 644 645 cell_1rw
* cell instance $865 r0 *1 65.565,2.73
X$865 251 4 252 644 645 cell_1rw
* cell instance $866 r0 *1 66.27,2.73
X$866 253 4 254 644 645 cell_1rw
* cell instance $867 r0 *1 66.975,2.73
X$867 255 4 256 644 645 cell_1rw
* cell instance $868 r0 *1 67.68,2.73
X$868 257 4 258 644 645 cell_1rw
* cell instance $869 r0 *1 68.385,2.73
X$869 259 4 260 644 645 cell_1rw
* cell instance $870 r0 *1 69.09,2.73
X$870 261 4 262 644 645 cell_1rw
* cell instance $871 r0 *1 69.795,2.73
X$871 263 4 264 644 645 cell_1rw
* cell instance $872 r0 *1 70.5,2.73
X$872 265 4 266 644 645 cell_1rw
* cell instance $873 r0 *1 71.205,2.73
X$873 267 4 268 644 645 cell_1rw
* cell instance $874 r0 *1 71.91,2.73
X$874 269 4 270 644 645 cell_1rw
* cell instance $875 r0 *1 72.615,2.73
X$875 271 4 272 644 645 cell_1rw
* cell instance $876 r0 *1 73.32,2.73
X$876 273 4 274 644 645 cell_1rw
* cell instance $877 r0 *1 74.025,2.73
X$877 275 4 276 644 645 cell_1rw
* cell instance $878 r0 *1 74.73,2.73
X$878 277 4 278 644 645 cell_1rw
* cell instance $879 r0 *1 75.435,2.73
X$879 279 4 280 644 645 cell_1rw
* cell instance $880 r0 *1 76.14,2.73
X$880 281 4 282 644 645 cell_1rw
* cell instance $881 r0 *1 76.845,2.73
X$881 283 4 284 644 645 cell_1rw
* cell instance $882 r0 *1 77.55,2.73
X$882 285 4 286 644 645 cell_1rw
* cell instance $883 r0 *1 78.255,2.73
X$883 287 4 288 644 645 cell_1rw
* cell instance $884 r0 *1 78.96,2.73
X$884 289 4 290 644 645 cell_1rw
* cell instance $885 r0 *1 79.665,2.73
X$885 291 4 292 644 645 cell_1rw
* cell instance $886 r0 *1 80.37,2.73
X$886 293 4 294 644 645 cell_1rw
* cell instance $887 r0 *1 81.075,2.73
X$887 295 4 296 644 645 cell_1rw
* cell instance $888 r0 *1 81.78,2.73
X$888 297 4 298 644 645 cell_1rw
* cell instance $889 r0 *1 82.485,2.73
X$889 299 4 300 644 645 cell_1rw
* cell instance $890 r0 *1 83.19,2.73
X$890 301 4 302 644 645 cell_1rw
* cell instance $891 r0 *1 83.895,2.73
X$891 303 4 304 644 645 cell_1rw
* cell instance $892 r0 *1 84.6,2.73
X$892 305 4 306 644 645 cell_1rw
* cell instance $893 r0 *1 85.305,2.73
X$893 307 4 308 644 645 cell_1rw
* cell instance $894 r0 *1 86.01,2.73
X$894 309 4 310 644 645 cell_1rw
* cell instance $895 r0 *1 86.715,2.73
X$895 311 4 312 644 645 cell_1rw
* cell instance $896 r0 *1 87.42,2.73
X$896 313 4 314 644 645 cell_1rw
* cell instance $897 r0 *1 88.125,2.73
X$897 315 4 316 644 645 cell_1rw
* cell instance $898 r0 *1 88.83,2.73
X$898 317 4 318 644 645 cell_1rw
* cell instance $899 r0 *1 89.535,2.73
X$899 319 4 320 644 645 cell_1rw
* cell instance $900 r0 *1 90.24,2.73
X$900 321 4 323 644 645 cell_1rw
* cell instance $901 r0 *1 90.945,2.73
X$901 324 4 325 644 645 cell_1rw
* cell instance $902 r0 *1 91.65,2.73
X$902 326 4 327 644 645 cell_1rw
* cell instance $903 r0 *1 92.355,2.73
X$903 328 4 329 644 645 cell_1rw
* cell instance $904 r0 *1 93.06,2.73
X$904 330 4 331 644 645 cell_1rw
* cell instance $905 r0 *1 93.765,2.73
X$905 332 4 333 644 645 cell_1rw
* cell instance $906 r0 *1 94.47,2.73
X$906 334 4 335 644 645 cell_1rw
* cell instance $907 r0 *1 95.175,2.73
X$907 336 4 337 644 645 cell_1rw
* cell instance $908 r0 *1 95.88,2.73
X$908 338 4 339 644 645 cell_1rw
* cell instance $909 r0 *1 96.585,2.73
X$909 340 4 341 644 645 cell_1rw
* cell instance $910 r0 *1 97.29,2.73
X$910 342 4 343 644 645 cell_1rw
* cell instance $911 r0 *1 97.995,2.73
X$911 344 4 345 644 645 cell_1rw
* cell instance $912 r0 *1 98.7,2.73
X$912 346 4 347 644 645 cell_1rw
* cell instance $913 r0 *1 99.405,2.73
X$913 348 4 349 644 645 cell_1rw
* cell instance $914 r0 *1 100.11,2.73
X$914 350 4 351 644 645 cell_1rw
* cell instance $915 r0 *1 100.815,2.73
X$915 352 4 353 644 645 cell_1rw
* cell instance $916 r0 *1 101.52,2.73
X$916 354 4 355 644 645 cell_1rw
* cell instance $917 r0 *1 102.225,2.73
X$917 356 4 357 644 645 cell_1rw
* cell instance $918 r0 *1 102.93,2.73
X$918 358 4 359 644 645 cell_1rw
* cell instance $919 r0 *1 103.635,2.73
X$919 360 4 361 644 645 cell_1rw
* cell instance $920 r0 *1 104.34,2.73
X$920 362 4 363 644 645 cell_1rw
* cell instance $921 r0 *1 105.045,2.73
X$921 364 4 365 644 645 cell_1rw
* cell instance $922 r0 *1 105.75,2.73
X$922 366 4 367 644 645 cell_1rw
* cell instance $923 r0 *1 106.455,2.73
X$923 368 4 369 644 645 cell_1rw
* cell instance $924 r0 *1 107.16,2.73
X$924 370 4 371 644 645 cell_1rw
* cell instance $925 r0 *1 107.865,2.73
X$925 372 4 373 644 645 cell_1rw
* cell instance $926 r0 *1 108.57,2.73
X$926 374 4 375 644 645 cell_1rw
* cell instance $927 r0 *1 109.275,2.73
X$927 376 4 377 644 645 cell_1rw
* cell instance $928 r0 *1 109.98,2.73
X$928 378 4 379 644 645 cell_1rw
* cell instance $929 r0 *1 110.685,2.73
X$929 380 4 381 644 645 cell_1rw
* cell instance $930 r0 *1 111.39,2.73
X$930 382 4 383 644 645 cell_1rw
* cell instance $931 r0 *1 112.095,2.73
X$931 384 4 385 644 645 cell_1rw
* cell instance $932 r0 *1 112.8,2.73
X$932 386 4 387 644 645 cell_1rw
* cell instance $933 r0 *1 113.505,2.73
X$933 388 4 389 644 645 cell_1rw
* cell instance $934 r0 *1 114.21,2.73
X$934 390 4 391 644 645 cell_1rw
* cell instance $935 r0 *1 114.915,2.73
X$935 392 4 393 644 645 cell_1rw
* cell instance $936 r0 *1 115.62,2.73
X$936 394 4 395 644 645 cell_1rw
* cell instance $937 r0 *1 116.325,2.73
X$937 396 4 397 644 645 cell_1rw
* cell instance $938 r0 *1 117.03,2.73
X$938 398 4 399 644 645 cell_1rw
* cell instance $939 r0 *1 117.735,2.73
X$939 400 4 401 644 645 cell_1rw
* cell instance $940 r0 *1 118.44,2.73
X$940 402 4 403 644 645 cell_1rw
* cell instance $941 r0 *1 119.145,2.73
X$941 404 4 405 644 645 cell_1rw
* cell instance $942 r0 *1 119.85,2.73
X$942 406 4 407 644 645 cell_1rw
* cell instance $943 r0 *1 120.555,2.73
X$943 408 4 409 644 645 cell_1rw
* cell instance $944 r0 *1 121.26,2.73
X$944 410 4 411 644 645 cell_1rw
* cell instance $945 r0 *1 121.965,2.73
X$945 412 4 413 644 645 cell_1rw
* cell instance $946 r0 *1 122.67,2.73
X$946 414 4 415 644 645 cell_1rw
* cell instance $947 r0 *1 123.375,2.73
X$947 416 4 417 644 645 cell_1rw
* cell instance $948 r0 *1 124.08,2.73
X$948 418 4 419 644 645 cell_1rw
* cell instance $949 r0 *1 124.785,2.73
X$949 420 4 421 644 645 cell_1rw
* cell instance $950 r0 *1 125.49,2.73
X$950 422 4 423 644 645 cell_1rw
* cell instance $951 r0 *1 126.195,2.73
X$951 424 4 425 644 645 cell_1rw
* cell instance $952 r0 *1 126.9,2.73
X$952 426 4 427 644 645 cell_1rw
* cell instance $953 r0 *1 127.605,2.73
X$953 428 4 429 644 645 cell_1rw
* cell instance $954 r0 *1 128.31,2.73
X$954 430 4 431 644 645 cell_1rw
* cell instance $955 r0 *1 129.015,2.73
X$955 432 4 433 644 645 cell_1rw
* cell instance $956 r0 *1 129.72,2.73
X$956 434 4 435 644 645 cell_1rw
* cell instance $957 r0 *1 130.425,2.73
X$957 436 4 437 644 645 cell_1rw
* cell instance $958 r0 *1 131.13,2.73
X$958 438 4 439 644 645 cell_1rw
* cell instance $959 r0 *1 131.835,2.73
X$959 440 4 441 644 645 cell_1rw
* cell instance $960 r0 *1 132.54,2.73
X$960 442 4 443 644 645 cell_1rw
* cell instance $961 r0 *1 133.245,2.73
X$961 444 4 445 644 645 cell_1rw
* cell instance $962 r0 *1 133.95,2.73
X$962 446 4 447 644 645 cell_1rw
* cell instance $963 r0 *1 134.655,2.73
X$963 448 4 449 644 645 cell_1rw
* cell instance $964 r0 *1 135.36,2.73
X$964 450 4 451 644 645 cell_1rw
* cell instance $965 r0 *1 136.065,2.73
X$965 452 4 453 644 645 cell_1rw
* cell instance $966 r0 *1 136.77,2.73
X$966 454 4 455 644 645 cell_1rw
* cell instance $967 r0 *1 137.475,2.73
X$967 456 4 457 644 645 cell_1rw
* cell instance $968 r0 *1 138.18,2.73
X$968 458 4 459 644 645 cell_1rw
* cell instance $969 r0 *1 138.885,2.73
X$969 460 4 461 644 645 cell_1rw
* cell instance $970 r0 *1 139.59,2.73
X$970 462 4 463 644 645 cell_1rw
* cell instance $971 r0 *1 140.295,2.73
X$971 464 4 465 644 645 cell_1rw
* cell instance $972 r0 *1 141,2.73
X$972 466 4 467 644 645 cell_1rw
* cell instance $973 r0 *1 141.705,2.73
X$973 468 4 469 644 645 cell_1rw
* cell instance $974 r0 *1 142.41,2.73
X$974 470 4 471 644 645 cell_1rw
* cell instance $975 r0 *1 143.115,2.73
X$975 472 4 473 644 645 cell_1rw
* cell instance $976 r0 *1 143.82,2.73
X$976 474 4 475 644 645 cell_1rw
* cell instance $977 r0 *1 144.525,2.73
X$977 476 4 477 644 645 cell_1rw
* cell instance $978 r0 *1 145.23,2.73
X$978 478 4 479 644 645 cell_1rw
* cell instance $979 r0 *1 145.935,2.73
X$979 480 4 481 644 645 cell_1rw
* cell instance $980 r0 *1 146.64,2.73
X$980 482 4 483 644 645 cell_1rw
* cell instance $981 r0 *1 147.345,2.73
X$981 484 4 485 644 645 cell_1rw
* cell instance $982 r0 *1 148.05,2.73
X$982 486 4 487 644 645 cell_1rw
* cell instance $983 r0 *1 148.755,2.73
X$983 488 4 489 644 645 cell_1rw
* cell instance $984 r0 *1 149.46,2.73
X$984 490 4 491 644 645 cell_1rw
* cell instance $985 r0 *1 150.165,2.73
X$985 492 4 493 644 645 cell_1rw
* cell instance $986 r0 *1 150.87,2.73
X$986 494 4 495 644 645 cell_1rw
* cell instance $987 r0 *1 151.575,2.73
X$987 496 4 497 644 645 cell_1rw
* cell instance $988 r0 *1 152.28,2.73
X$988 498 4 499 644 645 cell_1rw
* cell instance $989 r0 *1 152.985,2.73
X$989 500 4 501 644 645 cell_1rw
* cell instance $990 r0 *1 153.69,2.73
X$990 502 4 503 644 645 cell_1rw
* cell instance $991 r0 *1 154.395,2.73
X$991 504 4 505 644 645 cell_1rw
* cell instance $992 r0 *1 155.1,2.73
X$992 506 4 507 644 645 cell_1rw
* cell instance $993 r0 *1 155.805,2.73
X$993 508 4 509 644 645 cell_1rw
* cell instance $994 r0 *1 156.51,2.73
X$994 510 4 511 644 645 cell_1rw
* cell instance $995 r0 *1 157.215,2.73
X$995 512 4 513 644 645 cell_1rw
* cell instance $996 r0 *1 157.92,2.73
X$996 514 4 515 644 645 cell_1rw
* cell instance $997 r0 *1 158.625,2.73
X$997 516 4 517 644 645 cell_1rw
* cell instance $998 r0 *1 159.33,2.73
X$998 518 4 519 644 645 cell_1rw
* cell instance $999 r0 *1 160.035,2.73
X$999 520 4 521 644 645 cell_1rw
* cell instance $1000 r0 *1 160.74,2.73
X$1000 522 4 523 644 645 cell_1rw
* cell instance $1001 r0 *1 161.445,2.73
X$1001 524 4 525 644 645 cell_1rw
* cell instance $1002 r0 *1 162.15,2.73
X$1002 526 4 527 644 645 cell_1rw
* cell instance $1003 r0 *1 162.855,2.73
X$1003 528 4 529 644 645 cell_1rw
* cell instance $1004 r0 *1 163.56,2.73
X$1004 530 4 531 644 645 cell_1rw
* cell instance $1005 r0 *1 164.265,2.73
X$1005 532 4 533 644 645 cell_1rw
* cell instance $1006 r0 *1 164.97,2.73
X$1006 534 4 535 644 645 cell_1rw
* cell instance $1007 r0 *1 165.675,2.73
X$1007 536 4 537 644 645 cell_1rw
* cell instance $1008 r0 *1 166.38,2.73
X$1008 538 4 539 644 645 cell_1rw
* cell instance $1009 r0 *1 167.085,2.73
X$1009 540 4 541 644 645 cell_1rw
* cell instance $1010 r0 *1 167.79,2.73
X$1010 542 4 543 644 645 cell_1rw
* cell instance $1011 r0 *1 168.495,2.73
X$1011 544 4 545 644 645 cell_1rw
* cell instance $1012 r0 *1 169.2,2.73
X$1012 546 4 547 644 645 cell_1rw
* cell instance $1013 r0 *1 169.905,2.73
X$1013 548 4 549 644 645 cell_1rw
* cell instance $1014 r0 *1 170.61,2.73
X$1014 550 4 551 644 645 cell_1rw
* cell instance $1015 r0 *1 171.315,2.73
X$1015 552 4 553 644 645 cell_1rw
* cell instance $1016 r0 *1 172.02,2.73
X$1016 554 4 555 644 645 cell_1rw
* cell instance $1017 r0 *1 172.725,2.73
X$1017 556 4 557 644 645 cell_1rw
* cell instance $1018 r0 *1 173.43,2.73
X$1018 558 4 559 644 645 cell_1rw
* cell instance $1019 r0 *1 174.135,2.73
X$1019 560 4 561 644 645 cell_1rw
* cell instance $1020 r0 *1 174.84,2.73
X$1020 562 4 563 644 645 cell_1rw
* cell instance $1021 r0 *1 175.545,2.73
X$1021 564 4 565 644 645 cell_1rw
* cell instance $1022 r0 *1 176.25,2.73
X$1022 566 4 567 644 645 cell_1rw
* cell instance $1023 r0 *1 176.955,2.73
X$1023 568 4 569 644 645 cell_1rw
* cell instance $1024 r0 *1 177.66,2.73
X$1024 570 4 571 644 645 cell_1rw
* cell instance $1025 r0 *1 178.365,2.73
X$1025 572 4 573 644 645 cell_1rw
* cell instance $1026 r0 *1 179.07,2.73
X$1026 574 4 575 644 645 cell_1rw
* cell instance $1027 r0 *1 179.775,2.73
X$1027 576 4 577 644 645 cell_1rw
* cell instance $1028 r0 *1 180.48,2.73
X$1028 578 4 579 644 645 cell_1rw
* cell instance $1029 r0 *1 0.705,5.46
X$1029 67 5 68 644 645 cell_1rw
* cell instance $1030 r0 *1 0,5.46
X$1030 65 5 66 644 645 cell_1rw
* cell instance $1031 r0 *1 1.41,5.46
X$1031 69 5 70 644 645 cell_1rw
* cell instance $1032 r0 *1 2.115,5.46
X$1032 71 5 72 644 645 cell_1rw
* cell instance $1033 r0 *1 2.82,5.46
X$1033 73 5 74 644 645 cell_1rw
* cell instance $1034 r0 *1 3.525,5.46
X$1034 75 5 76 644 645 cell_1rw
* cell instance $1035 r0 *1 4.23,5.46
X$1035 77 5 78 644 645 cell_1rw
* cell instance $1036 r0 *1 4.935,5.46
X$1036 79 5 80 644 645 cell_1rw
* cell instance $1037 r0 *1 5.64,5.46
X$1037 81 5 82 644 645 cell_1rw
* cell instance $1038 r0 *1 6.345,5.46
X$1038 83 5 84 644 645 cell_1rw
* cell instance $1039 r0 *1 7.05,5.46
X$1039 85 5 86 644 645 cell_1rw
* cell instance $1040 r0 *1 7.755,5.46
X$1040 87 5 88 644 645 cell_1rw
* cell instance $1041 r0 *1 8.46,5.46
X$1041 89 5 90 644 645 cell_1rw
* cell instance $1042 r0 *1 9.165,5.46
X$1042 91 5 92 644 645 cell_1rw
* cell instance $1043 r0 *1 9.87,5.46
X$1043 93 5 94 644 645 cell_1rw
* cell instance $1044 r0 *1 10.575,5.46
X$1044 95 5 96 644 645 cell_1rw
* cell instance $1045 r0 *1 11.28,5.46
X$1045 97 5 98 644 645 cell_1rw
* cell instance $1046 r0 *1 11.985,5.46
X$1046 99 5 100 644 645 cell_1rw
* cell instance $1047 r0 *1 12.69,5.46
X$1047 101 5 102 644 645 cell_1rw
* cell instance $1048 r0 *1 13.395,5.46
X$1048 103 5 104 644 645 cell_1rw
* cell instance $1049 r0 *1 14.1,5.46
X$1049 105 5 106 644 645 cell_1rw
* cell instance $1050 r0 *1 14.805,5.46
X$1050 107 5 108 644 645 cell_1rw
* cell instance $1051 r0 *1 15.51,5.46
X$1051 109 5 110 644 645 cell_1rw
* cell instance $1052 r0 *1 16.215,5.46
X$1052 111 5 112 644 645 cell_1rw
* cell instance $1053 r0 *1 16.92,5.46
X$1053 113 5 114 644 645 cell_1rw
* cell instance $1054 r0 *1 17.625,5.46
X$1054 115 5 116 644 645 cell_1rw
* cell instance $1055 r0 *1 18.33,5.46
X$1055 117 5 118 644 645 cell_1rw
* cell instance $1056 r0 *1 19.035,5.46
X$1056 119 5 120 644 645 cell_1rw
* cell instance $1057 r0 *1 19.74,5.46
X$1057 121 5 122 644 645 cell_1rw
* cell instance $1058 r0 *1 20.445,5.46
X$1058 123 5 124 644 645 cell_1rw
* cell instance $1059 r0 *1 21.15,5.46
X$1059 125 5 126 644 645 cell_1rw
* cell instance $1060 r0 *1 21.855,5.46
X$1060 127 5 128 644 645 cell_1rw
* cell instance $1061 r0 *1 22.56,5.46
X$1061 129 5 130 644 645 cell_1rw
* cell instance $1062 r0 *1 23.265,5.46
X$1062 131 5 132 644 645 cell_1rw
* cell instance $1063 r0 *1 23.97,5.46
X$1063 133 5 134 644 645 cell_1rw
* cell instance $1064 r0 *1 24.675,5.46
X$1064 135 5 136 644 645 cell_1rw
* cell instance $1065 r0 *1 25.38,5.46
X$1065 137 5 138 644 645 cell_1rw
* cell instance $1066 r0 *1 26.085,5.46
X$1066 139 5 140 644 645 cell_1rw
* cell instance $1067 r0 *1 26.79,5.46
X$1067 141 5 142 644 645 cell_1rw
* cell instance $1068 r0 *1 27.495,5.46
X$1068 143 5 144 644 645 cell_1rw
* cell instance $1069 r0 *1 28.2,5.46
X$1069 145 5 146 644 645 cell_1rw
* cell instance $1070 r0 *1 28.905,5.46
X$1070 147 5 148 644 645 cell_1rw
* cell instance $1071 r0 *1 29.61,5.46
X$1071 149 5 150 644 645 cell_1rw
* cell instance $1072 r0 *1 30.315,5.46
X$1072 151 5 152 644 645 cell_1rw
* cell instance $1073 r0 *1 31.02,5.46
X$1073 153 5 154 644 645 cell_1rw
* cell instance $1074 r0 *1 31.725,5.46
X$1074 155 5 156 644 645 cell_1rw
* cell instance $1075 r0 *1 32.43,5.46
X$1075 157 5 158 644 645 cell_1rw
* cell instance $1076 r0 *1 33.135,5.46
X$1076 159 5 160 644 645 cell_1rw
* cell instance $1077 r0 *1 33.84,5.46
X$1077 161 5 162 644 645 cell_1rw
* cell instance $1078 r0 *1 34.545,5.46
X$1078 163 5 164 644 645 cell_1rw
* cell instance $1079 r0 *1 35.25,5.46
X$1079 165 5 166 644 645 cell_1rw
* cell instance $1080 r0 *1 35.955,5.46
X$1080 167 5 168 644 645 cell_1rw
* cell instance $1081 r0 *1 36.66,5.46
X$1081 169 5 170 644 645 cell_1rw
* cell instance $1082 r0 *1 37.365,5.46
X$1082 171 5 172 644 645 cell_1rw
* cell instance $1083 r0 *1 38.07,5.46
X$1083 173 5 174 644 645 cell_1rw
* cell instance $1084 r0 *1 38.775,5.46
X$1084 175 5 176 644 645 cell_1rw
* cell instance $1085 r0 *1 39.48,5.46
X$1085 177 5 178 644 645 cell_1rw
* cell instance $1086 r0 *1 40.185,5.46
X$1086 179 5 180 644 645 cell_1rw
* cell instance $1087 r0 *1 40.89,5.46
X$1087 181 5 182 644 645 cell_1rw
* cell instance $1088 r0 *1 41.595,5.46
X$1088 183 5 184 644 645 cell_1rw
* cell instance $1089 r0 *1 42.3,5.46
X$1089 185 5 186 644 645 cell_1rw
* cell instance $1090 r0 *1 43.005,5.46
X$1090 187 5 188 644 645 cell_1rw
* cell instance $1091 r0 *1 43.71,5.46
X$1091 189 5 190 644 645 cell_1rw
* cell instance $1092 r0 *1 44.415,5.46
X$1092 191 5 192 644 645 cell_1rw
* cell instance $1093 r0 *1 45.12,5.46
X$1093 193 5 194 644 645 cell_1rw
* cell instance $1094 r0 *1 45.825,5.46
X$1094 195 5 196 644 645 cell_1rw
* cell instance $1095 r0 *1 46.53,5.46
X$1095 197 5 198 644 645 cell_1rw
* cell instance $1096 r0 *1 47.235,5.46
X$1096 199 5 200 644 645 cell_1rw
* cell instance $1097 r0 *1 47.94,5.46
X$1097 201 5 202 644 645 cell_1rw
* cell instance $1098 r0 *1 48.645,5.46
X$1098 203 5 204 644 645 cell_1rw
* cell instance $1099 r0 *1 49.35,5.46
X$1099 205 5 206 644 645 cell_1rw
* cell instance $1100 r0 *1 50.055,5.46
X$1100 207 5 208 644 645 cell_1rw
* cell instance $1101 r0 *1 50.76,5.46
X$1101 209 5 210 644 645 cell_1rw
* cell instance $1102 r0 *1 51.465,5.46
X$1102 211 5 212 644 645 cell_1rw
* cell instance $1103 r0 *1 52.17,5.46
X$1103 213 5 214 644 645 cell_1rw
* cell instance $1104 r0 *1 52.875,5.46
X$1104 215 5 216 644 645 cell_1rw
* cell instance $1105 r0 *1 53.58,5.46
X$1105 217 5 218 644 645 cell_1rw
* cell instance $1106 r0 *1 54.285,5.46
X$1106 219 5 220 644 645 cell_1rw
* cell instance $1107 r0 *1 54.99,5.46
X$1107 221 5 222 644 645 cell_1rw
* cell instance $1108 r0 *1 55.695,5.46
X$1108 223 5 224 644 645 cell_1rw
* cell instance $1109 r0 *1 56.4,5.46
X$1109 225 5 226 644 645 cell_1rw
* cell instance $1110 r0 *1 57.105,5.46
X$1110 227 5 228 644 645 cell_1rw
* cell instance $1111 r0 *1 57.81,5.46
X$1111 229 5 230 644 645 cell_1rw
* cell instance $1112 r0 *1 58.515,5.46
X$1112 231 5 232 644 645 cell_1rw
* cell instance $1113 r0 *1 59.22,5.46
X$1113 233 5 234 644 645 cell_1rw
* cell instance $1114 r0 *1 59.925,5.46
X$1114 235 5 236 644 645 cell_1rw
* cell instance $1115 r0 *1 60.63,5.46
X$1115 237 5 238 644 645 cell_1rw
* cell instance $1116 r0 *1 61.335,5.46
X$1116 239 5 240 644 645 cell_1rw
* cell instance $1117 r0 *1 62.04,5.46
X$1117 241 5 242 644 645 cell_1rw
* cell instance $1118 r0 *1 62.745,5.46
X$1118 243 5 244 644 645 cell_1rw
* cell instance $1119 r0 *1 63.45,5.46
X$1119 245 5 246 644 645 cell_1rw
* cell instance $1120 r0 *1 64.155,5.46
X$1120 247 5 248 644 645 cell_1rw
* cell instance $1121 r0 *1 64.86,5.46
X$1121 249 5 250 644 645 cell_1rw
* cell instance $1122 r0 *1 65.565,5.46
X$1122 251 5 252 644 645 cell_1rw
* cell instance $1123 r0 *1 66.27,5.46
X$1123 253 5 254 644 645 cell_1rw
* cell instance $1124 r0 *1 66.975,5.46
X$1124 255 5 256 644 645 cell_1rw
* cell instance $1125 r0 *1 67.68,5.46
X$1125 257 5 258 644 645 cell_1rw
* cell instance $1126 r0 *1 68.385,5.46
X$1126 259 5 260 644 645 cell_1rw
* cell instance $1127 r0 *1 69.09,5.46
X$1127 261 5 262 644 645 cell_1rw
* cell instance $1128 r0 *1 69.795,5.46
X$1128 263 5 264 644 645 cell_1rw
* cell instance $1129 r0 *1 70.5,5.46
X$1129 265 5 266 644 645 cell_1rw
* cell instance $1130 r0 *1 71.205,5.46
X$1130 267 5 268 644 645 cell_1rw
* cell instance $1131 r0 *1 71.91,5.46
X$1131 269 5 270 644 645 cell_1rw
* cell instance $1132 r0 *1 72.615,5.46
X$1132 271 5 272 644 645 cell_1rw
* cell instance $1133 r0 *1 73.32,5.46
X$1133 273 5 274 644 645 cell_1rw
* cell instance $1134 r0 *1 74.025,5.46
X$1134 275 5 276 644 645 cell_1rw
* cell instance $1135 r0 *1 74.73,5.46
X$1135 277 5 278 644 645 cell_1rw
* cell instance $1136 r0 *1 75.435,5.46
X$1136 279 5 280 644 645 cell_1rw
* cell instance $1137 r0 *1 76.14,5.46
X$1137 281 5 282 644 645 cell_1rw
* cell instance $1138 r0 *1 76.845,5.46
X$1138 283 5 284 644 645 cell_1rw
* cell instance $1139 r0 *1 77.55,5.46
X$1139 285 5 286 644 645 cell_1rw
* cell instance $1140 r0 *1 78.255,5.46
X$1140 287 5 288 644 645 cell_1rw
* cell instance $1141 r0 *1 78.96,5.46
X$1141 289 5 290 644 645 cell_1rw
* cell instance $1142 r0 *1 79.665,5.46
X$1142 291 5 292 644 645 cell_1rw
* cell instance $1143 r0 *1 80.37,5.46
X$1143 293 5 294 644 645 cell_1rw
* cell instance $1144 r0 *1 81.075,5.46
X$1144 295 5 296 644 645 cell_1rw
* cell instance $1145 r0 *1 81.78,5.46
X$1145 297 5 298 644 645 cell_1rw
* cell instance $1146 r0 *1 82.485,5.46
X$1146 299 5 300 644 645 cell_1rw
* cell instance $1147 r0 *1 83.19,5.46
X$1147 301 5 302 644 645 cell_1rw
* cell instance $1148 r0 *1 83.895,5.46
X$1148 303 5 304 644 645 cell_1rw
* cell instance $1149 r0 *1 84.6,5.46
X$1149 305 5 306 644 645 cell_1rw
* cell instance $1150 r0 *1 85.305,5.46
X$1150 307 5 308 644 645 cell_1rw
* cell instance $1151 r0 *1 86.01,5.46
X$1151 309 5 310 644 645 cell_1rw
* cell instance $1152 r0 *1 86.715,5.46
X$1152 311 5 312 644 645 cell_1rw
* cell instance $1153 r0 *1 87.42,5.46
X$1153 313 5 314 644 645 cell_1rw
* cell instance $1154 r0 *1 88.125,5.46
X$1154 315 5 316 644 645 cell_1rw
* cell instance $1155 r0 *1 88.83,5.46
X$1155 317 5 318 644 645 cell_1rw
* cell instance $1156 r0 *1 89.535,5.46
X$1156 319 5 320 644 645 cell_1rw
* cell instance $1157 r0 *1 90.24,5.46
X$1157 321 5 323 644 645 cell_1rw
* cell instance $1158 r0 *1 90.945,5.46
X$1158 324 5 325 644 645 cell_1rw
* cell instance $1159 r0 *1 91.65,5.46
X$1159 326 5 327 644 645 cell_1rw
* cell instance $1160 r0 *1 92.355,5.46
X$1160 328 5 329 644 645 cell_1rw
* cell instance $1161 r0 *1 93.06,5.46
X$1161 330 5 331 644 645 cell_1rw
* cell instance $1162 r0 *1 93.765,5.46
X$1162 332 5 333 644 645 cell_1rw
* cell instance $1163 r0 *1 94.47,5.46
X$1163 334 5 335 644 645 cell_1rw
* cell instance $1164 r0 *1 95.175,5.46
X$1164 336 5 337 644 645 cell_1rw
* cell instance $1165 r0 *1 95.88,5.46
X$1165 338 5 339 644 645 cell_1rw
* cell instance $1166 r0 *1 96.585,5.46
X$1166 340 5 341 644 645 cell_1rw
* cell instance $1167 r0 *1 97.29,5.46
X$1167 342 5 343 644 645 cell_1rw
* cell instance $1168 r0 *1 97.995,5.46
X$1168 344 5 345 644 645 cell_1rw
* cell instance $1169 r0 *1 98.7,5.46
X$1169 346 5 347 644 645 cell_1rw
* cell instance $1170 r0 *1 99.405,5.46
X$1170 348 5 349 644 645 cell_1rw
* cell instance $1171 r0 *1 100.11,5.46
X$1171 350 5 351 644 645 cell_1rw
* cell instance $1172 r0 *1 100.815,5.46
X$1172 352 5 353 644 645 cell_1rw
* cell instance $1173 r0 *1 101.52,5.46
X$1173 354 5 355 644 645 cell_1rw
* cell instance $1174 r0 *1 102.225,5.46
X$1174 356 5 357 644 645 cell_1rw
* cell instance $1175 r0 *1 102.93,5.46
X$1175 358 5 359 644 645 cell_1rw
* cell instance $1176 r0 *1 103.635,5.46
X$1176 360 5 361 644 645 cell_1rw
* cell instance $1177 r0 *1 104.34,5.46
X$1177 362 5 363 644 645 cell_1rw
* cell instance $1178 r0 *1 105.045,5.46
X$1178 364 5 365 644 645 cell_1rw
* cell instance $1179 r0 *1 105.75,5.46
X$1179 366 5 367 644 645 cell_1rw
* cell instance $1180 r0 *1 106.455,5.46
X$1180 368 5 369 644 645 cell_1rw
* cell instance $1181 r0 *1 107.16,5.46
X$1181 370 5 371 644 645 cell_1rw
* cell instance $1182 r0 *1 107.865,5.46
X$1182 372 5 373 644 645 cell_1rw
* cell instance $1183 r0 *1 108.57,5.46
X$1183 374 5 375 644 645 cell_1rw
* cell instance $1184 r0 *1 109.275,5.46
X$1184 376 5 377 644 645 cell_1rw
* cell instance $1185 r0 *1 109.98,5.46
X$1185 378 5 379 644 645 cell_1rw
* cell instance $1186 r0 *1 110.685,5.46
X$1186 380 5 381 644 645 cell_1rw
* cell instance $1187 r0 *1 111.39,5.46
X$1187 382 5 383 644 645 cell_1rw
* cell instance $1188 r0 *1 112.095,5.46
X$1188 384 5 385 644 645 cell_1rw
* cell instance $1189 r0 *1 112.8,5.46
X$1189 386 5 387 644 645 cell_1rw
* cell instance $1190 r0 *1 113.505,5.46
X$1190 388 5 389 644 645 cell_1rw
* cell instance $1191 r0 *1 114.21,5.46
X$1191 390 5 391 644 645 cell_1rw
* cell instance $1192 r0 *1 114.915,5.46
X$1192 392 5 393 644 645 cell_1rw
* cell instance $1193 r0 *1 115.62,5.46
X$1193 394 5 395 644 645 cell_1rw
* cell instance $1194 r0 *1 116.325,5.46
X$1194 396 5 397 644 645 cell_1rw
* cell instance $1195 r0 *1 117.03,5.46
X$1195 398 5 399 644 645 cell_1rw
* cell instance $1196 r0 *1 117.735,5.46
X$1196 400 5 401 644 645 cell_1rw
* cell instance $1197 r0 *1 118.44,5.46
X$1197 402 5 403 644 645 cell_1rw
* cell instance $1198 r0 *1 119.145,5.46
X$1198 404 5 405 644 645 cell_1rw
* cell instance $1199 r0 *1 119.85,5.46
X$1199 406 5 407 644 645 cell_1rw
* cell instance $1200 r0 *1 120.555,5.46
X$1200 408 5 409 644 645 cell_1rw
* cell instance $1201 r0 *1 121.26,5.46
X$1201 410 5 411 644 645 cell_1rw
* cell instance $1202 r0 *1 121.965,5.46
X$1202 412 5 413 644 645 cell_1rw
* cell instance $1203 r0 *1 122.67,5.46
X$1203 414 5 415 644 645 cell_1rw
* cell instance $1204 r0 *1 123.375,5.46
X$1204 416 5 417 644 645 cell_1rw
* cell instance $1205 r0 *1 124.08,5.46
X$1205 418 5 419 644 645 cell_1rw
* cell instance $1206 r0 *1 124.785,5.46
X$1206 420 5 421 644 645 cell_1rw
* cell instance $1207 r0 *1 125.49,5.46
X$1207 422 5 423 644 645 cell_1rw
* cell instance $1208 r0 *1 126.195,5.46
X$1208 424 5 425 644 645 cell_1rw
* cell instance $1209 r0 *1 126.9,5.46
X$1209 426 5 427 644 645 cell_1rw
* cell instance $1210 r0 *1 127.605,5.46
X$1210 428 5 429 644 645 cell_1rw
* cell instance $1211 r0 *1 128.31,5.46
X$1211 430 5 431 644 645 cell_1rw
* cell instance $1212 r0 *1 129.015,5.46
X$1212 432 5 433 644 645 cell_1rw
* cell instance $1213 r0 *1 129.72,5.46
X$1213 434 5 435 644 645 cell_1rw
* cell instance $1214 r0 *1 130.425,5.46
X$1214 436 5 437 644 645 cell_1rw
* cell instance $1215 r0 *1 131.13,5.46
X$1215 438 5 439 644 645 cell_1rw
* cell instance $1216 r0 *1 131.835,5.46
X$1216 440 5 441 644 645 cell_1rw
* cell instance $1217 r0 *1 132.54,5.46
X$1217 442 5 443 644 645 cell_1rw
* cell instance $1218 r0 *1 133.245,5.46
X$1218 444 5 445 644 645 cell_1rw
* cell instance $1219 r0 *1 133.95,5.46
X$1219 446 5 447 644 645 cell_1rw
* cell instance $1220 r0 *1 134.655,5.46
X$1220 448 5 449 644 645 cell_1rw
* cell instance $1221 r0 *1 135.36,5.46
X$1221 450 5 451 644 645 cell_1rw
* cell instance $1222 r0 *1 136.065,5.46
X$1222 452 5 453 644 645 cell_1rw
* cell instance $1223 r0 *1 136.77,5.46
X$1223 454 5 455 644 645 cell_1rw
* cell instance $1224 r0 *1 137.475,5.46
X$1224 456 5 457 644 645 cell_1rw
* cell instance $1225 r0 *1 138.18,5.46
X$1225 458 5 459 644 645 cell_1rw
* cell instance $1226 r0 *1 138.885,5.46
X$1226 460 5 461 644 645 cell_1rw
* cell instance $1227 r0 *1 139.59,5.46
X$1227 462 5 463 644 645 cell_1rw
* cell instance $1228 r0 *1 140.295,5.46
X$1228 464 5 465 644 645 cell_1rw
* cell instance $1229 r0 *1 141,5.46
X$1229 466 5 467 644 645 cell_1rw
* cell instance $1230 r0 *1 141.705,5.46
X$1230 468 5 469 644 645 cell_1rw
* cell instance $1231 r0 *1 142.41,5.46
X$1231 470 5 471 644 645 cell_1rw
* cell instance $1232 r0 *1 143.115,5.46
X$1232 472 5 473 644 645 cell_1rw
* cell instance $1233 r0 *1 143.82,5.46
X$1233 474 5 475 644 645 cell_1rw
* cell instance $1234 r0 *1 144.525,5.46
X$1234 476 5 477 644 645 cell_1rw
* cell instance $1235 r0 *1 145.23,5.46
X$1235 478 5 479 644 645 cell_1rw
* cell instance $1236 r0 *1 145.935,5.46
X$1236 480 5 481 644 645 cell_1rw
* cell instance $1237 r0 *1 146.64,5.46
X$1237 482 5 483 644 645 cell_1rw
* cell instance $1238 r0 *1 147.345,5.46
X$1238 484 5 485 644 645 cell_1rw
* cell instance $1239 r0 *1 148.05,5.46
X$1239 486 5 487 644 645 cell_1rw
* cell instance $1240 r0 *1 148.755,5.46
X$1240 488 5 489 644 645 cell_1rw
* cell instance $1241 r0 *1 149.46,5.46
X$1241 490 5 491 644 645 cell_1rw
* cell instance $1242 r0 *1 150.165,5.46
X$1242 492 5 493 644 645 cell_1rw
* cell instance $1243 r0 *1 150.87,5.46
X$1243 494 5 495 644 645 cell_1rw
* cell instance $1244 r0 *1 151.575,5.46
X$1244 496 5 497 644 645 cell_1rw
* cell instance $1245 r0 *1 152.28,5.46
X$1245 498 5 499 644 645 cell_1rw
* cell instance $1246 r0 *1 152.985,5.46
X$1246 500 5 501 644 645 cell_1rw
* cell instance $1247 r0 *1 153.69,5.46
X$1247 502 5 503 644 645 cell_1rw
* cell instance $1248 r0 *1 154.395,5.46
X$1248 504 5 505 644 645 cell_1rw
* cell instance $1249 r0 *1 155.1,5.46
X$1249 506 5 507 644 645 cell_1rw
* cell instance $1250 r0 *1 155.805,5.46
X$1250 508 5 509 644 645 cell_1rw
* cell instance $1251 r0 *1 156.51,5.46
X$1251 510 5 511 644 645 cell_1rw
* cell instance $1252 r0 *1 157.215,5.46
X$1252 512 5 513 644 645 cell_1rw
* cell instance $1253 r0 *1 157.92,5.46
X$1253 514 5 515 644 645 cell_1rw
* cell instance $1254 r0 *1 158.625,5.46
X$1254 516 5 517 644 645 cell_1rw
* cell instance $1255 r0 *1 159.33,5.46
X$1255 518 5 519 644 645 cell_1rw
* cell instance $1256 r0 *1 160.035,5.46
X$1256 520 5 521 644 645 cell_1rw
* cell instance $1257 r0 *1 160.74,5.46
X$1257 522 5 523 644 645 cell_1rw
* cell instance $1258 r0 *1 161.445,5.46
X$1258 524 5 525 644 645 cell_1rw
* cell instance $1259 r0 *1 162.15,5.46
X$1259 526 5 527 644 645 cell_1rw
* cell instance $1260 r0 *1 162.855,5.46
X$1260 528 5 529 644 645 cell_1rw
* cell instance $1261 r0 *1 163.56,5.46
X$1261 530 5 531 644 645 cell_1rw
* cell instance $1262 r0 *1 164.265,5.46
X$1262 532 5 533 644 645 cell_1rw
* cell instance $1263 r0 *1 164.97,5.46
X$1263 534 5 535 644 645 cell_1rw
* cell instance $1264 r0 *1 165.675,5.46
X$1264 536 5 537 644 645 cell_1rw
* cell instance $1265 r0 *1 166.38,5.46
X$1265 538 5 539 644 645 cell_1rw
* cell instance $1266 r0 *1 167.085,5.46
X$1266 540 5 541 644 645 cell_1rw
* cell instance $1267 r0 *1 167.79,5.46
X$1267 542 5 543 644 645 cell_1rw
* cell instance $1268 r0 *1 168.495,5.46
X$1268 544 5 545 644 645 cell_1rw
* cell instance $1269 r0 *1 169.2,5.46
X$1269 546 5 547 644 645 cell_1rw
* cell instance $1270 r0 *1 169.905,5.46
X$1270 548 5 549 644 645 cell_1rw
* cell instance $1271 r0 *1 170.61,5.46
X$1271 550 5 551 644 645 cell_1rw
* cell instance $1272 r0 *1 171.315,5.46
X$1272 552 5 553 644 645 cell_1rw
* cell instance $1273 r0 *1 172.02,5.46
X$1273 554 5 555 644 645 cell_1rw
* cell instance $1274 r0 *1 172.725,5.46
X$1274 556 5 557 644 645 cell_1rw
* cell instance $1275 r0 *1 173.43,5.46
X$1275 558 5 559 644 645 cell_1rw
* cell instance $1276 r0 *1 174.135,5.46
X$1276 560 5 561 644 645 cell_1rw
* cell instance $1277 r0 *1 174.84,5.46
X$1277 562 5 563 644 645 cell_1rw
* cell instance $1278 r0 *1 175.545,5.46
X$1278 564 5 565 644 645 cell_1rw
* cell instance $1279 r0 *1 176.25,5.46
X$1279 566 5 567 644 645 cell_1rw
* cell instance $1280 r0 *1 176.955,5.46
X$1280 568 5 569 644 645 cell_1rw
* cell instance $1281 r0 *1 177.66,5.46
X$1281 570 5 571 644 645 cell_1rw
* cell instance $1282 r0 *1 178.365,5.46
X$1282 572 5 573 644 645 cell_1rw
* cell instance $1283 r0 *1 179.07,5.46
X$1283 574 5 575 644 645 cell_1rw
* cell instance $1284 r0 *1 179.775,5.46
X$1284 576 5 577 644 645 cell_1rw
* cell instance $1285 r0 *1 180.48,5.46
X$1285 578 5 579 644 645 cell_1rw
* cell instance $1286 m0 *1 0.705,8.19
X$1286 67 6 68 644 645 cell_1rw
* cell instance $1287 m0 *1 0,8.19
X$1287 65 6 66 644 645 cell_1rw
* cell instance $1288 m0 *1 1.41,8.19
X$1288 69 6 70 644 645 cell_1rw
* cell instance $1289 m0 *1 2.115,8.19
X$1289 71 6 72 644 645 cell_1rw
* cell instance $1290 m0 *1 2.82,8.19
X$1290 73 6 74 644 645 cell_1rw
* cell instance $1291 m0 *1 3.525,8.19
X$1291 75 6 76 644 645 cell_1rw
* cell instance $1292 m0 *1 4.23,8.19
X$1292 77 6 78 644 645 cell_1rw
* cell instance $1293 m0 *1 4.935,8.19
X$1293 79 6 80 644 645 cell_1rw
* cell instance $1294 m0 *1 5.64,8.19
X$1294 81 6 82 644 645 cell_1rw
* cell instance $1295 m0 *1 6.345,8.19
X$1295 83 6 84 644 645 cell_1rw
* cell instance $1296 m0 *1 7.05,8.19
X$1296 85 6 86 644 645 cell_1rw
* cell instance $1297 m0 *1 7.755,8.19
X$1297 87 6 88 644 645 cell_1rw
* cell instance $1298 m0 *1 8.46,8.19
X$1298 89 6 90 644 645 cell_1rw
* cell instance $1299 m0 *1 9.165,8.19
X$1299 91 6 92 644 645 cell_1rw
* cell instance $1300 m0 *1 9.87,8.19
X$1300 93 6 94 644 645 cell_1rw
* cell instance $1301 m0 *1 10.575,8.19
X$1301 95 6 96 644 645 cell_1rw
* cell instance $1302 m0 *1 11.28,8.19
X$1302 97 6 98 644 645 cell_1rw
* cell instance $1303 m0 *1 11.985,8.19
X$1303 99 6 100 644 645 cell_1rw
* cell instance $1304 m0 *1 12.69,8.19
X$1304 101 6 102 644 645 cell_1rw
* cell instance $1305 m0 *1 13.395,8.19
X$1305 103 6 104 644 645 cell_1rw
* cell instance $1306 m0 *1 14.1,8.19
X$1306 105 6 106 644 645 cell_1rw
* cell instance $1307 m0 *1 14.805,8.19
X$1307 107 6 108 644 645 cell_1rw
* cell instance $1308 m0 *1 15.51,8.19
X$1308 109 6 110 644 645 cell_1rw
* cell instance $1309 m0 *1 16.215,8.19
X$1309 111 6 112 644 645 cell_1rw
* cell instance $1310 m0 *1 16.92,8.19
X$1310 113 6 114 644 645 cell_1rw
* cell instance $1311 m0 *1 17.625,8.19
X$1311 115 6 116 644 645 cell_1rw
* cell instance $1312 m0 *1 18.33,8.19
X$1312 117 6 118 644 645 cell_1rw
* cell instance $1313 m0 *1 19.035,8.19
X$1313 119 6 120 644 645 cell_1rw
* cell instance $1314 m0 *1 19.74,8.19
X$1314 121 6 122 644 645 cell_1rw
* cell instance $1315 m0 *1 20.445,8.19
X$1315 123 6 124 644 645 cell_1rw
* cell instance $1316 m0 *1 21.15,8.19
X$1316 125 6 126 644 645 cell_1rw
* cell instance $1317 m0 *1 21.855,8.19
X$1317 127 6 128 644 645 cell_1rw
* cell instance $1318 m0 *1 22.56,8.19
X$1318 129 6 130 644 645 cell_1rw
* cell instance $1319 m0 *1 23.265,8.19
X$1319 131 6 132 644 645 cell_1rw
* cell instance $1320 m0 *1 23.97,8.19
X$1320 133 6 134 644 645 cell_1rw
* cell instance $1321 m0 *1 24.675,8.19
X$1321 135 6 136 644 645 cell_1rw
* cell instance $1322 m0 *1 25.38,8.19
X$1322 137 6 138 644 645 cell_1rw
* cell instance $1323 m0 *1 26.085,8.19
X$1323 139 6 140 644 645 cell_1rw
* cell instance $1324 m0 *1 26.79,8.19
X$1324 141 6 142 644 645 cell_1rw
* cell instance $1325 m0 *1 27.495,8.19
X$1325 143 6 144 644 645 cell_1rw
* cell instance $1326 m0 *1 28.2,8.19
X$1326 145 6 146 644 645 cell_1rw
* cell instance $1327 m0 *1 28.905,8.19
X$1327 147 6 148 644 645 cell_1rw
* cell instance $1328 m0 *1 29.61,8.19
X$1328 149 6 150 644 645 cell_1rw
* cell instance $1329 m0 *1 30.315,8.19
X$1329 151 6 152 644 645 cell_1rw
* cell instance $1330 m0 *1 31.02,8.19
X$1330 153 6 154 644 645 cell_1rw
* cell instance $1331 m0 *1 31.725,8.19
X$1331 155 6 156 644 645 cell_1rw
* cell instance $1332 m0 *1 32.43,8.19
X$1332 157 6 158 644 645 cell_1rw
* cell instance $1333 m0 *1 33.135,8.19
X$1333 159 6 160 644 645 cell_1rw
* cell instance $1334 m0 *1 33.84,8.19
X$1334 161 6 162 644 645 cell_1rw
* cell instance $1335 m0 *1 34.545,8.19
X$1335 163 6 164 644 645 cell_1rw
* cell instance $1336 m0 *1 35.25,8.19
X$1336 165 6 166 644 645 cell_1rw
* cell instance $1337 m0 *1 35.955,8.19
X$1337 167 6 168 644 645 cell_1rw
* cell instance $1338 m0 *1 36.66,8.19
X$1338 169 6 170 644 645 cell_1rw
* cell instance $1339 m0 *1 37.365,8.19
X$1339 171 6 172 644 645 cell_1rw
* cell instance $1340 m0 *1 38.07,8.19
X$1340 173 6 174 644 645 cell_1rw
* cell instance $1341 m0 *1 38.775,8.19
X$1341 175 6 176 644 645 cell_1rw
* cell instance $1342 m0 *1 39.48,8.19
X$1342 177 6 178 644 645 cell_1rw
* cell instance $1343 m0 *1 40.185,8.19
X$1343 179 6 180 644 645 cell_1rw
* cell instance $1344 m0 *1 40.89,8.19
X$1344 181 6 182 644 645 cell_1rw
* cell instance $1345 m0 *1 41.595,8.19
X$1345 183 6 184 644 645 cell_1rw
* cell instance $1346 m0 *1 42.3,8.19
X$1346 185 6 186 644 645 cell_1rw
* cell instance $1347 m0 *1 43.005,8.19
X$1347 187 6 188 644 645 cell_1rw
* cell instance $1348 m0 *1 43.71,8.19
X$1348 189 6 190 644 645 cell_1rw
* cell instance $1349 m0 *1 44.415,8.19
X$1349 191 6 192 644 645 cell_1rw
* cell instance $1350 m0 *1 45.12,8.19
X$1350 193 6 194 644 645 cell_1rw
* cell instance $1351 m0 *1 45.825,8.19
X$1351 195 6 196 644 645 cell_1rw
* cell instance $1352 m0 *1 46.53,8.19
X$1352 197 6 198 644 645 cell_1rw
* cell instance $1353 m0 *1 47.235,8.19
X$1353 199 6 200 644 645 cell_1rw
* cell instance $1354 m0 *1 47.94,8.19
X$1354 201 6 202 644 645 cell_1rw
* cell instance $1355 m0 *1 48.645,8.19
X$1355 203 6 204 644 645 cell_1rw
* cell instance $1356 m0 *1 49.35,8.19
X$1356 205 6 206 644 645 cell_1rw
* cell instance $1357 m0 *1 50.055,8.19
X$1357 207 6 208 644 645 cell_1rw
* cell instance $1358 m0 *1 50.76,8.19
X$1358 209 6 210 644 645 cell_1rw
* cell instance $1359 m0 *1 51.465,8.19
X$1359 211 6 212 644 645 cell_1rw
* cell instance $1360 m0 *1 52.17,8.19
X$1360 213 6 214 644 645 cell_1rw
* cell instance $1361 m0 *1 52.875,8.19
X$1361 215 6 216 644 645 cell_1rw
* cell instance $1362 m0 *1 53.58,8.19
X$1362 217 6 218 644 645 cell_1rw
* cell instance $1363 m0 *1 54.285,8.19
X$1363 219 6 220 644 645 cell_1rw
* cell instance $1364 m0 *1 54.99,8.19
X$1364 221 6 222 644 645 cell_1rw
* cell instance $1365 m0 *1 55.695,8.19
X$1365 223 6 224 644 645 cell_1rw
* cell instance $1366 m0 *1 56.4,8.19
X$1366 225 6 226 644 645 cell_1rw
* cell instance $1367 m0 *1 57.105,8.19
X$1367 227 6 228 644 645 cell_1rw
* cell instance $1368 m0 *1 57.81,8.19
X$1368 229 6 230 644 645 cell_1rw
* cell instance $1369 m0 *1 58.515,8.19
X$1369 231 6 232 644 645 cell_1rw
* cell instance $1370 m0 *1 59.22,8.19
X$1370 233 6 234 644 645 cell_1rw
* cell instance $1371 m0 *1 59.925,8.19
X$1371 235 6 236 644 645 cell_1rw
* cell instance $1372 m0 *1 60.63,8.19
X$1372 237 6 238 644 645 cell_1rw
* cell instance $1373 m0 *1 61.335,8.19
X$1373 239 6 240 644 645 cell_1rw
* cell instance $1374 m0 *1 62.04,8.19
X$1374 241 6 242 644 645 cell_1rw
* cell instance $1375 m0 *1 62.745,8.19
X$1375 243 6 244 644 645 cell_1rw
* cell instance $1376 m0 *1 63.45,8.19
X$1376 245 6 246 644 645 cell_1rw
* cell instance $1377 m0 *1 64.155,8.19
X$1377 247 6 248 644 645 cell_1rw
* cell instance $1378 m0 *1 64.86,8.19
X$1378 249 6 250 644 645 cell_1rw
* cell instance $1379 m0 *1 65.565,8.19
X$1379 251 6 252 644 645 cell_1rw
* cell instance $1380 m0 *1 66.27,8.19
X$1380 253 6 254 644 645 cell_1rw
* cell instance $1381 m0 *1 66.975,8.19
X$1381 255 6 256 644 645 cell_1rw
* cell instance $1382 m0 *1 67.68,8.19
X$1382 257 6 258 644 645 cell_1rw
* cell instance $1383 m0 *1 68.385,8.19
X$1383 259 6 260 644 645 cell_1rw
* cell instance $1384 m0 *1 69.09,8.19
X$1384 261 6 262 644 645 cell_1rw
* cell instance $1385 m0 *1 69.795,8.19
X$1385 263 6 264 644 645 cell_1rw
* cell instance $1386 m0 *1 70.5,8.19
X$1386 265 6 266 644 645 cell_1rw
* cell instance $1387 m0 *1 71.205,8.19
X$1387 267 6 268 644 645 cell_1rw
* cell instance $1388 m0 *1 71.91,8.19
X$1388 269 6 270 644 645 cell_1rw
* cell instance $1389 m0 *1 72.615,8.19
X$1389 271 6 272 644 645 cell_1rw
* cell instance $1390 m0 *1 73.32,8.19
X$1390 273 6 274 644 645 cell_1rw
* cell instance $1391 m0 *1 74.025,8.19
X$1391 275 6 276 644 645 cell_1rw
* cell instance $1392 m0 *1 74.73,8.19
X$1392 277 6 278 644 645 cell_1rw
* cell instance $1393 m0 *1 75.435,8.19
X$1393 279 6 280 644 645 cell_1rw
* cell instance $1394 m0 *1 76.14,8.19
X$1394 281 6 282 644 645 cell_1rw
* cell instance $1395 m0 *1 76.845,8.19
X$1395 283 6 284 644 645 cell_1rw
* cell instance $1396 m0 *1 77.55,8.19
X$1396 285 6 286 644 645 cell_1rw
* cell instance $1397 m0 *1 78.255,8.19
X$1397 287 6 288 644 645 cell_1rw
* cell instance $1398 m0 *1 78.96,8.19
X$1398 289 6 290 644 645 cell_1rw
* cell instance $1399 m0 *1 79.665,8.19
X$1399 291 6 292 644 645 cell_1rw
* cell instance $1400 m0 *1 80.37,8.19
X$1400 293 6 294 644 645 cell_1rw
* cell instance $1401 m0 *1 81.075,8.19
X$1401 295 6 296 644 645 cell_1rw
* cell instance $1402 m0 *1 81.78,8.19
X$1402 297 6 298 644 645 cell_1rw
* cell instance $1403 m0 *1 82.485,8.19
X$1403 299 6 300 644 645 cell_1rw
* cell instance $1404 m0 *1 83.19,8.19
X$1404 301 6 302 644 645 cell_1rw
* cell instance $1405 m0 *1 83.895,8.19
X$1405 303 6 304 644 645 cell_1rw
* cell instance $1406 m0 *1 84.6,8.19
X$1406 305 6 306 644 645 cell_1rw
* cell instance $1407 m0 *1 85.305,8.19
X$1407 307 6 308 644 645 cell_1rw
* cell instance $1408 m0 *1 86.01,8.19
X$1408 309 6 310 644 645 cell_1rw
* cell instance $1409 m0 *1 86.715,8.19
X$1409 311 6 312 644 645 cell_1rw
* cell instance $1410 m0 *1 87.42,8.19
X$1410 313 6 314 644 645 cell_1rw
* cell instance $1411 m0 *1 88.125,8.19
X$1411 315 6 316 644 645 cell_1rw
* cell instance $1412 m0 *1 88.83,8.19
X$1412 317 6 318 644 645 cell_1rw
* cell instance $1413 m0 *1 89.535,8.19
X$1413 319 6 320 644 645 cell_1rw
* cell instance $1414 m0 *1 90.24,8.19
X$1414 321 6 323 644 645 cell_1rw
* cell instance $1415 m0 *1 90.945,8.19
X$1415 324 6 325 644 645 cell_1rw
* cell instance $1416 m0 *1 91.65,8.19
X$1416 326 6 327 644 645 cell_1rw
* cell instance $1417 m0 *1 92.355,8.19
X$1417 328 6 329 644 645 cell_1rw
* cell instance $1418 m0 *1 93.06,8.19
X$1418 330 6 331 644 645 cell_1rw
* cell instance $1419 m0 *1 93.765,8.19
X$1419 332 6 333 644 645 cell_1rw
* cell instance $1420 m0 *1 94.47,8.19
X$1420 334 6 335 644 645 cell_1rw
* cell instance $1421 m0 *1 95.175,8.19
X$1421 336 6 337 644 645 cell_1rw
* cell instance $1422 m0 *1 95.88,8.19
X$1422 338 6 339 644 645 cell_1rw
* cell instance $1423 m0 *1 96.585,8.19
X$1423 340 6 341 644 645 cell_1rw
* cell instance $1424 m0 *1 97.29,8.19
X$1424 342 6 343 644 645 cell_1rw
* cell instance $1425 m0 *1 97.995,8.19
X$1425 344 6 345 644 645 cell_1rw
* cell instance $1426 m0 *1 98.7,8.19
X$1426 346 6 347 644 645 cell_1rw
* cell instance $1427 m0 *1 99.405,8.19
X$1427 348 6 349 644 645 cell_1rw
* cell instance $1428 m0 *1 100.11,8.19
X$1428 350 6 351 644 645 cell_1rw
* cell instance $1429 m0 *1 100.815,8.19
X$1429 352 6 353 644 645 cell_1rw
* cell instance $1430 m0 *1 101.52,8.19
X$1430 354 6 355 644 645 cell_1rw
* cell instance $1431 m0 *1 102.225,8.19
X$1431 356 6 357 644 645 cell_1rw
* cell instance $1432 m0 *1 102.93,8.19
X$1432 358 6 359 644 645 cell_1rw
* cell instance $1433 m0 *1 103.635,8.19
X$1433 360 6 361 644 645 cell_1rw
* cell instance $1434 m0 *1 104.34,8.19
X$1434 362 6 363 644 645 cell_1rw
* cell instance $1435 m0 *1 105.045,8.19
X$1435 364 6 365 644 645 cell_1rw
* cell instance $1436 m0 *1 105.75,8.19
X$1436 366 6 367 644 645 cell_1rw
* cell instance $1437 m0 *1 106.455,8.19
X$1437 368 6 369 644 645 cell_1rw
* cell instance $1438 m0 *1 107.16,8.19
X$1438 370 6 371 644 645 cell_1rw
* cell instance $1439 m0 *1 107.865,8.19
X$1439 372 6 373 644 645 cell_1rw
* cell instance $1440 m0 *1 108.57,8.19
X$1440 374 6 375 644 645 cell_1rw
* cell instance $1441 m0 *1 109.275,8.19
X$1441 376 6 377 644 645 cell_1rw
* cell instance $1442 m0 *1 109.98,8.19
X$1442 378 6 379 644 645 cell_1rw
* cell instance $1443 m0 *1 110.685,8.19
X$1443 380 6 381 644 645 cell_1rw
* cell instance $1444 m0 *1 111.39,8.19
X$1444 382 6 383 644 645 cell_1rw
* cell instance $1445 m0 *1 112.095,8.19
X$1445 384 6 385 644 645 cell_1rw
* cell instance $1446 m0 *1 112.8,8.19
X$1446 386 6 387 644 645 cell_1rw
* cell instance $1447 m0 *1 113.505,8.19
X$1447 388 6 389 644 645 cell_1rw
* cell instance $1448 m0 *1 114.21,8.19
X$1448 390 6 391 644 645 cell_1rw
* cell instance $1449 m0 *1 114.915,8.19
X$1449 392 6 393 644 645 cell_1rw
* cell instance $1450 m0 *1 115.62,8.19
X$1450 394 6 395 644 645 cell_1rw
* cell instance $1451 m0 *1 116.325,8.19
X$1451 396 6 397 644 645 cell_1rw
* cell instance $1452 m0 *1 117.03,8.19
X$1452 398 6 399 644 645 cell_1rw
* cell instance $1453 m0 *1 117.735,8.19
X$1453 400 6 401 644 645 cell_1rw
* cell instance $1454 m0 *1 118.44,8.19
X$1454 402 6 403 644 645 cell_1rw
* cell instance $1455 m0 *1 119.145,8.19
X$1455 404 6 405 644 645 cell_1rw
* cell instance $1456 m0 *1 119.85,8.19
X$1456 406 6 407 644 645 cell_1rw
* cell instance $1457 m0 *1 120.555,8.19
X$1457 408 6 409 644 645 cell_1rw
* cell instance $1458 m0 *1 121.26,8.19
X$1458 410 6 411 644 645 cell_1rw
* cell instance $1459 m0 *1 121.965,8.19
X$1459 412 6 413 644 645 cell_1rw
* cell instance $1460 m0 *1 122.67,8.19
X$1460 414 6 415 644 645 cell_1rw
* cell instance $1461 m0 *1 123.375,8.19
X$1461 416 6 417 644 645 cell_1rw
* cell instance $1462 m0 *1 124.08,8.19
X$1462 418 6 419 644 645 cell_1rw
* cell instance $1463 m0 *1 124.785,8.19
X$1463 420 6 421 644 645 cell_1rw
* cell instance $1464 m0 *1 125.49,8.19
X$1464 422 6 423 644 645 cell_1rw
* cell instance $1465 m0 *1 126.195,8.19
X$1465 424 6 425 644 645 cell_1rw
* cell instance $1466 m0 *1 126.9,8.19
X$1466 426 6 427 644 645 cell_1rw
* cell instance $1467 m0 *1 127.605,8.19
X$1467 428 6 429 644 645 cell_1rw
* cell instance $1468 m0 *1 128.31,8.19
X$1468 430 6 431 644 645 cell_1rw
* cell instance $1469 m0 *1 129.015,8.19
X$1469 432 6 433 644 645 cell_1rw
* cell instance $1470 m0 *1 129.72,8.19
X$1470 434 6 435 644 645 cell_1rw
* cell instance $1471 m0 *1 130.425,8.19
X$1471 436 6 437 644 645 cell_1rw
* cell instance $1472 m0 *1 131.13,8.19
X$1472 438 6 439 644 645 cell_1rw
* cell instance $1473 m0 *1 131.835,8.19
X$1473 440 6 441 644 645 cell_1rw
* cell instance $1474 m0 *1 132.54,8.19
X$1474 442 6 443 644 645 cell_1rw
* cell instance $1475 m0 *1 133.245,8.19
X$1475 444 6 445 644 645 cell_1rw
* cell instance $1476 m0 *1 133.95,8.19
X$1476 446 6 447 644 645 cell_1rw
* cell instance $1477 m0 *1 134.655,8.19
X$1477 448 6 449 644 645 cell_1rw
* cell instance $1478 m0 *1 135.36,8.19
X$1478 450 6 451 644 645 cell_1rw
* cell instance $1479 m0 *1 136.065,8.19
X$1479 452 6 453 644 645 cell_1rw
* cell instance $1480 m0 *1 136.77,8.19
X$1480 454 6 455 644 645 cell_1rw
* cell instance $1481 m0 *1 137.475,8.19
X$1481 456 6 457 644 645 cell_1rw
* cell instance $1482 m0 *1 138.18,8.19
X$1482 458 6 459 644 645 cell_1rw
* cell instance $1483 m0 *1 138.885,8.19
X$1483 460 6 461 644 645 cell_1rw
* cell instance $1484 m0 *1 139.59,8.19
X$1484 462 6 463 644 645 cell_1rw
* cell instance $1485 m0 *1 140.295,8.19
X$1485 464 6 465 644 645 cell_1rw
* cell instance $1486 m0 *1 141,8.19
X$1486 466 6 467 644 645 cell_1rw
* cell instance $1487 m0 *1 141.705,8.19
X$1487 468 6 469 644 645 cell_1rw
* cell instance $1488 m0 *1 142.41,8.19
X$1488 470 6 471 644 645 cell_1rw
* cell instance $1489 m0 *1 143.115,8.19
X$1489 472 6 473 644 645 cell_1rw
* cell instance $1490 m0 *1 143.82,8.19
X$1490 474 6 475 644 645 cell_1rw
* cell instance $1491 m0 *1 144.525,8.19
X$1491 476 6 477 644 645 cell_1rw
* cell instance $1492 m0 *1 145.23,8.19
X$1492 478 6 479 644 645 cell_1rw
* cell instance $1493 m0 *1 145.935,8.19
X$1493 480 6 481 644 645 cell_1rw
* cell instance $1494 m0 *1 146.64,8.19
X$1494 482 6 483 644 645 cell_1rw
* cell instance $1495 m0 *1 147.345,8.19
X$1495 484 6 485 644 645 cell_1rw
* cell instance $1496 m0 *1 148.05,8.19
X$1496 486 6 487 644 645 cell_1rw
* cell instance $1497 m0 *1 148.755,8.19
X$1497 488 6 489 644 645 cell_1rw
* cell instance $1498 m0 *1 149.46,8.19
X$1498 490 6 491 644 645 cell_1rw
* cell instance $1499 m0 *1 150.165,8.19
X$1499 492 6 493 644 645 cell_1rw
* cell instance $1500 m0 *1 150.87,8.19
X$1500 494 6 495 644 645 cell_1rw
* cell instance $1501 m0 *1 151.575,8.19
X$1501 496 6 497 644 645 cell_1rw
* cell instance $1502 m0 *1 152.28,8.19
X$1502 498 6 499 644 645 cell_1rw
* cell instance $1503 m0 *1 152.985,8.19
X$1503 500 6 501 644 645 cell_1rw
* cell instance $1504 m0 *1 153.69,8.19
X$1504 502 6 503 644 645 cell_1rw
* cell instance $1505 m0 *1 154.395,8.19
X$1505 504 6 505 644 645 cell_1rw
* cell instance $1506 m0 *1 155.1,8.19
X$1506 506 6 507 644 645 cell_1rw
* cell instance $1507 m0 *1 155.805,8.19
X$1507 508 6 509 644 645 cell_1rw
* cell instance $1508 m0 *1 156.51,8.19
X$1508 510 6 511 644 645 cell_1rw
* cell instance $1509 m0 *1 157.215,8.19
X$1509 512 6 513 644 645 cell_1rw
* cell instance $1510 m0 *1 157.92,8.19
X$1510 514 6 515 644 645 cell_1rw
* cell instance $1511 m0 *1 158.625,8.19
X$1511 516 6 517 644 645 cell_1rw
* cell instance $1512 m0 *1 159.33,8.19
X$1512 518 6 519 644 645 cell_1rw
* cell instance $1513 m0 *1 160.035,8.19
X$1513 520 6 521 644 645 cell_1rw
* cell instance $1514 m0 *1 160.74,8.19
X$1514 522 6 523 644 645 cell_1rw
* cell instance $1515 m0 *1 161.445,8.19
X$1515 524 6 525 644 645 cell_1rw
* cell instance $1516 m0 *1 162.15,8.19
X$1516 526 6 527 644 645 cell_1rw
* cell instance $1517 m0 *1 162.855,8.19
X$1517 528 6 529 644 645 cell_1rw
* cell instance $1518 m0 *1 163.56,8.19
X$1518 530 6 531 644 645 cell_1rw
* cell instance $1519 m0 *1 164.265,8.19
X$1519 532 6 533 644 645 cell_1rw
* cell instance $1520 m0 *1 164.97,8.19
X$1520 534 6 535 644 645 cell_1rw
* cell instance $1521 m0 *1 165.675,8.19
X$1521 536 6 537 644 645 cell_1rw
* cell instance $1522 m0 *1 166.38,8.19
X$1522 538 6 539 644 645 cell_1rw
* cell instance $1523 m0 *1 167.085,8.19
X$1523 540 6 541 644 645 cell_1rw
* cell instance $1524 m0 *1 167.79,8.19
X$1524 542 6 543 644 645 cell_1rw
* cell instance $1525 m0 *1 168.495,8.19
X$1525 544 6 545 644 645 cell_1rw
* cell instance $1526 m0 *1 169.2,8.19
X$1526 546 6 547 644 645 cell_1rw
* cell instance $1527 m0 *1 169.905,8.19
X$1527 548 6 549 644 645 cell_1rw
* cell instance $1528 m0 *1 170.61,8.19
X$1528 550 6 551 644 645 cell_1rw
* cell instance $1529 m0 *1 171.315,8.19
X$1529 552 6 553 644 645 cell_1rw
* cell instance $1530 m0 *1 172.02,8.19
X$1530 554 6 555 644 645 cell_1rw
* cell instance $1531 m0 *1 172.725,8.19
X$1531 556 6 557 644 645 cell_1rw
* cell instance $1532 m0 *1 173.43,8.19
X$1532 558 6 559 644 645 cell_1rw
* cell instance $1533 m0 *1 174.135,8.19
X$1533 560 6 561 644 645 cell_1rw
* cell instance $1534 m0 *1 174.84,8.19
X$1534 562 6 563 644 645 cell_1rw
* cell instance $1535 m0 *1 175.545,8.19
X$1535 564 6 565 644 645 cell_1rw
* cell instance $1536 m0 *1 176.25,8.19
X$1536 566 6 567 644 645 cell_1rw
* cell instance $1537 m0 *1 176.955,8.19
X$1537 568 6 569 644 645 cell_1rw
* cell instance $1538 m0 *1 177.66,8.19
X$1538 570 6 571 644 645 cell_1rw
* cell instance $1539 m0 *1 178.365,8.19
X$1539 572 6 573 644 645 cell_1rw
* cell instance $1540 m0 *1 179.07,8.19
X$1540 574 6 575 644 645 cell_1rw
* cell instance $1541 m0 *1 179.775,8.19
X$1541 576 6 577 644 645 cell_1rw
* cell instance $1542 m0 *1 180.48,8.19
X$1542 578 6 579 644 645 cell_1rw
* cell instance $1543 r0 *1 0.705,8.19
X$1543 67 7 68 644 645 cell_1rw
* cell instance $1544 r0 *1 0,8.19
X$1544 65 7 66 644 645 cell_1rw
* cell instance $1545 r0 *1 1.41,8.19
X$1545 69 7 70 644 645 cell_1rw
* cell instance $1546 r0 *1 2.115,8.19
X$1546 71 7 72 644 645 cell_1rw
* cell instance $1547 r0 *1 2.82,8.19
X$1547 73 7 74 644 645 cell_1rw
* cell instance $1548 r0 *1 3.525,8.19
X$1548 75 7 76 644 645 cell_1rw
* cell instance $1549 r0 *1 4.23,8.19
X$1549 77 7 78 644 645 cell_1rw
* cell instance $1550 r0 *1 4.935,8.19
X$1550 79 7 80 644 645 cell_1rw
* cell instance $1551 r0 *1 5.64,8.19
X$1551 81 7 82 644 645 cell_1rw
* cell instance $1552 r0 *1 6.345,8.19
X$1552 83 7 84 644 645 cell_1rw
* cell instance $1553 r0 *1 7.05,8.19
X$1553 85 7 86 644 645 cell_1rw
* cell instance $1554 r0 *1 7.755,8.19
X$1554 87 7 88 644 645 cell_1rw
* cell instance $1555 r0 *1 8.46,8.19
X$1555 89 7 90 644 645 cell_1rw
* cell instance $1556 r0 *1 9.165,8.19
X$1556 91 7 92 644 645 cell_1rw
* cell instance $1557 r0 *1 9.87,8.19
X$1557 93 7 94 644 645 cell_1rw
* cell instance $1558 r0 *1 10.575,8.19
X$1558 95 7 96 644 645 cell_1rw
* cell instance $1559 r0 *1 11.28,8.19
X$1559 97 7 98 644 645 cell_1rw
* cell instance $1560 r0 *1 11.985,8.19
X$1560 99 7 100 644 645 cell_1rw
* cell instance $1561 r0 *1 12.69,8.19
X$1561 101 7 102 644 645 cell_1rw
* cell instance $1562 r0 *1 13.395,8.19
X$1562 103 7 104 644 645 cell_1rw
* cell instance $1563 r0 *1 14.1,8.19
X$1563 105 7 106 644 645 cell_1rw
* cell instance $1564 r0 *1 14.805,8.19
X$1564 107 7 108 644 645 cell_1rw
* cell instance $1565 r0 *1 15.51,8.19
X$1565 109 7 110 644 645 cell_1rw
* cell instance $1566 r0 *1 16.215,8.19
X$1566 111 7 112 644 645 cell_1rw
* cell instance $1567 r0 *1 16.92,8.19
X$1567 113 7 114 644 645 cell_1rw
* cell instance $1568 r0 *1 17.625,8.19
X$1568 115 7 116 644 645 cell_1rw
* cell instance $1569 r0 *1 18.33,8.19
X$1569 117 7 118 644 645 cell_1rw
* cell instance $1570 r0 *1 19.035,8.19
X$1570 119 7 120 644 645 cell_1rw
* cell instance $1571 r0 *1 19.74,8.19
X$1571 121 7 122 644 645 cell_1rw
* cell instance $1572 r0 *1 20.445,8.19
X$1572 123 7 124 644 645 cell_1rw
* cell instance $1573 r0 *1 21.15,8.19
X$1573 125 7 126 644 645 cell_1rw
* cell instance $1574 r0 *1 21.855,8.19
X$1574 127 7 128 644 645 cell_1rw
* cell instance $1575 r0 *1 22.56,8.19
X$1575 129 7 130 644 645 cell_1rw
* cell instance $1576 r0 *1 23.265,8.19
X$1576 131 7 132 644 645 cell_1rw
* cell instance $1577 r0 *1 23.97,8.19
X$1577 133 7 134 644 645 cell_1rw
* cell instance $1578 r0 *1 24.675,8.19
X$1578 135 7 136 644 645 cell_1rw
* cell instance $1579 r0 *1 25.38,8.19
X$1579 137 7 138 644 645 cell_1rw
* cell instance $1580 r0 *1 26.085,8.19
X$1580 139 7 140 644 645 cell_1rw
* cell instance $1581 r0 *1 26.79,8.19
X$1581 141 7 142 644 645 cell_1rw
* cell instance $1582 r0 *1 27.495,8.19
X$1582 143 7 144 644 645 cell_1rw
* cell instance $1583 r0 *1 28.2,8.19
X$1583 145 7 146 644 645 cell_1rw
* cell instance $1584 r0 *1 28.905,8.19
X$1584 147 7 148 644 645 cell_1rw
* cell instance $1585 r0 *1 29.61,8.19
X$1585 149 7 150 644 645 cell_1rw
* cell instance $1586 r0 *1 30.315,8.19
X$1586 151 7 152 644 645 cell_1rw
* cell instance $1587 r0 *1 31.02,8.19
X$1587 153 7 154 644 645 cell_1rw
* cell instance $1588 r0 *1 31.725,8.19
X$1588 155 7 156 644 645 cell_1rw
* cell instance $1589 r0 *1 32.43,8.19
X$1589 157 7 158 644 645 cell_1rw
* cell instance $1590 r0 *1 33.135,8.19
X$1590 159 7 160 644 645 cell_1rw
* cell instance $1591 r0 *1 33.84,8.19
X$1591 161 7 162 644 645 cell_1rw
* cell instance $1592 r0 *1 34.545,8.19
X$1592 163 7 164 644 645 cell_1rw
* cell instance $1593 r0 *1 35.25,8.19
X$1593 165 7 166 644 645 cell_1rw
* cell instance $1594 r0 *1 35.955,8.19
X$1594 167 7 168 644 645 cell_1rw
* cell instance $1595 r0 *1 36.66,8.19
X$1595 169 7 170 644 645 cell_1rw
* cell instance $1596 r0 *1 37.365,8.19
X$1596 171 7 172 644 645 cell_1rw
* cell instance $1597 r0 *1 38.07,8.19
X$1597 173 7 174 644 645 cell_1rw
* cell instance $1598 r0 *1 38.775,8.19
X$1598 175 7 176 644 645 cell_1rw
* cell instance $1599 r0 *1 39.48,8.19
X$1599 177 7 178 644 645 cell_1rw
* cell instance $1600 r0 *1 40.185,8.19
X$1600 179 7 180 644 645 cell_1rw
* cell instance $1601 r0 *1 40.89,8.19
X$1601 181 7 182 644 645 cell_1rw
* cell instance $1602 r0 *1 41.595,8.19
X$1602 183 7 184 644 645 cell_1rw
* cell instance $1603 r0 *1 42.3,8.19
X$1603 185 7 186 644 645 cell_1rw
* cell instance $1604 r0 *1 43.005,8.19
X$1604 187 7 188 644 645 cell_1rw
* cell instance $1605 r0 *1 43.71,8.19
X$1605 189 7 190 644 645 cell_1rw
* cell instance $1606 r0 *1 44.415,8.19
X$1606 191 7 192 644 645 cell_1rw
* cell instance $1607 r0 *1 45.12,8.19
X$1607 193 7 194 644 645 cell_1rw
* cell instance $1608 r0 *1 45.825,8.19
X$1608 195 7 196 644 645 cell_1rw
* cell instance $1609 r0 *1 46.53,8.19
X$1609 197 7 198 644 645 cell_1rw
* cell instance $1610 r0 *1 47.235,8.19
X$1610 199 7 200 644 645 cell_1rw
* cell instance $1611 r0 *1 47.94,8.19
X$1611 201 7 202 644 645 cell_1rw
* cell instance $1612 r0 *1 48.645,8.19
X$1612 203 7 204 644 645 cell_1rw
* cell instance $1613 r0 *1 49.35,8.19
X$1613 205 7 206 644 645 cell_1rw
* cell instance $1614 r0 *1 50.055,8.19
X$1614 207 7 208 644 645 cell_1rw
* cell instance $1615 r0 *1 50.76,8.19
X$1615 209 7 210 644 645 cell_1rw
* cell instance $1616 r0 *1 51.465,8.19
X$1616 211 7 212 644 645 cell_1rw
* cell instance $1617 r0 *1 52.17,8.19
X$1617 213 7 214 644 645 cell_1rw
* cell instance $1618 r0 *1 52.875,8.19
X$1618 215 7 216 644 645 cell_1rw
* cell instance $1619 r0 *1 53.58,8.19
X$1619 217 7 218 644 645 cell_1rw
* cell instance $1620 r0 *1 54.285,8.19
X$1620 219 7 220 644 645 cell_1rw
* cell instance $1621 r0 *1 54.99,8.19
X$1621 221 7 222 644 645 cell_1rw
* cell instance $1622 r0 *1 55.695,8.19
X$1622 223 7 224 644 645 cell_1rw
* cell instance $1623 r0 *1 56.4,8.19
X$1623 225 7 226 644 645 cell_1rw
* cell instance $1624 r0 *1 57.105,8.19
X$1624 227 7 228 644 645 cell_1rw
* cell instance $1625 r0 *1 57.81,8.19
X$1625 229 7 230 644 645 cell_1rw
* cell instance $1626 r0 *1 58.515,8.19
X$1626 231 7 232 644 645 cell_1rw
* cell instance $1627 r0 *1 59.22,8.19
X$1627 233 7 234 644 645 cell_1rw
* cell instance $1628 r0 *1 59.925,8.19
X$1628 235 7 236 644 645 cell_1rw
* cell instance $1629 r0 *1 60.63,8.19
X$1629 237 7 238 644 645 cell_1rw
* cell instance $1630 r0 *1 61.335,8.19
X$1630 239 7 240 644 645 cell_1rw
* cell instance $1631 r0 *1 62.04,8.19
X$1631 241 7 242 644 645 cell_1rw
* cell instance $1632 r0 *1 62.745,8.19
X$1632 243 7 244 644 645 cell_1rw
* cell instance $1633 r0 *1 63.45,8.19
X$1633 245 7 246 644 645 cell_1rw
* cell instance $1634 r0 *1 64.155,8.19
X$1634 247 7 248 644 645 cell_1rw
* cell instance $1635 r0 *1 64.86,8.19
X$1635 249 7 250 644 645 cell_1rw
* cell instance $1636 r0 *1 65.565,8.19
X$1636 251 7 252 644 645 cell_1rw
* cell instance $1637 r0 *1 66.27,8.19
X$1637 253 7 254 644 645 cell_1rw
* cell instance $1638 r0 *1 66.975,8.19
X$1638 255 7 256 644 645 cell_1rw
* cell instance $1639 r0 *1 67.68,8.19
X$1639 257 7 258 644 645 cell_1rw
* cell instance $1640 r0 *1 68.385,8.19
X$1640 259 7 260 644 645 cell_1rw
* cell instance $1641 r0 *1 69.09,8.19
X$1641 261 7 262 644 645 cell_1rw
* cell instance $1642 r0 *1 69.795,8.19
X$1642 263 7 264 644 645 cell_1rw
* cell instance $1643 r0 *1 70.5,8.19
X$1643 265 7 266 644 645 cell_1rw
* cell instance $1644 r0 *1 71.205,8.19
X$1644 267 7 268 644 645 cell_1rw
* cell instance $1645 r0 *1 71.91,8.19
X$1645 269 7 270 644 645 cell_1rw
* cell instance $1646 r0 *1 72.615,8.19
X$1646 271 7 272 644 645 cell_1rw
* cell instance $1647 r0 *1 73.32,8.19
X$1647 273 7 274 644 645 cell_1rw
* cell instance $1648 r0 *1 74.025,8.19
X$1648 275 7 276 644 645 cell_1rw
* cell instance $1649 r0 *1 74.73,8.19
X$1649 277 7 278 644 645 cell_1rw
* cell instance $1650 r0 *1 75.435,8.19
X$1650 279 7 280 644 645 cell_1rw
* cell instance $1651 r0 *1 76.14,8.19
X$1651 281 7 282 644 645 cell_1rw
* cell instance $1652 r0 *1 76.845,8.19
X$1652 283 7 284 644 645 cell_1rw
* cell instance $1653 r0 *1 77.55,8.19
X$1653 285 7 286 644 645 cell_1rw
* cell instance $1654 r0 *1 78.255,8.19
X$1654 287 7 288 644 645 cell_1rw
* cell instance $1655 r0 *1 78.96,8.19
X$1655 289 7 290 644 645 cell_1rw
* cell instance $1656 r0 *1 79.665,8.19
X$1656 291 7 292 644 645 cell_1rw
* cell instance $1657 r0 *1 80.37,8.19
X$1657 293 7 294 644 645 cell_1rw
* cell instance $1658 r0 *1 81.075,8.19
X$1658 295 7 296 644 645 cell_1rw
* cell instance $1659 r0 *1 81.78,8.19
X$1659 297 7 298 644 645 cell_1rw
* cell instance $1660 r0 *1 82.485,8.19
X$1660 299 7 300 644 645 cell_1rw
* cell instance $1661 r0 *1 83.19,8.19
X$1661 301 7 302 644 645 cell_1rw
* cell instance $1662 r0 *1 83.895,8.19
X$1662 303 7 304 644 645 cell_1rw
* cell instance $1663 r0 *1 84.6,8.19
X$1663 305 7 306 644 645 cell_1rw
* cell instance $1664 r0 *1 85.305,8.19
X$1664 307 7 308 644 645 cell_1rw
* cell instance $1665 r0 *1 86.01,8.19
X$1665 309 7 310 644 645 cell_1rw
* cell instance $1666 r0 *1 86.715,8.19
X$1666 311 7 312 644 645 cell_1rw
* cell instance $1667 r0 *1 87.42,8.19
X$1667 313 7 314 644 645 cell_1rw
* cell instance $1668 r0 *1 88.125,8.19
X$1668 315 7 316 644 645 cell_1rw
* cell instance $1669 r0 *1 88.83,8.19
X$1669 317 7 318 644 645 cell_1rw
* cell instance $1670 r0 *1 89.535,8.19
X$1670 319 7 320 644 645 cell_1rw
* cell instance $1671 r0 *1 90.24,8.19
X$1671 321 7 323 644 645 cell_1rw
* cell instance $1672 r0 *1 90.945,8.19
X$1672 324 7 325 644 645 cell_1rw
* cell instance $1673 r0 *1 91.65,8.19
X$1673 326 7 327 644 645 cell_1rw
* cell instance $1674 r0 *1 92.355,8.19
X$1674 328 7 329 644 645 cell_1rw
* cell instance $1675 r0 *1 93.06,8.19
X$1675 330 7 331 644 645 cell_1rw
* cell instance $1676 r0 *1 93.765,8.19
X$1676 332 7 333 644 645 cell_1rw
* cell instance $1677 r0 *1 94.47,8.19
X$1677 334 7 335 644 645 cell_1rw
* cell instance $1678 r0 *1 95.175,8.19
X$1678 336 7 337 644 645 cell_1rw
* cell instance $1679 r0 *1 95.88,8.19
X$1679 338 7 339 644 645 cell_1rw
* cell instance $1680 r0 *1 96.585,8.19
X$1680 340 7 341 644 645 cell_1rw
* cell instance $1681 r0 *1 97.29,8.19
X$1681 342 7 343 644 645 cell_1rw
* cell instance $1682 r0 *1 97.995,8.19
X$1682 344 7 345 644 645 cell_1rw
* cell instance $1683 r0 *1 98.7,8.19
X$1683 346 7 347 644 645 cell_1rw
* cell instance $1684 r0 *1 99.405,8.19
X$1684 348 7 349 644 645 cell_1rw
* cell instance $1685 r0 *1 100.11,8.19
X$1685 350 7 351 644 645 cell_1rw
* cell instance $1686 r0 *1 100.815,8.19
X$1686 352 7 353 644 645 cell_1rw
* cell instance $1687 r0 *1 101.52,8.19
X$1687 354 7 355 644 645 cell_1rw
* cell instance $1688 r0 *1 102.225,8.19
X$1688 356 7 357 644 645 cell_1rw
* cell instance $1689 r0 *1 102.93,8.19
X$1689 358 7 359 644 645 cell_1rw
* cell instance $1690 r0 *1 103.635,8.19
X$1690 360 7 361 644 645 cell_1rw
* cell instance $1691 r0 *1 104.34,8.19
X$1691 362 7 363 644 645 cell_1rw
* cell instance $1692 r0 *1 105.045,8.19
X$1692 364 7 365 644 645 cell_1rw
* cell instance $1693 r0 *1 105.75,8.19
X$1693 366 7 367 644 645 cell_1rw
* cell instance $1694 r0 *1 106.455,8.19
X$1694 368 7 369 644 645 cell_1rw
* cell instance $1695 r0 *1 107.16,8.19
X$1695 370 7 371 644 645 cell_1rw
* cell instance $1696 r0 *1 107.865,8.19
X$1696 372 7 373 644 645 cell_1rw
* cell instance $1697 r0 *1 108.57,8.19
X$1697 374 7 375 644 645 cell_1rw
* cell instance $1698 r0 *1 109.275,8.19
X$1698 376 7 377 644 645 cell_1rw
* cell instance $1699 r0 *1 109.98,8.19
X$1699 378 7 379 644 645 cell_1rw
* cell instance $1700 r0 *1 110.685,8.19
X$1700 380 7 381 644 645 cell_1rw
* cell instance $1701 r0 *1 111.39,8.19
X$1701 382 7 383 644 645 cell_1rw
* cell instance $1702 r0 *1 112.095,8.19
X$1702 384 7 385 644 645 cell_1rw
* cell instance $1703 r0 *1 112.8,8.19
X$1703 386 7 387 644 645 cell_1rw
* cell instance $1704 r0 *1 113.505,8.19
X$1704 388 7 389 644 645 cell_1rw
* cell instance $1705 r0 *1 114.21,8.19
X$1705 390 7 391 644 645 cell_1rw
* cell instance $1706 r0 *1 114.915,8.19
X$1706 392 7 393 644 645 cell_1rw
* cell instance $1707 r0 *1 115.62,8.19
X$1707 394 7 395 644 645 cell_1rw
* cell instance $1708 r0 *1 116.325,8.19
X$1708 396 7 397 644 645 cell_1rw
* cell instance $1709 r0 *1 117.03,8.19
X$1709 398 7 399 644 645 cell_1rw
* cell instance $1710 r0 *1 117.735,8.19
X$1710 400 7 401 644 645 cell_1rw
* cell instance $1711 r0 *1 118.44,8.19
X$1711 402 7 403 644 645 cell_1rw
* cell instance $1712 r0 *1 119.145,8.19
X$1712 404 7 405 644 645 cell_1rw
* cell instance $1713 r0 *1 119.85,8.19
X$1713 406 7 407 644 645 cell_1rw
* cell instance $1714 r0 *1 120.555,8.19
X$1714 408 7 409 644 645 cell_1rw
* cell instance $1715 r0 *1 121.26,8.19
X$1715 410 7 411 644 645 cell_1rw
* cell instance $1716 r0 *1 121.965,8.19
X$1716 412 7 413 644 645 cell_1rw
* cell instance $1717 r0 *1 122.67,8.19
X$1717 414 7 415 644 645 cell_1rw
* cell instance $1718 r0 *1 123.375,8.19
X$1718 416 7 417 644 645 cell_1rw
* cell instance $1719 r0 *1 124.08,8.19
X$1719 418 7 419 644 645 cell_1rw
* cell instance $1720 r0 *1 124.785,8.19
X$1720 420 7 421 644 645 cell_1rw
* cell instance $1721 r0 *1 125.49,8.19
X$1721 422 7 423 644 645 cell_1rw
* cell instance $1722 r0 *1 126.195,8.19
X$1722 424 7 425 644 645 cell_1rw
* cell instance $1723 r0 *1 126.9,8.19
X$1723 426 7 427 644 645 cell_1rw
* cell instance $1724 r0 *1 127.605,8.19
X$1724 428 7 429 644 645 cell_1rw
* cell instance $1725 r0 *1 128.31,8.19
X$1725 430 7 431 644 645 cell_1rw
* cell instance $1726 r0 *1 129.015,8.19
X$1726 432 7 433 644 645 cell_1rw
* cell instance $1727 r0 *1 129.72,8.19
X$1727 434 7 435 644 645 cell_1rw
* cell instance $1728 r0 *1 130.425,8.19
X$1728 436 7 437 644 645 cell_1rw
* cell instance $1729 r0 *1 131.13,8.19
X$1729 438 7 439 644 645 cell_1rw
* cell instance $1730 r0 *1 131.835,8.19
X$1730 440 7 441 644 645 cell_1rw
* cell instance $1731 r0 *1 132.54,8.19
X$1731 442 7 443 644 645 cell_1rw
* cell instance $1732 r0 *1 133.245,8.19
X$1732 444 7 445 644 645 cell_1rw
* cell instance $1733 r0 *1 133.95,8.19
X$1733 446 7 447 644 645 cell_1rw
* cell instance $1734 r0 *1 134.655,8.19
X$1734 448 7 449 644 645 cell_1rw
* cell instance $1735 r0 *1 135.36,8.19
X$1735 450 7 451 644 645 cell_1rw
* cell instance $1736 r0 *1 136.065,8.19
X$1736 452 7 453 644 645 cell_1rw
* cell instance $1737 r0 *1 136.77,8.19
X$1737 454 7 455 644 645 cell_1rw
* cell instance $1738 r0 *1 137.475,8.19
X$1738 456 7 457 644 645 cell_1rw
* cell instance $1739 r0 *1 138.18,8.19
X$1739 458 7 459 644 645 cell_1rw
* cell instance $1740 r0 *1 138.885,8.19
X$1740 460 7 461 644 645 cell_1rw
* cell instance $1741 r0 *1 139.59,8.19
X$1741 462 7 463 644 645 cell_1rw
* cell instance $1742 r0 *1 140.295,8.19
X$1742 464 7 465 644 645 cell_1rw
* cell instance $1743 r0 *1 141,8.19
X$1743 466 7 467 644 645 cell_1rw
* cell instance $1744 r0 *1 141.705,8.19
X$1744 468 7 469 644 645 cell_1rw
* cell instance $1745 r0 *1 142.41,8.19
X$1745 470 7 471 644 645 cell_1rw
* cell instance $1746 r0 *1 143.115,8.19
X$1746 472 7 473 644 645 cell_1rw
* cell instance $1747 r0 *1 143.82,8.19
X$1747 474 7 475 644 645 cell_1rw
* cell instance $1748 r0 *1 144.525,8.19
X$1748 476 7 477 644 645 cell_1rw
* cell instance $1749 r0 *1 145.23,8.19
X$1749 478 7 479 644 645 cell_1rw
* cell instance $1750 r0 *1 145.935,8.19
X$1750 480 7 481 644 645 cell_1rw
* cell instance $1751 r0 *1 146.64,8.19
X$1751 482 7 483 644 645 cell_1rw
* cell instance $1752 r0 *1 147.345,8.19
X$1752 484 7 485 644 645 cell_1rw
* cell instance $1753 r0 *1 148.05,8.19
X$1753 486 7 487 644 645 cell_1rw
* cell instance $1754 r0 *1 148.755,8.19
X$1754 488 7 489 644 645 cell_1rw
* cell instance $1755 r0 *1 149.46,8.19
X$1755 490 7 491 644 645 cell_1rw
* cell instance $1756 r0 *1 150.165,8.19
X$1756 492 7 493 644 645 cell_1rw
* cell instance $1757 r0 *1 150.87,8.19
X$1757 494 7 495 644 645 cell_1rw
* cell instance $1758 r0 *1 151.575,8.19
X$1758 496 7 497 644 645 cell_1rw
* cell instance $1759 r0 *1 152.28,8.19
X$1759 498 7 499 644 645 cell_1rw
* cell instance $1760 r0 *1 152.985,8.19
X$1760 500 7 501 644 645 cell_1rw
* cell instance $1761 r0 *1 153.69,8.19
X$1761 502 7 503 644 645 cell_1rw
* cell instance $1762 r0 *1 154.395,8.19
X$1762 504 7 505 644 645 cell_1rw
* cell instance $1763 r0 *1 155.1,8.19
X$1763 506 7 507 644 645 cell_1rw
* cell instance $1764 r0 *1 155.805,8.19
X$1764 508 7 509 644 645 cell_1rw
* cell instance $1765 r0 *1 156.51,8.19
X$1765 510 7 511 644 645 cell_1rw
* cell instance $1766 r0 *1 157.215,8.19
X$1766 512 7 513 644 645 cell_1rw
* cell instance $1767 r0 *1 157.92,8.19
X$1767 514 7 515 644 645 cell_1rw
* cell instance $1768 r0 *1 158.625,8.19
X$1768 516 7 517 644 645 cell_1rw
* cell instance $1769 r0 *1 159.33,8.19
X$1769 518 7 519 644 645 cell_1rw
* cell instance $1770 r0 *1 160.035,8.19
X$1770 520 7 521 644 645 cell_1rw
* cell instance $1771 r0 *1 160.74,8.19
X$1771 522 7 523 644 645 cell_1rw
* cell instance $1772 r0 *1 161.445,8.19
X$1772 524 7 525 644 645 cell_1rw
* cell instance $1773 r0 *1 162.15,8.19
X$1773 526 7 527 644 645 cell_1rw
* cell instance $1774 r0 *1 162.855,8.19
X$1774 528 7 529 644 645 cell_1rw
* cell instance $1775 r0 *1 163.56,8.19
X$1775 530 7 531 644 645 cell_1rw
* cell instance $1776 r0 *1 164.265,8.19
X$1776 532 7 533 644 645 cell_1rw
* cell instance $1777 r0 *1 164.97,8.19
X$1777 534 7 535 644 645 cell_1rw
* cell instance $1778 r0 *1 165.675,8.19
X$1778 536 7 537 644 645 cell_1rw
* cell instance $1779 r0 *1 166.38,8.19
X$1779 538 7 539 644 645 cell_1rw
* cell instance $1780 r0 *1 167.085,8.19
X$1780 540 7 541 644 645 cell_1rw
* cell instance $1781 r0 *1 167.79,8.19
X$1781 542 7 543 644 645 cell_1rw
* cell instance $1782 r0 *1 168.495,8.19
X$1782 544 7 545 644 645 cell_1rw
* cell instance $1783 r0 *1 169.2,8.19
X$1783 546 7 547 644 645 cell_1rw
* cell instance $1784 r0 *1 169.905,8.19
X$1784 548 7 549 644 645 cell_1rw
* cell instance $1785 r0 *1 170.61,8.19
X$1785 550 7 551 644 645 cell_1rw
* cell instance $1786 r0 *1 171.315,8.19
X$1786 552 7 553 644 645 cell_1rw
* cell instance $1787 r0 *1 172.02,8.19
X$1787 554 7 555 644 645 cell_1rw
* cell instance $1788 r0 *1 172.725,8.19
X$1788 556 7 557 644 645 cell_1rw
* cell instance $1789 r0 *1 173.43,8.19
X$1789 558 7 559 644 645 cell_1rw
* cell instance $1790 r0 *1 174.135,8.19
X$1790 560 7 561 644 645 cell_1rw
* cell instance $1791 r0 *1 174.84,8.19
X$1791 562 7 563 644 645 cell_1rw
* cell instance $1792 r0 *1 175.545,8.19
X$1792 564 7 565 644 645 cell_1rw
* cell instance $1793 r0 *1 176.25,8.19
X$1793 566 7 567 644 645 cell_1rw
* cell instance $1794 r0 *1 176.955,8.19
X$1794 568 7 569 644 645 cell_1rw
* cell instance $1795 r0 *1 177.66,8.19
X$1795 570 7 571 644 645 cell_1rw
* cell instance $1796 r0 *1 178.365,8.19
X$1796 572 7 573 644 645 cell_1rw
* cell instance $1797 r0 *1 179.07,8.19
X$1797 574 7 575 644 645 cell_1rw
* cell instance $1798 r0 *1 179.775,8.19
X$1798 576 7 577 644 645 cell_1rw
* cell instance $1799 r0 *1 180.48,8.19
X$1799 578 7 579 644 645 cell_1rw
* cell instance $1800 m0 *1 0.705,10.92
X$1800 67 8 68 644 645 cell_1rw
* cell instance $1801 m0 *1 0,10.92
X$1801 65 8 66 644 645 cell_1rw
* cell instance $1802 m0 *1 1.41,10.92
X$1802 69 8 70 644 645 cell_1rw
* cell instance $1803 m0 *1 2.115,10.92
X$1803 71 8 72 644 645 cell_1rw
* cell instance $1804 m0 *1 2.82,10.92
X$1804 73 8 74 644 645 cell_1rw
* cell instance $1805 m0 *1 3.525,10.92
X$1805 75 8 76 644 645 cell_1rw
* cell instance $1806 m0 *1 4.23,10.92
X$1806 77 8 78 644 645 cell_1rw
* cell instance $1807 m0 *1 4.935,10.92
X$1807 79 8 80 644 645 cell_1rw
* cell instance $1808 m0 *1 5.64,10.92
X$1808 81 8 82 644 645 cell_1rw
* cell instance $1809 m0 *1 6.345,10.92
X$1809 83 8 84 644 645 cell_1rw
* cell instance $1810 m0 *1 7.05,10.92
X$1810 85 8 86 644 645 cell_1rw
* cell instance $1811 m0 *1 7.755,10.92
X$1811 87 8 88 644 645 cell_1rw
* cell instance $1812 m0 *1 8.46,10.92
X$1812 89 8 90 644 645 cell_1rw
* cell instance $1813 m0 *1 9.165,10.92
X$1813 91 8 92 644 645 cell_1rw
* cell instance $1814 m0 *1 9.87,10.92
X$1814 93 8 94 644 645 cell_1rw
* cell instance $1815 m0 *1 10.575,10.92
X$1815 95 8 96 644 645 cell_1rw
* cell instance $1816 m0 *1 11.28,10.92
X$1816 97 8 98 644 645 cell_1rw
* cell instance $1817 m0 *1 11.985,10.92
X$1817 99 8 100 644 645 cell_1rw
* cell instance $1818 m0 *1 12.69,10.92
X$1818 101 8 102 644 645 cell_1rw
* cell instance $1819 m0 *1 13.395,10.92
X$1819 103 8 104 644 645 cell_1rw
* cell instance $1820 m0 *1 14.1,10.92
X$1820 105 8 106 644 645 cell_1rw
* cell instance $1821 m0 *1 14.805,10.92
X$1821 107 8 108 644 645 cell_1rw
* cell instance $1822 m0 *1 15.51,10.92
X$1822 109 8 110 644 645 cell_1rw
* cell instance $1823 m0 *1 16.215,10.92
X$1823 111 8 112 644 645 cell_1rw
* cell instance $1824 m0 *1 16.92,10.92
X$1824 113 8 114 644 645 cell_1rw
* cell instance $1825 m0 *1 17.625,10.92
X$1825 115 8 116 644 645 cell_1rw
* cell instance $1826 m0 *1 18.33,10.92
X$1826 117 8 118 644 645 cell_1rw
* cell instance $1827 m0 *1 19.035,10.92
X$1827 119 8 120 644 645 cell_1rw
* cell instance $1828 m0 *1 19.74,10.92
X$1828 121 8 122 644 645 cell_1rw
* cell instance $1829 m0 *1 20.445,10.92
X$1829 123 8 124 644 645 cell_1rw
* cell instance $1830 m0 *1 21.15,10.92
X$1830 125 8 126 644 645 cell_1rw
* cell instance $1831 m0 *1 21.855,10.92
X$1831 127 8 128 644 645 cell_1rw
* cell instance $1832 m0 *1 22.56,10.92
X$1832 129 8 130 644 645 cell_1rw
* cell instance $1833 m0 *1 23.265,10.92
X$1833 131 8 132 644 645 cell_1rw
* cell instance $1834 m0 *1 23.97,10.92
X$1834 133 8 134 644 645 cell_1rw
* cell instance $1835 m0 *1 24.675,10.92
X$1835 135 8 136 644 645 cell_1rw
* cell instance $1836 m0 *1 25.38,10.92
X$1836 137 8 138 644 645 cell_1rw
* cell instance $1837 m0 *1 26.085,10.92
X$1837 139 8 140 644 645 cell_1rw
* cell instance $1838 m0 *1 26.79,10.92
X$1838 141 8 142 644 645 cell_1rw
* cell instance $1839 m0 *1 27.495,10.92
X$1839 143 8 144 644 645 cell_1rw
* cell instance $1840 m0 *1 28.2,10.92
X$1840 145 8 146 644 645 cell_1rw
* cell instance $1841 m0 *1 28.905,10.92
X$1841 147 8 148 644 645 cell_1rw
* cell instance $1842 m0 *1 29.61,10.92
X$1842 149 8 150 644 645 cell_1rw
* cell instance $1843 m0 *1 30.315,10.92
X$1843 151 8 152 644 645 cell_1rw
* cell instance $1844 m0 *1 31.02,10.92
X$1844 153 8 154 644 645 cell_1rw
* cell instance $1845 m0 *1 31.725,10.92
X$1845 155 8 156 644 645 cell_1rw
* cell instance $1846 m0 *1 32.43,10.92
X$1846 157 8 158 644 645 cell_1rw
* cell instance $1847 m0 *1 33.135,10.92
X$1847 159 8 160 644 645 cell_1rw
* cell instance $1848 m0 *1 33.84,10.92
X$1848 161 8 162 644 645 cell_1rw
* cell instance $1849 m0 *1 34.545,10.92
X$1849 163 8 164 644 645 cell_1rw
* cell instance $1850 m0 *1 35.25,10.92
X$1850 165 8 166 644 645 cell_1rw
* cell instance $1851 m0 *1 35.955,10.92
X$1851 167 8 168 644 645 cell_1rw
* cell instance $1852 m0 *1 36.66,10.92
X$1852 169 8 170 644 645 cell_1rw
* cell instance $1853 m0 *1 37.365,10.92
X$1853 171 8 172 644 645 cell_1rw
* cell instance $1854 m0 *1 38.07,10.92
X$1854 173 8 174 644 645 cell_1rw
* cell instance $1855 m0 *1 38.775,10.92
X$1855 175 8 176 644 645 cell_1rw
* cell instance $1856 m0 *1 39.48,10.92
X$1856 177 8 178 644 645 cell_1rw
* cell instance $1857 m0 *1 40.185,10.92
X$1857 179 8 180 644 645 cell_1rw
* cell instance $1858 m0 *1 40.89,10.92
X$1858 181 8 182 644 645 cell_1rw
* cell instance $1859 m0 *1 41.595,10.92
X$1859 183 8 184 644 645 cell_1rw
* cell instance $1860 m0 *1 42.3,10.92
X$1860 185 8 186 644 645 cell_1rw
* cell instance $1861 m0 *1 43.005,10.92
X$1861 187 8 188 644 645 cell_1rw
* cell instance $1862 m0 *1 43.71,10.92
X$1862 189 8 190 644 645 cell_1rw
* cell instance $1863 m0 *1 44.415,10.92
X$1863 191 8 192 644 645 cell_1rw
* cell instance $1864 m0 *1 45.12,10.92
X$1864 193 8 194 644 645 cell_1rw
* cell instance $1865 m0 *1 45.825,10.92
X$1865 195 8 196 644 645 cell_1rw
* cell instance $1866 m0 *1 46.53,10.92
X$1866 197 8 198 644 645 cell_1rw
* cell instance $1867 m0 *1 47.235,10.92
X$1867 199 8 200 644 645 cell_1rw
* cell instance $1868 m0 *1 47.94,10.92
X$1868 201 8 202 644 645 cell_1rw
* cell instance $1869 m0 *1 48.645,10.92
X$1869 203 8 204 644 645 cell_1rw
* cell instance $1870 m0 *1 49.35,10.92
X$1870 205 8 206 644 645 cell_1rw
* cell instance $1871 m0 *1 50.055,10.92
X$1871 207 8 208 644 645 cell_1rw
* cell instance $1872 m0 *1 50.76,10.92
X$1872 209 8 210 644 645 cell_1rw
* cell instance $1873 m0 *1 51.465,10.92
X$1873 211 8 212 644 645 cell_1rw
* cell instance $1874 m0 *1 52.17,10.92
X$1874 213 8 214 644 645 cell_1rw
* cell instance $1875 m0 *1 52.875,10.92
X$1875 215 8 216 644 645 cell_1rw
* cell instance $1876 m0 *1 53.58,10.92
X$1876 217 8 218 644 645 cell_1rw
* cell instance $1877 m0 *1 54.285,10.92
X$1877 219 8 220 644 645 cell_1rw
* cell instance $1878 m0 *1 54.99,10.92
X$1878 221 8 222 644 645 cell_1rw
* cell instance $1879 m0 *1 55.695,10.92
X$1879 223 8 224 644 645 cell_1rw
* cell instance $1880 m0 *1 56.4,10.92
X$1880 225 8 226 644 645 cell_1rw
* cell instance $1881 m0 *1 57.105,10.92
X$1881 227 8 228 644 645 cell_1rw
* cell instance $1882 m0 *1 57.81,10.92
X$1882 229 8 230 644 645 cell_1rw
* cell instance $1883 m0 *1 58.515,10.92
X$1883 231 8 232 644 645 cell_1rw
* cell instance $1884 m0 *1 59.22,10.92
X$1884 233 8 234 644 645 cell_1rw
* cell instance $1885 m0 *1 59.925,10.92
X$1885 235 8 236 644 645 cell_1rw
* cell instance $1886 m0 *1 60.63,10.92
X$1886 237 8 238 644 645 cell_1rw
* cell instance $1887 m0 *1 61.335,10.92
X$1887 239 8 240 644 645 cell_1rw
* cell instance $1888 m0 *1 62.04,10.92
X$1888 241 8 242 644 645 cell_1rw
* cell instance $1889 m0 *1 62.745,10.92
X$1889 243 8 244 644 645 cell_1rw
* cell instance $1890 m0 *1 63.45,10.92
X$1890 245 8 246 644 645 cell_1rw
* cell instance $1891 m0 *1 64.155,10.92
X$1891 247 8 248 644 645 cell_1rw
* cell instance $1892 m0 *1 64.86,10.92
X$1892 249 8 250 644 645 cell_1rw
* cell instance $1893 m0 *1 65.565,10.92
X$1893 251 8 252 644 645 cell_1rw
* cell instance $1894 m0 *1 66.27,10.92
X$1894 253 8 254 644 645 cell_1rw
* cell instance $1895 m0 *1 66.975,10.92
X$1895 255 8 256 644 645 cell_1rw
* cell instance $1896 m0 *1 67.68,10.92
X$1896 257 8 258 644 645 cell_1rw
* cell instance $1897 m0 *1 68.385,10.92
X$1897 259 8 260 644 645 cell_1rw
* cell instance $1898 m0 *1 69.09,10.92
X$1898 261 8 262 644 645 cell_1rw
* cell instance $1899 m0 *1 69.795,10.92
X$1899 263 8 264 644 645 cell_1rw
* cell instance $1900 m0 *1 70.5,10.92
X$1900 265 8 266 644 645 cell_1rw
* cell instance $1901 m0 *1 71.205,10.92
X$1901 267 8 268 644 645 cell_1rw
* cell instance $1902 m0 *1 71.91,10.92
X$1902 269 8 270 644 645 cell_1rw
* cell instance $1903 m0 *1 72.615,10.92
X$1903 271 8 272 644 645 cell_1rw
* cell instance $1904 m0 *1 73.32,10.92
X$1904 273 8 274 644 645 cell_1rw
* cell instance $1905 m0 *1 74.025,10.92
X$1905 275 8 276 644 645 cell_1rw
* cell instance $1906 m0 *1 74.73,10.92
X$1906 277 8 278 644 645 cell_1rw
* cell instance $1907 m0 *1 75.435,10.92
X$1907 279 8 280 644 645 cell_1rw
* cell instance $1908 m0 *1 76.14,10.92
X$1908 281 8 282 644 645 cell_1rw
* cell instance $1909 m0 *1 76.845,10.92
X$1909 283 8 284 644 645 cell_1rw
* cell instance $1910 m0 *1 77.55,10.92
X$1910 285 8 286 644 645 cell_1rw
* cell instance $1911 m0 *1 78.255,10.92
X$1911 287 8 288 644 645 cell_1rw
* cell instance $1912 m0 *1 78.96,10.92
X$1912 289 8 290 644 645 cell_1rw
* cell instance $1913 m0 *1 79.665,10.92
X$1913 291 8 292 644 645 cell_1rw
* cell instance $1914 m0 *1 80.37,10.92
X$1914 293 8 294 644 645 cell_1rw
* cell instance $1915 m0 *1 81.075,10.92
X$1915 295 8 296 644 645 cell_1rw
* cell instance $1916 m0 *1 81.78,10.92
X$1916 297 8 298 644 645 cell_1rw
* cell instance $1917 m0 *1 82.485,10.92
X$1917 299 8 300 644 645 cell_1rw
* cell instance $1918 m0 *1 83.19,10.92
X$1918 301 8 302 644 645 cell_1rw
* cell instance $1919 m0 *1 83.895,10.92
X$1919 303 8 304 644 645 cell_1rw
* cell instance $1920 m0 *1 84.6,10.92
X$1920 305 8 306 644 645 cell_1rw
* cell instance $1921 m0 *1 85.305,10.92
X$1921 307 8 308 644 645 cell_1rw
* cell instance $1922 m0 *1 86.01,10.92
X$1922 309 8 310 644 645 cell_1rw
* cell instance $1923 m0 *1 86.715,10.92
X$1923 311 8 312 644 645 cell_1rw
* cell instance $1924 m0 *1 87.42,10.92
X$1924 313 8 314 644 645 cell_1rw
* cell instance $1925 m0 *1 88.125,10.92
X$1925 315 8 316 644 645 cell_1rw
* cell instance $1926 m0 *1 88.83,10.92
X$1926 317 8 318 644 645 cell_1rw
* cell instance $1927 m0 *1 89.535,10.92
X$1927 319 8 320 644 645 cell_1rw
* cell instance $1928 m0 *1 90.24,10.92
X$1928 321 8 323 644 645 cell_1rw
* cell instance $1929 m0 *1 90.945,10.92
X$1929 324 8 325 644 645 cell_1rw
* cell instance $1930 m0 *1 91.65,10.92
X$1930 326 8 327 644 645 cell_1rw
* cell instance $1931 m0 *1 92.355,10.92
X$1931 328 8 329 644 645 cell_1rw
* cell instance $1932 m0 *1 93.06,10.92
X$1932 330 8 331 644 645 cell_1rw
* cell instance $1933 m0 *1 93.765,10.92
X$1933 332 8 333 644 645 cell_1rw
* cell instance $1934 m0 *1 94.47,10.92
X$1934 334 8 335 644 645 cell_1rw
* cell instance $1935 m0 *1 95.175,10.92
X$1935 336 8 337 644 645 cell_1rw
* cell instance $1936 m0 *1 95.88,10.92
X$1936 338 8 339 644 645 cell_1rw
* cell instance $1937 m0 *1 96.585,10.92
X$1937 340 8 341 644 645 cell_1rw
* cell instance $1938 m0 *1 97.29,10.92
X$1938 342 8 343 644 645 cell_1rw
* cell instance $1939 m0 *1 97.995,10.92
X$1939 344 8 345 644 645 cell_1rw
* cell instance $1940 m0 *1 98.7,10.92
X$1940 346 8 347 644 645 cell_1rw
* cell instance $1941 m0 *1 99.405,10.92
X$1941 348 8 349 644 645 cell_1rw
* cell instance $1942 m0 *1 100.11,10.92
X$1942 350 8 351 644 645 cell_1rw
* cell instance $1943 m0 *1 100.815,10.92
X$1943 352 8 353 644 645 cell_1rw
* cell instance $1944 m0 *1 101.52,10.92
X$1944 354 8 355 644 645 cell_1rw
* cell instance $1945 m0 *1 102.225,10.92
X$1945 356 8 357 644 645 cell_1rw
* cell instance $1946 m0 *1 102.93,10.92
X$1946 358 8 359 644 645 cell_1rw
* cell instance $1947 m0 *1 103.635,10.92
X$1947 360 8 361 644 645 cell_1rw
* cell instance $1948 m0 *1 104.34,10.92
X$1948 362 8 363 644 645 cell_1rw
* cell instance $1949 m0 *1 105.045,10.92
X$1949 364 8 365 644 645 cell_1rw
* cell instance $1950 m0 *1 105.75,10.92
X$1950 366 8 367 644 645 cell_1rw
* cell instance $1951 m0 *1 106.455,10.92
X$1951 368 8 369 644 645 cell_1rw
* cell instance $1952 m0 *1 107.16,10.92
X$1952 370 8 371 644 645 cell_1rw
* cell instance $1953 m0 *1 107.865,10.92
X$1953 372 8 373 644 645 cell_1rw
* cell instance $1954 m0 *1 108.57,10.92
X$1954 374 8 375 644 645 cell_1rw
* cell instance $1955 m0 *1 109.275,10.92
X$1955 376 8 377 644 645 cell_1rw
* cell instance $1956 m0 *1 109.98,10.92
X$1956 378 8 379 644 645 cell_1rw
* cell instance $1957 m0 *1 110.685,10.92
X$1957 380 8 381 644 645 cell_1rw
* cell instance $1958 m0 *1 111.39,10.92
X$1958 382 8 383 644 645 cell_1rw
* cell instance $1959 m0 *1 112.095,10.92
X$1959 384 8 385 644 645 cell_1rw
* cell instance $1960 m0 *1 112.8,10.92
X$1960 386 8 387 644 645 cell_1rw
* cell instance $1961 m0 *1 113.505,10.92
X$1961 388 8 389 644 645 cell_1rw
* cell instance $1962 m0 *1 114.21,10.92
X$1962 390 8 391 644 645 cell_1rw
* cell instance $1963 m0 *1 114.915,10.92
X$1963 392 8 393 644 645 cell_1rw
* cell instance $1964 m0 *1 115.62,10.92
X$1964 394 8 395 644 645 cell_1rw
* cell instance $1965 m0 *1 116.325,10.92
X$1965 396 8 397 644 645 cell_1rw
* cell instance $1966 m0 *1 117.03,10.92
X$1966 398 8 399 644 645 cell_1rw
* cell instance $1967 m0 *1 117.735,10.92
X$1967 400 8 401 644 645 cell_1rw
* cell instance $1968 m0 *1 118.44,10.92
X$1968 402 8 403 644 645 cell_1rw
* cell instance $1969 m0 *1 119.145,10.92
X$1969 404 8 405 644 645 cell_1rw
* cell instance $1970 m0 *1 119.85,10.92
X$1970 406 8 407 644 645 cell_1rw
* cell instance $1971 m0 *1 120.555,10.92
X$1971 408 8 409 644 645 cell_1rw
* cell instance $1972 m0 *1 121.26,10.92
X$1972 410 8 411 644 645 cell_1rw
* cell instance $1973 m0 *1 121.965,10.92
X$1973 412 8 413 644 645 cell_1rw
* cell instance $1974 m0 *1 122.67,10.92
X$1974 414 8 415 644 645 cell_1rw
* cell instance $1975 m0 *1 123.375,10.92
X$1975 416 8 417 644 645 cell_1rw
* cell instance $1976 m0 *1 124.08,10.92
X$1976 418 8 419 644 645 cell_1rw
* cell instance $1977 m0 *1 124.785,10.92
X$1977 420 8 421 644 645 cell_1rw
* cell instance $1978 m0 *1 125.49,10.92
X$1978 422 8 423 644 645 cell_1rw
* cell instance $1979 m0 *1 126.195,10.92
X$1979 424 8 425 644 645 cell_1rw
* cell instance $1980 m0 *1 126.9,10.92
X$1980 426 8 427 644 645 cell_1rw
* cell instance $1981 m0 *1 127.605,10.92
X$1981 428 8 429 644 645 cell_1rw
* cell instance $1982 m0 *1 128.31,10.92
X$1982 430 8 431 644 645 cell_1rw
* cell instance $1983 m0 *1 129.015,10.92
X$1983 432 8 433 644 645 cell_1rw
* cell instance $1984 m0 *1 129.72,10.92
X$1984 434 8 435 644 645 cell_1rw
* cell instance $1985 m0 *1 130.425,10.92
X$1985 436 8 437 644 645 cell_1rw
* cell instance $1986 m0 *1 131.13,10.92
X$1986 438 8 439 644 645 cell_1rw
* cell instance $1987 m0 *1 131.835,10.92
X$1987 440 8 441 644 645 cell_1rw
* cell instance $1988 m0 *1 132.54,10.92
X$1988 442 8 443 644 645 cell_1rw
* cell instance $1989 m0 *1 133.245,10.92
X$1989 444 8 445 644 645 cell_1rw
* cell instance $1990 m0 *1 133.95,10.92
X$1990 446 8 447 644 645 cell_1rw
* cell instance $1991 m0 *1 134.655,10.92
X$1991 448 8 449 644 645 cell_1rw
* cell instance $1992 m0 *1 135.36,10.92
X$1992 450 8 451 644 645 cell_1rw
* cell instance $1993 m0 *1 136.065,10.92
X$1993 452 8 453 644 645 cell_1rw
* cell instance $1994 m0 *1 136.77,10.92
X$1994 454 8 455 644 645 cell_1rw
* cell instance $1995 m0 *1 137.475,10.92
X$1995 456 8 457 644 645 cell_1rw
* cell instance $1996 m0 *1 138.18,10.92
X$1996 458 8 459 644 645 cell_1rw
* cell instance $1997 m0 *1 138.885,10.92
X$1997 460 8 461 644 645 cell_1rw
* cell instance $1998 m0 *1 139.59,10.92
X$1998 462 8 463 644 645 cell_1rw
* cell instance $1999 m0 *1 140.295,10.92
X$1999 464 8 465 644 645 cell_1rw
* cell instance $2000 m0 *1 141,10.92
X$2000 466 8 467 644 645 cell_1rw
* cell instance $2001 m0 *1 141.705,10.92
X$2001 468 8 469 644 645 cell_1rw
* cell instance $2002 m0 *1 142.41,10.92
X$2002 470 8 471 644 645 cell_1rw
* cell instance $2003 m0 *1 143.115,10.92
X$2003 472 8 473 644 645 cell_1rw
* cell instance $2004 m0 *1 143.82,10.92
X$2004 474 8 475 644 645 cell_1rw
* cell instance $2005 m0 *1 144.525,10.92
X$2005 476 8 477 644 645 cell_1rw
* cell instance $2006 m0 *1 145.23,10.92
X$2006 478 8 479 644 645 cell_1rw
* cell instance $2007 m0 *1 145.935,10.92
X$2007 480 8 481 644 645 cell_1rw
* cell instance $2008 m0 *1 146.64,10.92
X$2008 482 8 483 644 645 cell_1rw
* cell instance $2009 m0 *1 147.345,10.92
X$2009 484 8 485 644 645 cell_1rw
* cell instance $2010 m0 *1 148.05,10.92
X$2010 486 8 487 644 645 cell_1rw
* cell instance $2011 m0 *1 148.755,10.92
X$2011 488 8 489 644 645 cell_1rw
* cell instance $2012 m0 *1 149.46,10.92
X$2012 490 8 491 644 645 cell_1rw
* cell instance $2013 m0 *1 150.165,10.92
X$2013 492 8 493 644 645 cell_1rw
* cell instance $2014 m0 *1 150.87,10.92
X$2014 494 8 495 644 645 cell_1rw
* cell instance $2015 m0 *1 151.575,10.92
X$2015 496 8 497 644 645 cell_1rw
* cell instance $2016 m0 *1 152.28,10.92
X$2016 498 8 499 644 645 cell_1rw
* cell instance $2017 m0 *1 152.985,10.92
X$2017 500 8 501 644 645 cell_1rw
* cell instance $2018 m0 *1 153.69,10.92
X$2018 502 8 503 644 645 cell_1rw
* cell instance $2019 m0 *1 154.395,10.92
X$2019 504 8 505 644 645 cell_1rw
* cell instance $2020 m0 *1 155.1,10.92
X$2020 506 8 507 644 645 cell_1rw
* cell instance $2021 m0 *1 155.805,10.92
X$2021 508 8 509 644 645 cell_1rw
* cell instance $2022 m0 *1 156.51,10.92
X$2022 510 8 511 644 645 cell_1rw
* cell instance $2023 m0 *1 157.215,10.92
X$2023 512 8 513 644 645 cell_1rw
* cell instance $2024 m0 *1 157.92,10.92
X$2024 514 8 515 644 645 cell_1rw
* cell instance $2025 m0 *1 158.625,10.92
X$2025 516 8 517 644 645 cell_1rw
* cell instance $2026 m0 *1 159.33,10.92
X$2026 518 8 519 644 645 cell_1rw
* cell instance $2027 m0 *1 160.035,10.92
X$2027 520 8 521 644 645 cell_1rw
* cell instance $2028 m0 *1 160.74,10.92
X$2028 522 8 523 644 645 cell_1rw
* cell instance $2029 m0 *1 161.445,10.92
X$2029 524 8 525 644 645 cell_1rw
* cell instance $2030 m0 *1 162.15,10.92
X$2030 526 8 527 644 645 cell_1rw
* cell instance $2031 m0 *1 162.855,10.92
X$2031 528 8 529 644 645 cell_1rw
* cell instance $2032 m0 *1 163.56,10.92
X$2032 530 8 531 644 645 cell_1rw
* cell instance $2033 m0 *1 164.265,10.92
X$2033 532 8 533 644 645 cell_1rw
* cell instance $2034 m0 *1 164.97,10.92
X$2034 534 8 535 644 645 cell_1rw
* cell instance $2035 m0 *1 165.675,10.92
X$2035 536 8 537 644 645 cell_1rw
* cell instance $2036 m0 *1 166.38,10.92
X$2036 538 8 539 644 645 cell_1rw
* cell instance $2037 m0 *1 167.085,10.92
X$2037 540 8 541 644 645 cell_1rw
* cell instance $2038 m0 *1 167.79,10.92
X$2038 542 8 543 644 645 cell_1rw
* cell instance $2039 m0 *1 168.495,10.92
X$2039 544 8 545 644 645 cell_1rw
* cell instance $2040 m0 *1 169.2,10.92
X$2040 546 8 547 644 645 cell_1rw
* cell instance $2041 m0 *1 169.905,10.92
X$2041 548 8 549 644 645 cell_1rw
* cell instance $2042 m0 *1 170.61,10.92
X$2042 550 8 551 644 645 cell_1rw
* cell instance $2043 m0 *1 171.315,10.92
X$2043 552 8 553 644 645 cell_1rw
* cell instance $2044 m0 *1 172.02,10.92
X$2044 554 8 555 644 645 cell_1rw
* cell instance $2045 m0 *1 172.725,10.92
X$2045 556 8 557 644 645 cell_1rw
* cell instance $2046 m0 *1 173.43,10.92
X$2046 558 8 559 644 645 cell_1rw
* cell instance $2047 m0 *1 174.135,10.92
X$2047 560 8 561 644 645 cell_1rw
* cell instance $2048 m0 *1 174.84,10.92
X$2048 562 8 563 644 645 cell_1rw
* cell instance $2049 m0 *1 175.545,10.92
X$2049 564 8 565 644 645 cell_1rw
* cell instance $2050 m0 *1 176.25,10.92
X$2050 566 8 567 644 645 cell_1rw
* cell instance $2051 m0 *1 176.955,10.92
X$2051 568 8 569 644 645 cell_1rw
* cell instance $2052 m0 *1 177.66,10.92
X$2052 570 8 571 644 645 cell_1rw
* cell instance $2053 m0 *1 178.365,10.92
X$2053 572 8 573 644 645 cell_1rw
* cell instance $2054 m0 *1 179.07,10.92
X$2054 574 8 575 644 645 cell_1rw
* cell instance $2055 m0 *1 179.775,10.92
X$2055 576 8 577 644 645 cell_1rw
* cell instance $2056 m0 *1 180.48,10.92
X$2056 578 8 579 644 645 cell_1rw
* cell instance $2057 m0 *1 0.705,13.65
X$2057 67 9 68 644 645 cell_1rw
* cell instance $2058 m0 *1 0,13.65
X$2058 65 9 66 644 645 cell_1rw
* cell instance $2059 m0 *1 1.41,13.65
X$2059 69 9 70 644 645 cell_1rw
* cell instance $2060 m0 *1 2.115,13.65
X$2060 71 9 72 644 645 cell_1rw
* cell instance $2061 m0 *1 2.82,13.65
X$2061 73 9 74 644 645 cell_1rw
* cell instance $2062 m0 *1 3.525,13.65
X$2062 75 9 76 644 645 cell_1rw
* cell instance $2063 m0 *1 4.23,13.65
X$2063 77 9 78 644 645 cell_1rw
* cell instance $2064 m0 *1 4.935,13.65
X$2064 79 9 80 644 645 cell_1rw
* cell instance $2065 m0 *1 5.64,13.65
X$2065 81 9 82 644 645 cell_1rw
* cell instance $2066 m0 *1 6.345,13.65
X$2066 83 9 84 644 645 cell_1rw
* cell instance $2067 m0 *1 7.05,13.65
X$2067 85 9 86 644 645 cell_1rw
* cell instance $2068 m0 *1 7.755,13.65
X$2068 87 9 88 644 645 cell_1rw
* cell instance $2069 m0 *1 8.46,13.65
X$2069 89 9 90 644 645 cell_1rw
* cell instance $2070 m0 *1 9.165,13.65
X$2070 91 9 92 644 645 cell_1rw
* cell instance $2071 m0 *1 9.87,13.65
X$2071 93 9 94 644 645 cell_1rw
* cell instance $2072 m0 *1 10.575,13.65
X$2072 95 9 96 644 645 cell_1rw
* cell instance $2073 m0 *1 11.28,13.65
X$2073 97 9 98 644 645 cell_1rw
* cell instance $2074 m0 *1 11.985,13.65
X$2074 99 9 100 644 645 cell_1rw
* cell instance $2075 m0 *1 12.69,13.65
X$2075 101 9 102 644 645 cell_1rw
* cell instance $2076 m0 *1 13.395,13.65
X$2076 103 9 104 644 645 cell_1rw
* cell instance $2077 m0 *1 14.1,13.65
X$2077 105 9 106 644 645 cell_1rw
* cell instance $2078 m0 *1 14.805,13.65
X$2078 107 9 108 644 645 cell_1rw
* cell instance $2079 m0 *1 15.51,13.65
X$2079 109 9 110 644 645 cell_1rw
* cell instance $2080 m0 *1 16.215,13.65
X$2080 111 9 112 644 645 cell_1rw
* cell instance $2081 m0 *1 16.92,13.65
X$2081 113 9 114 644 645 cell_1rw
* cell instance $2082 m0 *1 17.625,13.65
X$2082 115 9 116 644 645 cell_1rw
* cell instance $2083 m0 *1 18.33,13.65
X$2083 117 9 118 644 645 cell_1rw
* cell instance $2084 m0 *1 19.035,13.65
X$2084 119 9 120 644 645 cell_1rw
* cell instance $2085 m0 *1 19.74,13.65
X$2085 121 9 122 644 645 cell_1rw
* cell instance $2086 m0 *1 20.445,13.65
X$2086 123 9 124 644 645 cell_1rw
* cell instance $2087 m0 *1 21.15,13.65
X$2087 125 9 126 644 645 cell_1rw
* cell instance $2088 m0 *1 21.855,13.65
X$2088 127 9 128 644 645 cell_1rw
* cell instance $2089 m0 *1 22.56,13.65
X$2089 129 9 130 644 645 cell_1rw
* cell instance $2090 m0 *1 23.265,13.65
X$2090 131 9 132 644 645 cell_1rw
* cell instance $2091 m0 *1 23.97,13.65
X$2091 133 9 134 644 645 cell_1rw
* cell instance $2092 m0 *1 24.675,13.65
X$2092 135 9 136 644 645 cell_1rw
* cell instance $2093 m0 *1 25.38,13.65
X$2093 137 9 138 644 645 cell_1rw
* cell instance $2094 m0 *1 26.085,13.65
X$2094 139 9 140 644 645 cell_1rw
* cell instance $2095 m0 *1 26.79,13.65
X$2095 141 9 142 644 645 cell_1rw
* cell instance $2096 m0 *1 27.495,13.65
X$2096 143 9 144 644 645 cell_1rw
* cell instance $2097 m0 *1 28.2,13.65
X$2097 145 9 146 644 645 cell_1rw
* cell instance $2098 m0 *1 28.905,13.65
X$2098 147 9 148 644 645 cell_1rw
* cell instance $2099 m0 *1 29.61,13.65
X$2099 149 9 150 644 645 cell_1rw
* cell instance $2100 m0 *1 30.315,13.65
X$2100 151 9 152 644 645 cell_1rw
* cell instance $2101 m0 *1 31.02,13.65
X$2101 153 9 154 644 645 cell_1rw
* cell instance $2102 m0 *1 31.725,13.65
X$2102 155 9 156 644 645 cell_1rw
* cell instance $2103 m0 *1 32.43,13.65
X$2103 157 9 158 644 645 cell_1rw
* cell instance $2104 m0 *1 33.135,13.65
X$2104 159 9 160 644 645 cell_1rw
* cell instance $2105 m0 *1 33.84,13.65
X$2105 161 9 162 644 645 cell_1rw
* cell instance $2106 m0 *1 34.545,13.65
X$2106 163 9 164 644 645 cell_1rw
* cell instance $2107 m0 *1 35.25,13.65
X$2107 165 9 166 644 645 cell_1rw
* cell instance $2108 m0 *1 35.955,13.65
X$2108 167 9 168 644 645 cell_1rw
* cell instance $2109 m0 *1 36.66,13.65
X$2109 169 9 170 644 645 cell_1rw
* cell instance $2110 m0 *1 37.365,13.65
X$2110 171 9 172 644 645 cell_1rw
* cell instance $2111 m0 *1 38.07,13.65
X$2111 173 9 174 644 645 cell_1rw
* cell instance $2112 m0 *1 38.775,13.65
X$2112 175 9 176 644 645 cell_1rw
* cell instance $2113 m0 *1 39.48,13.65
X$2113 177 9 178 644 645 cell_1rw
* cell instance $2114 m0 *1 40.185,13.65
X$2114 179 9 180 644 645 cell_1rw
* cell instance $2115 m0 *1 40.89,13.65
X$2115 181 9 182 644 645 cell_1rw
* cell instance $2116 m0 *1 41.595,13.65
X$2116 183 9 184 644 645 cell_1rw
* cell instance $2117 m0 *1 42.3,13.65
X$2117 185 9 186 644 645 cell_1rw
* cell instance $2118 m0 *1 43.005,13.65
X$2118 187 9 188 644 645 cell_1rw
* cell instance $2119 m0 *1 43.71,13.65
X$2119 189 9 190 644 645 cell_1rw
* cell instance $2120 m0 *1 44.415,13.65
X$2120 191 9 192 644 645 cell_1rw
* cell instance $2121 m0 *1 45.12,13.65
X$2121 193 9 194 644 645 cell_1rw
* cell instance $2122 m0 *1 45.825,13.65
X$2122 195 9 196 644 645 cell_1rw
* cell instance $2123 m0 *1 46.53,13.65
X$2123 197 9 198 644 645 cell_1rw
* cell instance $2124 m0 *1 47.235,13.65
X$2124 199 9 200 644 645 cell_1rw
* cell instance $2125 m0 *1 47.94,13.65
X$2125 201 9 202 644 645 cell_1rw
* cell instance $2126 m0 *1 48.645,13.65
X$2126 203 9 204 644 645 cell_1rw
* cell instance $2127 m0 *1 49.35,13.65
X$2127 205 9 206 644 645 cell_1rw
* cell instance $2128 m0 *1 50.055,13.65
X$2128 207 9 208 644 645 cell_1rw
* cell instance $2129 m0 *1 50.76,13.65
X$2129 209 9 210 644 645 cell_1rw
* cell instance $2130 m0 *1 51.465,13.65
X$2130 211 9 212 644 645 cell_1rw
* cell instance $2131 m0 *1 52.17,13.65
X$2131 213 9 214 644 645 cell_1rw
* cell instance $2132 m0 *1 52.875,13.65
X$2132 215 9 216 644 645 cell_1rw
* cell instance $2133 m0 *1 53.58,13.65
X$2133 217 9 218 644 645 cell_1rw
* cell instance $2134 m0 *1 54.285,13.65
X$2134 219 9 220 644 645 cell_1rw
* cell instance $2135 m0 *1 54.99,13.65
X$2135 221 9 222 644 645 cell_1rw
* cell instance $2136 m0 *1 55.695,13.65
X$2136 223 9 224 644 645 cell_1rw
* cell instance $2137 m0 *1 56.4,13.65
X$2137 225 9 226 644 645 cell_1rw
* cell instance $2138 m0 *1 57.105,13.65
X$2138 227 9 228 644 645 cell_1rw
* cell instance $2139 m0 *1 57.81,13.65
X$2139 229 9 230 644 645 cell_1rw
* cell instance $2140 m0 *1 58.515,13.65
X$2140 231 9 232 644 645 cell_1rw
* cell instance $2141 m0 *1 59.22,13.65
X$2141 233 9 234 644 645 cell_1rw
* cell instance $2142 m0 *1 59.925,13.65
X$2142 235 9 236 644 645 cell_1rw
* cell instance $2143 m0 *1 60.63,13.65
X$2143 237 9 238 644 645 cell_1rw
* cell instance $2144 m0 *1 61.335,13.65
X$2144 239 9 240 644 645 cell_1rw
* cell instance $2145 m0 *1 62.04,13.65
X$2145 241 9 242 644 645 cell_1rw
* cell instance $2146 m0 *1 62.745,13.65
X$2146 243 9 244 644 645 cell_1rw
* cell instance $2147 m0 *1 63.45,13.65
X$2147 245 9 246 644 645 cell_1rw
* cell instance $2148 m0 *1 64.155,13.65
X$2148 247 9 248 644 645 cell_1rw
* cell instance $2149 m0 *1 64.86,13.65
X$2149 249 9 250 644 645 cell_1rw
* cell instance $2150 m0 *1 65.565,13.65
X$2150 251 9 252 644 645 cell_1rw
* cell instance $2151 m0 *1 66.27,13.65
X$2151 253 9 254 644 645 cell_1rw
* cell instance $2152 m0 *1 66.975,13.65
X$2152 255 9 256 644 645 cell_1rw
* cell instance $2153 m0 *1 67.68,13.65
X$2153 257 9 258 644 645 cell_1rw
* cell instance $2154 m0 *1 68.385,13.65
X$2154 259 9 260 644 645 cell_1rw
* cell instance $2155 m0 *1 69.09,13.65
X$2155 261 9 262 644 645 cell_1rw
* cell instance $2156 m0 *1 69.795,13.65
X$2156 263 9 264 644 645 cell_1rw
* cell instance $2157 m0 *1 70.5,13.65
X$2157 265 9 266 644 645 cell_1rw
* cell instance $2158 m0 *1 71.205,13.65
X$2158 267 9 268 644 645 cell_1rw
* cell instance $2159 m0 *1 71.91,13.65
X$2159 269 9 270 644 645 cell_1rw
* cell instance $2160 m0 *1 72.615,13.65
X$2160 271 9 272 644 645 cell_1rw
* cell instance $2161 m0 *1 73.32,13.65
X$2161 273 9 274 644 645 cell_1rw
* cell instance $2162 m0 *1 74.025,13.65
X$2162 275 9 276 644 645 cell_1rw
* cell instance $2163 m0 *1 74.73,13.65
X$2163 277 9 278 644 645 cell_1rw
* cell instance $2164 m0 *1 75.435,13.65
X$2164 279 9 280 644 645 cell_1rw
* cell instance $2165 m0 *1 76.14,13.65
X$2165 281 9 282 644 645 cell_1rw
* cell instance $2166 m0 *1 76.845,13.65
X$2166 283 9 284 644 645 cell_1rw
* cell instance $2167 m0 *1 77.55,13.65
X$2167 285 9 286 644 645 cell_1rw
* cell instance $2168 m0 *1 78.255,13.65
X$2168 287 9 288 644 645 cell_1rw
* cell instance $2169 m0 *1 78.96,13.65
X$2169 289 9 290 644 645 cell_1rw
* cell instance $2170 m0 *1 79.665,13.65
X$2170 291 9 292 644 645 cell_1rw
* cell instance $2171 m0 *1 80.37,13.65
X$2171 293 9 294 644 645 cell_1rw
* cell instance $2172 m0 *1 81.075,13.65
X$2172 295 9 296 644 645 cell_1rw
* cell instance $2173 m0 *1 81.78,13.65
X$2173 297 9 298 644 645 cell_1rw
* cell instance $2174 m0 *1 82.485,13.65
X$2174 299 9 300 644 645 cell_1rw
* cell instance $2175 m0 *1 83.19,13.65
X$2175 301 9 302 644 645 cell_1rw
* cell instance $2176 m0 *1 83.895,13.65
X$2176 303 9 304 644 645 cell_1rw
* cell instance $2177 m0 *1 84.6,13.65
X$2177 305 9 306 644 645 cell_1rw
* cell instance $2178 m0 *1 85.305,13.65
X$2178 307 9 308 644 645 cell_1rw
* cell instance $2179 m0 *1 86.01,13.65
X$2179 309 9 310 644 645 cell_1rw
* cell instance $2180 m0 *1 86.715,13.65
X$2180 311 9 312 644 645 cell_1rw
* cell instance $2181 m0 *1 87.42,13.65
X$2181 313 9 314 644 645 cell_1rw
* cell instance $2182 m0 *1 88.125,13.65
X$2182 315 9 316 644 645 cell_1rw
* cell instance $2183 m0 *1 88.83,13.65
X$2183 317 9 318 644 645 cell_1rw
* cell instance $2184 m0 *1 89.535,13.65
X$2184 319 9 320 644 645 cell_1rw
* cell instance $2185 m0 *1 90.24,13.65
X$2185 321 9 323 644 645 cell_1rw
* cell instance $2186 m0 *1 90.945,13.65
X$2186 324 9 325 644 645 cell_1rw
* cell instance $2187 m0 *1 91.65,13.65
X$2187 326 9 327 644 645 cell_1rw
* cell instance $2188 m0 *1 92.355,13.65
X$2188 328 9 329 644 645 cell_1rw
* cell instance $2189 m0 *1 93.06,13.65
X$2189 330 9 331 644 645 cell_1rw
* cell instance $2190 m0 *1 93.765,13.65
X$2190 332 9 333 644 645 cell_1rw
* cell instance $2191 m0 *1 94.47,13.65
X$2191 334 9 335 644 645 cell_1rw
* cell instance $2192 m0 *1 95.175,13.65
X$2192 336 9 337 644 645 cell_1rw
* cell instance $2193 m0 *1 95.88,13.65
X$2193 338 9 339 644 645 cell_1rw
* cell instance $2194 m0 *1 96.585,13.65
X$2194 340 9 341 644 645 cell_1rw
* cell instance $2195 m0 *1 97.29,13.65
X$2195 342 9 343 644 645 cell_1rw
* cell instance $2196 m0 *1 97.995,13.65
X$2196 344 9 345 644 645 cell_1rw
* cell instance $2197 m0 *1 98.7,13.65
X$2197 346 9 347 644 645 cell_1rw
* cell instance $2198 m0 *1 99.405,13.65
X$2198 348 9 349 644 645 cell_1rw
* cell instance $2199 m0 *1 100.11,13.65
X$2199 350 9 351 644 645 cell_1rw
* cell instance $2200 m0 *1 100.815,13.65
X$2200 352 9 353 644 645 cell_1rw
* cell instance $2201 m0 *1 101.52,13.65
X$2201 354 9 355 644 645 cell_1rw
* cell instance $2202 m0 *1 102.225,13.65
X$2202 356 9 357 644 645 cell_1rw
* cell instance $2203 m0 *1 102.93,13.65
X$2203 358 9 359 644 645 cell_1rw
* cell instance $2204 m0 *1 103.635,13.65
X$2204 360 9 361 644 645 cell_1rw
* cell instance $2205 m0 *1 104.34,13.65
X$2205 362 9 363 644 645 cell_1rw
* cell instance $2206 m0 *1 105.045,13.65
X$2206 364 9 365 644 645 cell_1rw
* cell instance $2207 m0 *1 105.75,13.65
X$2207 366 9 367 644 645 cell_1rw
* cell instance $2208 m0 *1 106.455,13.65
X$2208 368 9 369 644 645 cell_1rw
* cell instance $2209 m0 *1 107.16,13.65
X$2209 370 9 371 644 645 cell_1rw
* cell instance $2210 m0 *1 107.865,13.65
X$2210 372 9 373 644 645 cell_1rw
* cell instance $2211 m0 *1 108.57,13.65
X$2211 374 9 375 644 645 cell_1rw
* cell instance $2212 m0 *1 109.275,13.65
X$2212 376 9 377 644 645 cell_1rw
* cell instance $2213 m0 *1 109.98,13.65
X$2213 378 9 379 644 645 cell_1rw
* cell instance $2214 m0 *1 110.685,13.65
X$2214 380 9 381 644 645 cell_1rw
* cell instance $2215 m0 *1 111.39,13.65
X$2215 382 9 383 644 645 cell_1rw
* cell instance $2216 m0 *1 112.095,13.65
X$2216 384 9 385 644 645 cell_1rw
* cell instance $2217 m0 *1 112.8,13.65
X$2217 386 9 387 644 645 cell_1rw
* cell instance $2218 m0 *1 113.505,13.65
X$2218 388 9 389 644 645 cell_1rw
* cell instance $2219 m0 *1 114.21,13.65
X$2219 390 9 391 644 645 cell_1rw
* cell instance $2220 m0 *1 114.915,13.65
X$2220 392 9 393 644 645 cell_1rw
* cell instance $2221 m0 *1 115.62,13.65
X$2221 394 9 395 644 645 cell_1rw
* cell instance $2222 m0 *1 116.325,13.65
X$2222 396 9 397 644 645 cell_1rw
* cell instance $2223 m0 *1 117.03,13.65
X$2223 398 9 399 644 645 cell_1rw
* cell instance $2224 m0 *1 117.735,13.65
X$2224 400 9 401 644 645 cell_1rw
* cell instance $2225 m0 *1 118.44,13.65
X$2225 402 9 403 644 645 cell_1rw
* cell instance $2226 m0 *1 119.145,13.65
X$2226 404 9 405 644 645 cell_1rw
* cell instance $2227 m0 *1 119.85,13.65
X$2227 406 9 407 644 645 cell_1rw
* cell instance $2228 m0 *1 120.555,13.65
X$2228 408 9 409 644 645 cell_1rw
* cell instance $2229 m0 *1 121.26,13.65
X$2229 410 9 411 644 645 cell_1rw
* cell instance $2230 m0 *1 121.965,13.65
X$2230 412 9 413 644 645 cell_1rw
* cell instance $2231 m0 *1 122.67,13.65
X$2231 414 9 415 644 645 cell_1rw
* cell instance $2232 m0 *1 123.375,13.65
X$2232 416 9 417 644 645 cell_1rw
* cell instance $2233 m0 *1 124.08,13.65
X$2233 418 9 419 644 645 cell_1rw
* cell instance $2234 m0 *1 124.785,13.65
X$2234 420 9 421 644 645 cell_1rw
* cell instance $2235 m0 *1 125.49,13.65
X$2235 422 9 423 644 645 cell_1rw
* cell instance $2236 m0 *1 126.195,13.65
X$2236 424 9 425 644 645 cell_1rw
* cell instance $2237 m0 *1 126.9,13.65
X$2237 426 9 427 644 645 cell_1rw
* cell instance $2238 m0 *1 127.605,13.65
X$2238 428 9 429 644 645 cell_1rw
* cell instance $2239 m0 *1 128.31,13.65
X$2239 430 9 431 644 645 cell_1rw
* cell instance $2240 m0 *1 129.015,13.65
X$2240 432 9 433 644 645 cell_1rw
* cell instance $2241 m0 *1 129.72,13.65
X$2241 434 9 435 644 645 cell_1rw
* cell instance $2242 m0 *1 130.425,13.65
X$2242 436 9 437 644 645 cell_1rw
* cell instance $2243 m0 *1 131.13,13.65
X$2243 438 9 439 644 645 cell_1rw
* cell instance $2244 m0 *1 131.835,13.65
X$2244 440 9 441 644 645 cell_1rw
* cell instance $2245 m0 *1 132.54,13.65
X$2245 442 9 443 644 645 cell_1rw
* cell instance $2246 m0 *1 133.245,13.65
X$2246 444 9 445 644 645 cell_1rw
* cell instance $2247 m0 *1 133.95,13.65
X$2247 446 9 447 644 645 cell_1rw
* cell instance $2248 m0 *1 134.655,13.65
X$2248 448 9 449 644 645 cell_1rw
* cell instance $2249 m0 *1 135.36,13.65
X$2249 450 9 451 644 645 cell_1rw
* cell instance $2250 m0 *1 136.065,13.65
X$2250 452 9 453 644 645 cell_1rw
* cell instance $2251 m0 *1 136.77,13.65
X$2251 454 9 455 644 645 cell_1rw
* cell instance $2252 m0 *1 137.475,13.65
X$2252 456 9 457 644 645 cell_1rw
* cell instance $2253 m0 *1 138.18,13.65
X$2253 458 9 459 644 645 cell_1rw
* cell instance $2254 m0 *1 138.885,13.65
X$2254 460 9 461 644 645 cell_1rw
* cell instance $2255 m0 *1 139.59,13.65
X$2255 462 9 463 644 645 cell_1rw
* cell instance $2256 m0 *1 140.295,13.65
X$2256 464 9 465 644 645 cell_1rw
* cell instance $2257 m0 *1 141,13.65
X$2257 466 9 467 644 645 cell_1rw
* cell instance $2258 m0 *1 141.705,13.65
X$2258 468 9 469 644 645 cell_1rw
* cell instance $2259 m0 *1 142.41,13.65
X$2259 470 9 471 644 645 cell_1rw
* cell instance $2260 m0 *1 143.115,13.65
X$2260 472 9 473 644 645 cell_1rw
* cell instance $2261 m0 *1 143.82,13.65
X$2261 474 9 475 644 645 cell_1rw
* cell instance $2262 m0 *1 144.525,13.65
X$2262 476 9 477 644 645 cell_1rw
* cell instance $2263 m0 *1 145.23,13.65
X$2263 478 9 479 644 645 cell_1rw
* cell instance $2264 m0 *1 145.935,13.65
X$2264 480 9 481 644 645 cell_1rw
* cell instance $2265 m0 *1 146.64,13.65
X$2265 482 9 483 644 645 cell_1rw
* cell instance $2266 m0 *1 147.345,13.65
X$2266 484 9 485 644 645 cell_1rw
* cell instance $2267 m0 *1 148.05,13.65
X$2267 486 9 487 644 645 cell_1rw
* cell instance $2268 m0 *1 148.755,13.65
X$2268 488 9 489 644 645 cell_1rw
* cell instance $2269 m0 *1 149.46,13.65
X$2269 490 9 491 644 645 cell_1rw
* cell instance $2270 m0 *1 150.165,13.65
X$2270 492 9 493 644 645 cell_1rw
* cell instance $2271 m0 *1 150.87,13.65
X$2271 494 9 495 644 645 cell_1rw
* cell instance $2272 m0 *1 151.575,13.65
X$2272 496 9 497 644 645 cell_1rw
* cell instance $2273 m0 *1 152.28,13.65
X$2273 498 9 499 644 645 cell_1rw
* cell instance $2274 m0 *1 152.985,13.65
X$2274 500 9 501 644 645 cell_1rw
* cell instance $2275 m0 *1 153.69,13.65
X$2275 502 9 503 644 645 cell_1rw
* cell instance $2276 m0 *1 154.395,13.65
X$2276 504 9 505 644 645 cell_1rw
* cell instance $2277 m0 *1 155.1,13.65
X$2277 506 9 507 644 645 cell_1rw
* cell instance $2278 m0 *1 155.805,13.65
X$2278 508 9 509 644 645 cell_1rw
* cell instance $2279 m0 *1 156.51,13.65
X$2279 510 9 511 644 645 cell_1rw
* cell instance $2280 m0 *1 157.215,13.65
X$2280 512 9 513 644 645 cell_1rw
* cell instance $2281 m0 *1 157.92,13.65
X$2281 514 9 515 644 645 cell_1rw
* cell instance $2282 m0 *1 158.625,13.65
X$2282 516 9 517 644 645 cell_1rw
* cell instance $2283 m0 *1 159.33,13.65
X$2283 518 9 519 644 645 cell_1rw
* cell instance $2284 m0 *1 160.035,13.65
X$2284 520 9 521 644 645 cell_1rw
* cell instance $2285 m0 *1 160.74,13.65
X$2285 522 9 523 644 645 cell_1rw
* cell instance $2286 m0 *1 161.445,13.65
X$2286 524 9 525 644 645 cell_1rw
* cell instance $2287 m0 *1 162.15,13.65
X$2287 526 9 527 644 645 cell_1rw
* cell instance $2288 m0 *1 162.855,13.65
X$2288 528 9 529 644 645 cell_1rw
* cell instance $2289 m0 *1 163.56,13.65
X$2289 530 9 531 644 645 cell_1rw
* cell instance $2290 m0 *1 164.265,13.65
X$2290 532 9 533 644 645 cell_1rw
* cell instance $2291 m0 *1 164.97,13.65
X$2291 534 9 535 644 645 cell_1rw
* cell instance $2292 m0 *1 165.675,13.65
X$2292 536 9 537 644 645 cell_1rw
* cell instance $2293 m0 *1 166.38,13.65
X$2293 538 9 539 644 645 cell_1rw
* cell instance $2294 m0 *1 167.085,13.65
X$2294 540 9 541 644 645 cell_1rw
* cell instance $2295 m0 *1 167.79,13.65
X$2295 542 9 543 644 645 cell_1rw
* cell instance $2296 m0 *1 168.495,13.65
X$2296 544 9 545 644 645 cell_1rw
* cell instance $2297 m0 *1 169.2,13.65
X$2297 546 9 547 644 645 cell_1rw
* cell instance $2298 m0 *1 169.905,13.65
X$2298 548 9 549 644 645 cell_1rw
* cell instance $2299 m0 *1 170.61,13.65
X$2299 550 9 551 644 645 cell_1rw
* cell instance $2300 m0 *1 171.315,13.65
X$2300 552 9 553 644 645 cell_1rw
* cell instance $2301 m0 *1 172.02,13.65
X$2301 554 9 555 644 645 cell_1rw
* cell instance $2302 m0 *1 172.725,13.65
X$2302 556 9 557 644 645 cell_1rw
* cell instance $2303 m0 *1 173.43,13.65
X$2303 558 9 559 644 645 cell_1rw
* cell instance $2304 m0 *1 174.135,13.65
X$2304 560 9 561 644 645 cell_1rw
* cell instance $2305 m0 *1 174.84,13.65
X$2305 562 9 563 644 645 cell_1rw
* cell instance $2306 m0 *1 175.545,13.65
X$2306 564 9 565 644 645 cell_1rw
* cell instance $2307 m0 *1 176.25,13.65
X$2307 566 9 567 644 645 cell_1rw
* cell instance $2308 m0 *1 176.955,13.65
X$2308 568 9 569 644 645 cell_1rw
* cell instance $2309 m0 *1 177.66,13.65
X$2309 570 9 571 644 645 cell_1rw
* cell instance $2310 m0 *1 178.365,13.65
X$2310 572 9 573 644 645 cell_1rw
* cell instance $2311 m0 *1 179.07,13.65
X$2311 574 9 575 644 645 cell_1rw
* cell instance $2312 m0 *1 179.775,13.65
X$2312 576 9 577 644 645 cell_1rw
* cell instance $2313 m0 *1 180.48,13.65
X$2313 578 9 579 644 645 cell_1rw
* cell instance $2314 r0 *1 0.705,10.92
X$2314 67 10 68 644 645 cell_1rw
* cell instance $2315 r0 *1 0,10.92
X$2315 65 10 66 644 645 cell_1rw
* cell instance $2316 r0 *1 1.41,10.92
X$2316 69 10 70 644 645 cell_1rw
* cell instance $2317 r0 *1 2.115,10.92
X$2317 71 10 72 644 645 cell_1rw
* cell instance $2318 r0 *1 2.82,10.92
X$2318 73 10 74 644 645 cell_1rw
* cell instance $2319 r0 *1 3.525,10.92
X$2319 75 10 76 644 645 cell_1rw
* cell instance $2320 r0 *1 4.23,10.92
X$2320 77 10 78 644 645 cell_1rw
* cell instance $2321 r0 *1 4.935,10.92
X$2321 79 10 80 644 645 cell_1rw
* cell instance $2322 r0 *1 5.64,10.92
X$2322 81 10 82 644 645 cell_1rw
* cell instance $2323 r0 *1 6.345,10.92
X$2323 83 10 84 644 645 cell_1rw
* cell instance $2324 r0 *1 7.05,10.92
X$2324 85 10 86 644 645 cell_1rw
* cell instance $2325 r0 *1 7.755,10.92
X$2325 87 10 88 644 645 cell_1rw
* cell instance $2326 r0 *1 8.46,10.92
X$2326 89 10 90 644 645 cell_1rw
* cell instance $2327 r0 *1 9.165,10.92
X$2327 91 10 92 644 645 cell_1rw
* cell instance $2328 r0 *1 9.87,10.92
X$2328 93 10 94 644 645 cell_1rw
* cell instance $2329 r0 *1 10.575,10.92
X$2329 95 10 96 644 645 cell_1rw
* cell instance $2330 r0 *1 11.28,10.92
X$2330 97 10 98 644 645 cell_1rw
* cell instance $2331 r0 *1 11.985,10.92
X$2331 99 10 100 644 645 cell_1rw
* cell instance $2332 r0 *1 12.69,10.92
X$2332 101 10 102 644 645 cell_1rw
* cell instance $2333 r0 *1 13.395,10.92
X$2333 103 10 104 644 645 cell_1rw
* cell instance $2334 r0 *1 14.1,10.92
X$2334 105 10 106 644 645 cell_1rw
* cell instance $2335 r0 *1 14.805,10.92
X$2335 107 10 108 644 645 cell_1rw
* cell instance $2336 r0 *1 15.51,10.92
X$2336 109 10 110 644 645 cell_1rw
* cell instance $2337 r0 *1 16.215,10.92
X$2337 111 10 112 644 645 cell_1rw
* cell instance $2338 r0 *1 16.92,10.92
X$2338 113 10 114 644 645 cell_1rw
* cell instance $2339 r0 *1 17.625,10.92
X$2339 115 10 116 644 645 cell_1rw
* cell instance $2340 r0 *1 18.33,10.92
X$2340 117 10 118 644 645 cell_1rw
* cell instance $2341 r0 *1 19.035,10.92
X$2341 119 10 120 644 645 cell_1rw
* cell instance $2342 r0 *1 19.74,10.92
X$2342 121 10 122 644 645 cell_1rw
* cell instance $2343 r0 *1 20.445,10.92
X$2343 123 10 124 644 645 cell_1rw
* cell instance $2344 r0 *1 21.15,10.92
X$2344 125 10 126 644 645 cell_1rw
* cell instance $2345 r0 *1 21.855,10.92
X$2345 127 10 128 644 645 cell_1rw
* cell instance $2346 r0 *1 22.56,10.92
X$2346 129 10 130 644 645 cell_1rw
* cell instance $2347 r0 *1 23.265,10.92
X$2347 131 10 132 644 645 cell_1rw
* cell instance $2348 r0 *1 23.97,10.92
X$2348 133 10 134 644 645 cell_1rw
* cell instance $2349 r0 *1 24.675,10.92
X$2349 135 10 136 644 645 cell_1rw
* cell instance $2350 r0 *1 25.38,10.92
X$2350 137 10 138 644 645 cell_1rw
* cell instance $2351 r0 *1 26.085,10.92
X$2351 139 10 140 644 645 cell_1rw
* cell instance $2352 r0 *1 26.79,10.92
X$2352 141 10 142 644 645 cell_1rw
* cell instance $2353 r0 *1 27.495,10.92
X$2353 143 10 144 644 645 cell_1rw
* cell instance $2354 r0 *1 28.2,10.92
X$2354 145 10 146 644 645 cell_1rw
* cell instance $2355 r0 *1 28.905,10.92
X$2355 147 10 148 644 645 cell_1rw
* cell instance $2356 r0 *1 29.61,10.92
X$2356 149 10 150 644 645 cell_1rw
* cell instance $2357 r0 *1 30.315,10.92
X$2357 151 10 152 644 645 cell_1rw
* cell instance $2358 r0 *1 31.02,10.92
X$2358 153 10 154 644 645 cell_1rw
* cell instance $2359 r0 *1 31.725,10.92
X$2359 155 10 156 644 645 cell_1rw
* cell instance $2360 r0 *1 32.43,10.92
X$2360 157 10 158 644 645 cell_1rw
* cell instance $2361 r0 *1 33.135,10.92
X$2361 159 10 160 644 645 cell_1rw
* cell instance $2362 r0 *1 33.84,10.92
X$2362 161 10 162 644 645 cell_1rw
* cell instance $2363 r0 *1 34.545,10.92
X$2363 163 10 164 644 645 cell_1rw
* cell instance $2364 r0 *1 35.25,10.92
X$2364 165 10 166 644 645 cell_1rw
* cell instance $2365 r0 *1 35.955,10.92
X$2365 167 10 168 644 645 cell_1rw
* cell instance $2366 r0 *1 36.66,10.92
X$2366 169 10 170 644 645 cell_1rw
* cell instance $2367 r0 *1 37.365,10.92
X$2367 171 10 172 644 645 cell_1rw
* cell instance $2368 r0 *1 38.07,10.92
X$2368 173 10 174 644 645 cell_1rw
* cell instance $2369 r0 *1 38.775,10.92
X$2369 175 10 176 644 645 cell_1rw
* cell instance $2370 r0 *1 39.48,10.92
X$2370 177 10 178 644 645 cell_1rw
* cell instance $2371 r0 *1 40.185,10.92
X$2371 179 10 180 644 645 cell_1rw
* cell instance $2372 r0 *1 40.89,10.92
X$2372 181 10 182 644 645 cell_1rw
* cell instance $2373 r0 *1 41.595,10.92
X$2373 183 10 184 644 645 cell_1rw
* cell instance $2374 r0 *1 42.3,10.92
X$2374 185 10 186 644 645 cell_1rw
* cell instance $2375 r0 *1 43.005,10.92
X$2375 187 10 188 644 645 cell_1rw
* cell instance $2376 r0 *1 43.71,10.92
X$2376 189 10 190 644 645 cell_1rw
* cell instance $2377 r0 *1 44.415,10.92
X$2377 191 10 192 644 645 cell_1rw
* cell instance $2378 r0 *1 45.12,10.92
X$2378 193 10 194 644 645 cell_1rw
* cell instance $2379 r0 *1 45.825,10.92
X$2379 195 10 196 644 645 cell_1rw
* cell instance $2380 r0 *1 46.53,10.92
X$2380 197 10 198 644 645 cell_1rw
* cell instance $2381 r0 *1 47.235,10.92
X$2381 199 10 200 644 645 cell_1rw
* cell instance $2382 r0 *1 47.94,10.92
X$2382 201 10 202 644 645 cell_1rw
* cell instance $2383 r0 *1 48.645,10.92
X$2383 203 10 204 644 645 cell_1rw
* cell instance $2384 r0 *1 49.35,10.92
X$2384 205 10 206 644 645 cell_1rw
* cell instance $2385 r0 *1 50.055,10.92
X$2385 207 10 208 644 645 cell_1rw
* cell instance $2386 r0 *1 50.76,10.92
X$2386 209 10 210 644 645 cell_1rw
* cell instance $2387 r0 *1 51.465,10.92
X$2387 211 10 212 644 645 cell_1rw
* cell instance $2388 r0 *1 52.17,10.92
X$2388 213 10 214 644 645 cell_1rw
* cell instance $2389 r0 *1 52.875,10.92
X$2389 215 10 216 644 645 cell_1rw
* cell instance $2390 r0 *1 53.58,10.92
X$2390 217 10 218 644 645 cell_1rw
* cell instance $2391 r0 *1 54.285,10.92
X$2391 219 10 220 644 645 cell_1rw
* cell instance $2392 r0 *1 54.99,10.92
X$2392 221 10 222 644 645 cell_1rw
* cell instance $2393 r0 *1 55.695,10.92
X$2393 223 10 224 644 645 cell_1rw
* cell instance $2394 r0 *1 56.4,10.92
X$2394 225 10 226 644 645 cell_1rw
* cell instance $2395 r0 *1 57.105,10.92
X$2395 227 10 228 644 645 cell_1rw
* cell instance $2396 r0 *1 57.81,10.92
X$2396 229 10 230 644 645 cell_1rw
* cell instance $2397 r0 *1 58.515,10.92
X$2397 231 10 232 644 645 cell_1rw
* cell instance $2398 r0 *1 59.22,10.92
X$2398 233 10 234 644 645 cell_1rw
* cell instance $2399 r0 *1 59.925,10.92
X$2399 235 10 236 644 645 cell_1rw
* cell instance $2400 r0 *1 60.63,10.92
X$2400 237 10 238 644 645 cell_1rw
* cell instance $2401 r0 *1 61.335,10.92
X$2401 239 10 240 644 645 cell_1rw
* cell instance $2402 r0 *1 62.04,10.92
X$2402 241 10 242 644 645 cell_1rw
* cell instance $2403 r0 *1 62.745,10.92
X$2403 243 10 244 644 645 cell_1rw
* cell instance $2404 r0 *1 63.45,10.92
X$2404 245 10 246 644 645 cell_1rw
* cell instance $2405 r0 *1 64.155,10.92
X$2405 247 10 248 644 645 cell_1rw
* cell instance $2406 r0 *1 64.86,10.92
X$2406 249 10 250 644 645 cell_1rw
* cell instance $2407 r0 *1 65.565,10.92
X$2407 251 10 252 644 645 cell_1rw
* cell instance $2408 r0 *1 66.27,10.92
X$2408 253 10 254 644 645 cell_1rw
* cell instance $2409 r0 *1 66.975,10.92
X$2409 255 10 256 644 645 cell_1rw
* cell instance $2410 r0 *1 67.68,10.92
X$2410 257 10 258 644 645 cell_1rw
* cell instance $2411 r0 *1 68.385,10.92
X$2411 259 10 260 644 645 cell_1rw
* cell instance $2412 r0 *1 69.09,10.92
X$2412 261 10 262 644 645 cell_1rw
* cell instance $2413 r0 *1 69.795,10.92
X$2413 263 10 264 644 645 cell_1rw
* cell instance $2414 r0 *1 70.5,10.92
X$2414 265 10 266 644 645 cell_1rw
* cell instance $2415 r0 *1 71.205,10.92
X$2415 267 10 268 644 645 cell_1rw
* cell instance $2416 r0 *1 71.91,10.92
X$2416 269 10 270 644 645 cell_1rw
* cell instance $2417 r0 *1 72.615,10.92
X$2417 271 10 272 644 645 cell_1rw
* cell instance $2418 r0 *1 73.32,10.92
X$2418 273 10 274 644 645 cell_1rw
* cell instance $2419 r0 *1 74.025,10.92
X$2419 275 10 276 644 645 cell_1rw
* cell instance $2420 r0 *1 74.73,10.92
X$2420 277 10 278 644 645 cell_1rw
* cell instance $2421 r0 *1 75.435,10.92
X$2421 279 10 280 644 645 cell_1rw
* cell instance $2422 r0 *1 76.14,10.92
X$2422 281 10 282 644 645 cell_1rw
* cell instance $2423 r0 *1 76.845,10.92
X$2423 283 10 284 644 645 cell_1rw
* cell instance $2424 r0 *1 77.55,10.92
X$2424 285 10 286 644 645 cell_1rw
* cell instance $2425 r0 *1 78.255,10.92
X$2425 287 10 288 644 645 cell_1rw
* cell instance $2426 r0 *1 78.96,10.92
X$2426 289 10 290 644 645 cell_1rw
* cell instance $2427 r0 *1 79.665,10.92
X$2427 291 10 292 644 645 cell_1rw
* cell instance $2428 r0 *1 80.37,10.92
X$2428 293 10 294 644 645 cell_1rw
* cell instance $2429 r0 *1 81.075,10.92
X$2429 295 10 296 644 645 cell_1rw
* cell instance $2430 r0 *1 81.78,10.92
X$2430 297 10 298 644 645 cell_1rw
* cell instance $2431 r0 *1 82.485,10.92
X$2431 299 10 300 644 645 cell_1rw
* cell instance $2432 r0 *1 83.19,10.92
X$2432 301 10 302 644 645 cell_1rw
* cell instance $2433 r0 *1 83.895,10.92
X$2433 303 10 304 644 645 cell_1rw
* cell instance $2434 r0 *1 84.6,10.92
X$2434 305 10 306 644 645 cell_1rw
* cell instance $2435 r0 *1 85.305,10.92
X$2435 307 10 308 644 645 cell_1rw
* cell instance $2436 r0 *1 86.01,10.92
X$2436 309 10 310 644 645 cell_1rw
* cell instance $2437 r0 *1 86.715,10.92
X$2437 311 10 312 644 645 cell_1rw
* cell instance $2438 r0 *1 87.42,10.92
X$2438 313 10 314 644 645 cell_1rw
* cell instance $2439 r0 *1 88.125,10.92
X$2439 315 10 316 644 645 cell_1rw
* cell instance $2440 r0 *1 88.83,10.92
X$2440 317 10 318 644 645 cell_1rw
* cell instance $2441 r0 *1 89.535,10.92
X$2441 319 10 320 644 645 cell_1rw
* cell instance $2442 r0 *1 90.24,10.92
X$2442 321 10 323 644 645 cell_1rw
* cell instance $2443 r0 *1 90.945,10.92
X$2443 324 10 325 644 645 cell_1rw
* cell instance $2444 r0 *1 91.65,10.92
X$2444 326 10 327 644 645 cell_1rw
* cell instance $2445 r0 *1 92.355,10.92
X$2445 328 10 329 644 645 cell_1rw
* cell instance $2446 r0 *1 93.06,10.92
X$2446 330 10 331 644 645 cell_1rw
* cell instance $2447 r0 *1 93.765,10.92
X$2447 332 10 333 644 645 cell_1rw
* cell instance $2448 r0 *1 94.47,10.92
X$2448 334 10 335 644 645 cell_1rw
* cell instance $2449 r0 *1 95.175,10.92
X$2449 336 10 337 644 645 cell_1rw
* cell instance $2450 r0 *1 95.88,10.92
X$2450 338 10 339 644 645 cell_1rw
* cell instance $2451 r0 *1 96.585,10.92
X$2451 340 10 341 644 645 cell_1rw
* cell instance $2452 r0 *1 97.29,10.92
X$2452 342 10 343 644 645 cell_1rw
* cell instance $2453 r0 *1 97.995,10.92
X$2453 344 10 345 644 645 cell_1rw
* cell instance $2454 r0 *1 98.7,10.92
X$2454 346 10 347 644 645 cell_1rw
* cell instance $2455 r0 *1 99.405,10.92
X$2455 348 10 349 644 645 cell_1rw
* cell instance $2456 r0 *1 100.11,10.92
X$2456 350 10 351 644 645 cell_1rw
* cell instance $2457 r0 *1 100.815,10.92
X$2457 352 10 353 644 645 cell_1rw
* cell instance $2458 r0 *1 101.52,10.92
X$2458 354 10 355 644 645 cell_1rw
* cell instance $2459 r0 *1 102.225,10.92
X$2459 356 10 357 644 645 cell_1rw
* cell instance $2460 r0 *1 102.93,10.92
X$2460 358 10 359 644 645 cell_1rw
* cell instance $2461 r0 *1 103.635,10.92
X$2461 360 10 361 644 645 cell_1rw
* cell instance $2462 r0 *1 104.34,10.92
X$2462 362 10 363 644 645 cell_1rw
* cell instance $2463 r0 *1 105.045,10.92
X$2463 364 10 365 644 645 cell_1rw
* cell instance $2464 r0 *1 105.75,10.92
X$2464 366 10 367 644 645 cell_1rw
* cell instance $2465 r0 *1 106.455,10.92
X$2465 368 10 369 644 645 cell_1rw
* cell instance $2466 r0 *1 107.16,10.92
X$2466 370 10 371 644 645 cell_1rw
* cell instance $2467 r0 *1 107.865,10.92
X$2467 372 10 373 644 645 cell_1rw
* cell instance $2468 r0 *1 108.57,10.92
X$2468 374 10 375 644 645 cell_1rw
* cell instance $2469 r0 *1 109.275,10.92
X$2469 376 10 377 644 645 cell_1rw
* cell instance $2470 r0 *1 109.98,10.92
X$2470 378 10 379 644 645 cell_1rw
* cell instance $2471 r0 *1 110.685,10.92
X$2471 380 10 381 644 645 cell_1rw
* cell instance $2472 r0 *1 111.39,10.92
X$2472 382 10 383 644 645 cell_1rw
* cell instance $2473 r0 *1 112.095,10.92
X$2473 384 10 385 644 645 cell_1rw
* cell instance $2474 r0 *1 112.8,10.92
X$2474 386 10 387 644 645 cell_1rw
* cell instance $2475 r0 *1 113.505,10.92
X$2475 388 10 389 644 645 cell_1rw
* cell instance $2476 r0 *1 114.21,10.92
X$2476 390 10 391 644 645 cell_1rw
* cell instance $2477 r0 *1 114.915,10.92
X$2477 392 10 393 644 645 cell_1rw
* cell instance $2478 r0 *1 115.62,10.92
X$2478 394 10 395 644 645 cell_1rw
* cell instance $2479 r0 *1 116.325,10.92
X$2479 396 10 397 644 645 cell_1rw
* cell instance $2480 r0 *1 117.03,10.92
X$2480 398 10 399 644 645 cell_1rw
* cell instance $2481 r0 *1 117.735,10.92
X$2481 400 10 401 644 645 cell_1rw
* cell instance $2482 r0 *1 118.44,10.92
X$2482 402 10 403 644 645 cell_1rw
* cell instance $2483 r0 *1 119.145,10.92
X$2483 404 10 405 644 645 cell_1rw
* cell instance $2484 r0 *1 119.85,10.92
X$2484 406 10 407 644 645 cell_1rw
* cell instance $2485 r0 *1 120.555,10.92
X$2485 408 10 409 644 645 cell_1rw
* cell instance $2486 r0 *1 121.26,10.92
X$2486 410 10 411 644 645 cell_1rw
* cell instance $2487 r0 *1 121.965,10.92
X$2487 412 10 413 644 645 cell_1rw
* cell instance $2488 r0 *1 122.67,10.92
X$2488 414 10 415 644 645 cell_1rw
* cell instance $2489 r0 *1 123.375,10.92
X$2489 416 10 417 644 645 cell_1rw
* cell instance $2490 r0 *1 124.08,10.92
X$2490 418 10 419 644 645 cell_1rw
* cell instance $2491 r0 *1 124.785,10.92
X$2491 420 10 421 644 645 cell_1rw
* cell instance $2492 r0 *1 125.49,10.92
X$2492 422 10 423 644 645 cell_1rw
* cell instance $2493 r0 *1 126.195,10.92
X$2493 424 10 425 644 645 cell_1rw
* cell instance $2494 r0 *1 126.9,10.92
X$2494 426 10 427 644 645 cell_1rw
* cell instance $2495 r0 *1 127.605,10.92
X$2495 428 10 429 644 645 cell_1rw
* cell instance $2496 r0 *1 128.31,10.92
X$2496 430 10 431 644 645 cell_1rw
* cell instance $2497 r0 *1 129.015,10.92
X$2497 432 10 433 644 645 cell_1rw
* cell instance $2498 r0 *1 129.72,10.92
X$2498 434 10 435 644 645 cell_1rw
* cell instance $2499 r0 *1 130.425,10.92
X$2499 436 10 437 644 645 cell_1rw
* cell instance $2500 r0 *1 131.13,10.92
X$2500 438 10 439 644 645 cell_1rw
* cell instance $2501 r0 *1 131.835,10.92
X$2501 440 10 441 644 645 cell_1rw
* cell instance $2502 r0 *1 132.54,10.92
X$2502 442 10 443 644 645 cell_1rw
* cell instance $2503 r0 *1 133.245,10.92
X$2503 444 10 445 644 645 cell_1rw
* cell instance $2504 r0 *1 133.95,10.92
X$2504 446 10 447 644 645 cell_1rw
* cell instance $2505 r0 *1 134.655,10.92
X$2505 448 10 449 644 645 cell_1rw
* cell instance $2506 r0 *1 135.36,10.92
X$2506 450 10 451 644 645 cell_1rw
* cell instance $2507 r0 *1 136.065,10.92
X$2507 452 10 453 644 645 cell_1rw
* cell instance $2508 r0 *1 136.77,10.92
X$2508 454 10 455 644 645 cell_1rw
* cell instance $2509 r0 *1 137.475,10.92
X$2509 456 10 457 644 645 cell_1rw
* cell instance $2510 r0 *1 138.18,10.92
X$2510 458 10 459 644 645 cell_1rw
* cell instance $2511 r0 *1 138.885,10.92
X$2511 460 10 461 644 645 cell_1rw
* cell instance $2512 r0 *1 139.59,10.92
X$2512 462 10 463 644 645 cell_1rw
* cell instance $2513 r0 *1 140.295,10.92
X$2513 464 10 465 644 645 cell_1rw
* cell instance $2514 r0 *1 141,10.92
X$2514 466 10 467 644 645 cell_1rw
* cell instance $2515 r0 *1 141.705,10.92
X$2515 468 10 469 644 645 cell_1rw
* cell instance $2516 r0 *1 142.41,10.92
X$2516 470 10 471 644 645 cell_1rw
* cell instance $2517 r0 *1 143.115,10.92
X$2517 472 10 473 644 645 cell_1rw
* cell instance $2518 r0 *1 143.82,10.92
X$2518 474 10 475 644 645 cell_1rw
* cell instance $2519 r0 *1 144.525,10.92
X$2519 476 10 477 644 645 cell_1rw
* cell instance $2520 r0 *1 145.23,10.92
X$2520 478 10 479 644 645 cell_1rw
* cell instance $2521 r0 *1 145.935,10.92
X$2521 480 10 481 644 645 cell_1rw
* cell instance $2522 r0 *1 146.64,10.92
X$2522 482 10 483 644 645 cell_1rw
* cell instance $2523 r0 *1 147.345,10.92
X$2523 484 10 485 644 645 cell_1rw
* cell instance $2524 r0 *1 148.05,10.92
X$2524 486 10 487 644 645 cell_1rw
* cell instance $2525 r0 *1 148.755,10.92
X$2525 488 10 489 644 645 cell_1rw
* cell instance $2526 r0 *1 149.46,10.92
X$2526 490 10 491 644 645 cell_1rw
* cell instance $2527 r0 *1 150.165,10.92
X$2527 492 10 493 644 645 cell_1rw
* cell instance $2528 r0 *1 150.87,10.92
X$2528 494 10 495 644 645 cell_1rw
* cell instance $2529 r0 *1 151.575,10.92
X$2529 496 10 497 644 645 cell_1rw
* cell instance $2530 r0 *1 152.28,10.92
X$2530 498 10 499 644 645 cell_1rw
* cell instance $2531 r0 *1 152.985,10.92
X$2531 500 10 501 644 645 cell_1rw
* cell instance $2532 r0 *1 153.69,10.92
X$2532 502 10 503 644 645 cell_1rw
* cell instance $2533 r0 *1 154.395,10.92
X$2533 504 10 505 644 645 cell_1rw
* cell instance $2534 r0 *1 155.1,10.92
X$2534 506 10 507 644 645 cell_1rw
* cell instance $2535 r0 *1 155.805,10.92
X$2535 508 10 509 644 645 cell_1rw
* cell instance $2536 r0 *1 156.51,10.92
X$2536 510 10 511 644 645 cell_1rw
* cell instance $2537 r0 *1 157.215,10.92
X$2537 512 10 513 644 645 cell_1rw
* cell instance $2538 r0 *1 157.92,10.92
X$2538 514 10 515 644 645 cell_1rw
* cell instance $2539 r0 *1 158.625,10.92
X$2539 516 10 517 644 645 cell_1rw
* cell instance $2540 r0 *1 159.33,10.92
X$2540 518 10 519 644 645 cell_1rw
* cell instance $2541 r0 *1 160.035,10.92
X$2541 520 10 521 644 645 cell_1rw
* cell instance $2542 r0 *1 160.74,10.92
X$2542 522 10 523 644 645 cell_1rw
* cell instance $2543 r0 *1 161.445,10.92
X$2543 524 10 525 644 645 cell_1rw
* cell instance $2544 r0 *1 162.15,10.92
X$2544 526 10 527 644 645 cell_1rw
* cell instance $2545 r0 *1 162.855,10.92
X$2545 528 10 529 644 645 cell_1rw
* cell instance $2546 r0 *1 163.56,10.92
X$2546 530 10 531 644 645 cell_1rw
* cell instance $2547 r0 *1 164.265,10.92
X$2547 532 10 533 644 645 cell_1rw
* cell instance $2548 r0 *1 164.97,10.92
X$2548 534 10 535 644 645 cell_1rw
* cell instance $2549 r0 *1 165.675,10.92
X$2549 536 10 537 644 645 cell_1rw
* cell instance $2550 r0 *1 166.38,10.92
X$2550 538 10 539 644 645 cell_1rw
* cell instance $2551 r0 *1 167.085,10.92
X$2551 540 10 541 644 645 cell_1rw
* cell instance $2552 r0 *1 167.79,10.92
X$2552 542 10 543 644 645 cell_1rw
* cell instance $2553 r0 *1 168.495,10.92
X$2553 544 10 545 644 645 cell_1rw
* cell instance $2554 r0 *1 169.2,10.92
X$2554 546 10 547 644 645 cell_1rw
* cell instance $2555 r0 *1 169.905,10.92
X$2555 548 10 549 644 645 cell_1rw
* cell instance $2556 r0 *1 170.61,10.92
X$2556 550 10 551 644 645 cell_1rw
* cell instance $2557 r0 *1 171.315,10.92
X$2557 552 10 553 644 645 cell_1rw
* cell instance $2558 r0 *1 172.02,10.92
X$2558 554 10 555 644 645 cell_1rw
* cell instance $2559 r0 *1 172.725,10.92
X$2559 556 10 557 644 645 cell_1rw
* cell instance $2560 r0 *1 173.43,10.92
X$2560 558 10 559 644 645 cell_1rw
* cell instance $2561 r0 *1 174.135,10.92
X$2561 560 10 561 644 645 cell_1rw
* cell instance $2562 r0 *1 174.84,10.92
X$2562 562 10 563 644 645 cell_1rw
* cell instance $2563 r0 *1 175.545,10.92
X$2563 564 10 565 644 645 cell_1rw
* cell instance $2564 r0 *1 176.25,10.92
X$2564 566 10 567 644 645 cell_1rw
* cell instance $2565 r0 *1 176.955,10.92
X$2565 568 10 569 644 645 cell_1rw
* cell instance $2566 r0 *1 177.66,10.92
X$2566 570 10 571 644 645 cell_1rw
* cell instance $2567 r0 *1 178.365,10.92
X$2567 572 10 573 644 645 cell_1rw
* cell instance $2568 r0 *1 179.07,10.92
X$2568 574 10 575 644 645 cell_1rw
* cell instance $2569 r0 *1 179.775,10.92
X$2569 576 10 577 644 645 cell_1rw
* cell instance $2570 r0 *1 180.48,10.92
X$2570 578 10 579 644 645 cell_1rw
* cell instance $2571 r0 *1 0.705,13.65
X$2571 67 11 68 644 645 cell_1rw
* cell instance $2572 r0 *1 0,13.65
X$2572 65 11 66 644 645 cell_1rw
* cell instance $2573 r0 *1 1.41,13.65
X$2573 69 11 70 644 645 cell_1rw
* cell instance $2574 r0 *1 2.115,13.65
X$2574 71 11 72 644 645 cell_1rw
* cell instance $2575 r0 *1 2.82,13.65
X$2575 73 11 74 644 645 cell_1rw
* cell instance $2576 r0 *1 3.525,13.65
X$2576 75 11 76 644 645 cell_1rw
* cell instance $2577 r0 *1 4.23,13.65
X$2577 77 11 78 644 645 cell_1rw
* cell instance $2578 r0 *1 4.935,13.65
X$2578 79 11 80 644 645 cell_1rw
* cell instance $2579 r0 *1 5.64,13.65
X$2579 81 11 82 644 645 cell_1rw
* cell instance $2580 r0 *1 6.345,13.65
X$2580 83 11 84 644 645 cell_1rw
* cell instance $2581 r0 *1 7.05,13.65
X$2581 85 11 86 644 645 cell_1rw
* cell instance $2582 r0 *1 7.755,13.65
X$2582 87 11 88 644 645 cell_1rw
* cell instance $2583 r0 *1 8.46,13.65
X$2583 89 11 90 644 645 cell_1rw
* cell instance $2584 r0 *1 9.165,13.65
X$2584 91 11 92 644 645 cell_1rw
* cell instance $2585 r0 *1 9.87,13.65
X$2585 93 11 94 644 645 cell_1rw
* cell instance $2586 r0 *1 10.575,13.65
X$2586 95 11 96 644 645 cell_1rw
* cell instance $2587 r0 *1 11.28,13.65
X$2587 97 11 98 644 645 cell_1rw
* cell instance $2588 r0 *1 11.985,13.65
X$2588 99 11 100 644 645 cell_1rw
* cell instance $2589 r0 *1 12.69,13.65
X$2589 101 11 102 644 645 cell_1rw
* cell instance $2590 r0 *1 13.395,13.65
X$2590 103 11 104 644 645 cell_1rw
* cell instance $2591 r0 *1 14.1,13.65
X$2591 105 11 106 644 645 cell_1rw
* cell instance $2592 r0 *1 14.805,13.65
X$2592 107 11 108 644 645 cell_1rw
* cell instance $2593 r0 *1 15.51,13.65
X$2593 109 11 110 644 645 cell_1rw
* cell instance $2594 r0 *1 16.215,13.65
X$2594 111 11 112 644 645 cell_1rw
* cell instance $2595 r0 *1 16.92,13.65
X$2595 113 11 114 644 645 cell_1rw
* cell instance $2596 r0 *1 17.625,13.65
X$2596 115 11 116 644 645 cell_1rw
* cell instance $2597 r0 *1 18.33,13.65
X$2597 117 11 118 644 645 cell_1rw
* cell instance $2598 r0 *1 19.035,13.65
X$2598 119 11 120 644 645 cell_1rw
* cell instance $2599 r0 *1 19.74,13.65
X$2599 121 11 122 644 645 cell_1rw
* cell instance $2600 r0 *1 20.445,13.65
X$2600 123 11 124 644 645 cell_1rw
* cell instance $2601 r0 *1 21.15,13.65
X$2601 125 11 126 644 645 cell_1rw
* cell instance $2602 r0 *1 21.855,13.65
X$2602 127 11 128 644 645 cell_1rw
* cell instance $2603 r0 *1 22.56,13.65
X$2603 129 11 130 644 645 cell_1rw
* cell instance $2604 r0 *1 23.265,13.65
X$2604 131 11 132 644 645 cell_1rw
* cell instance $2605 r0 *1 23.97,13.65
X$2605 133 11 134 644 645 cell_1rw
* cell instance $2606 r0 *1 24.675,13.65
X$2606 135 11 136 644 645 cell_1rw
* cell instance $2607 r0 *1 25.38,13.65
X$2607 137 11 138 644 645 cell_1rw
* cell instance $2608 r0 *1 26.085,13.65
X$2608 139 11 140 644 645 cell_1rw
* cell instance $2609 r0 *1 26.79,13.65
X$2609 141 11 142 644 645 cell_1rw
* cell instance $2610 r0 *1 27.495,13.65
X$2610 143 11 144 644 645 cell_1rw
* cell instance $2611 r0 *1 28.2,13.65
X$2611 145 11 146 644 645 cell_1rw
* cell instance $2612 r0 *1 28.905,13.65
X$2612 147 11 148 644 645 cell_1rw
* cell instance $2613 r0 *1 29.61,13.65
X$2613 149 11 150 644 645 cell_1rw
* cell instance $2614 r0 *1 30.315,13.65
X$2614 151 11 152 644 645 cell_1rw
* cell instance $2615 r0 *1 31.02,13.65
X$2615 153 11 154 644 645 cell_1rw
* cell instance $2616 r0 *1 31.725,13.65
X$2616 155 11 156 644 645 cell_1rw
* cell instance $2617 r0 *1 32.43,13.65
X$2617 157 11 158 644 645 cell_1rw
* cell instance $2618 r0 *1 33.135,13.65
X$2618 159 11 160 644 645 cell_1rw
* cell instance $2619 r0 *1 33.84,13.65
X$2619 161 11 162 644 645 cell_1rw
* cell instance $2620 r0 *1 34.545,13.65
X$2620 163 11 164 644 645 cell_1rw
* cell instance $2621 r0 *1 35.25,13.65
X$2621 165 11 166 644 645 cell_1rw
* cell instance $2622 r0 *1 35.955,13.65
X$2622 167 11 168 644 645 cell_1rw
* cell instance $2623 r0 *1 36.66,13.65
X$2623 169 11 170 644 645 cell_1rw
* cell instance $2624 r0 *1 37.365,13.65
X$2624 171 11 172 644 645 cell_1rw
* cell instance $2625 r0 *1 38.07,13.65
X$2625 173 11 174 644 645 cell_1rw
* cell instance $2626 r0 *1 38.775,13.65
X$2626 175 11 176 644 645 cell_1rw
* cell instance $2627 r0 *1 39.48,13.65
X$2627 177 11 178 644 645 cell_1rw
* cell instance $2628 r0 *1 40.185,13.65
X$2628 179 11 180 644 645 cell_1rw
* cell instance $2629 r0 *1 40.89,13.65
X$2629 181 11 182 644 645 cell_1rw
* cell instance $2630 r0 *1 41.595,13.65
X$2630 183 11 184 644 645 cell_1rw
* cell instance $2631 r0 *1 42.3,13.65
X$2631 185 11 186 644 645 cell_1rw
* cell instance $2632 r0 *1 43.005,13.65
X$2632 187 11 188 644 645 cell_1rw
* cell instance $2633 r0 *1 43.71,13.65
X$2633 189 11 190 644 645 cell_1rw
* cell instance $2634 r0 *1 44.415,13.65
X$2634 191 11 192 644 645 cell_1rw
* cell instance $2635 r0 *1 45.12,13.65
X$2635 193 11 194 644 645 cell_1rw
* cell instance $2636 r0 *1 45.825,13.65
X$2636 195 11 196 644 645 cell_1rw
* cell instance $2637 r0 *1 46.53,13.65
X$2637 197 11 198 644 645 cell_1rw
* cell instance $2638 r0 *1 47.235,13.65
X$2638 199 11 200 644 645 cell_1rw
* cell instance $2639 r0 *1 47.94,13.65
X$2639 201 11 202 644 645 cell_1rw
* cell instance $2640 r0 *1 48.645,13.65
X$2640 203 11 204 644 645 cell_1rw
* cell instance $2641 r0 *1 49.35,13.65
X$2641 205 11 206 644 645 cell_1rw
* cell instance $2642 r0 *1 50.055,13.65
X$2642 207 11 208 644 645 cell_1rw
* cell instance $2643 r0 *1 50.76,13.65
X$2643 209 11 210 644 645 cell_1rw
* cell instance $2644 r0 *1 51.465,13.65
X$2644 211 11 212 644 645 cell_1rw
* cell instance $2645 r0 *1 52.17,13.65
X$2645 213 11 214 644 645 cell_1rw
* cell instance $2646 r0 *1 52.875,13.65
X$2646 215 11 216 644 645 cell_1rw
* cell instance $2647 r0 *1 53.58,13.65
X$2647 217 11 218 644 645 cell_1rw
* cell instance $2648 r0 *1 54.285,13.65
X$2648 219 11 220 644 645 cell_1rw
* cell instance $2649 r0 *1 54.99,13.65
X$2649 221 11 222 644 645 cell_1rw
* cell instance $2650 r0 *1 55.695,13.65
X$2650 223 11 224 644 645 cell_1rw
* cell instance $2651 r0 *1 56.4,13.65
X$2651 225 11 226 644 645 cell_1rw
* cell instance $2652 r0 *1 57.105,13.65
X$2652 227 11 228 644 645 cell_1rw
* cell instance $2653 r0 *1 57.81,13.65
X$2653 229 11 230 644 645 cell_1rw
* cell instance $2654 r0 *1 58.515,13.65
X$2654 231 11 232 644 645 cell_1rw
* cell instance $2655 r0 *1 59.22,13.65
X$2655 233 11 234 644 645 cell_1rw
* cell instance $2656 r0 *1 59.925,13.65
X$2656 235 11 236 644 645 cell_1rw
* cell instance $2657 r0 *1 60.63,13.65
X$2657 237 11 238 644 645 cell_1rw
* cell instance $2658 r0 *1 61.335,13.65
X$2658 239 11 240 644 645 cell_1rw
* cell instance $2659 r0 *1 62.04,13.65
X$2659 241 11 242 644 645 cell_1rw
* cell instance $2660 r0 *1 62.745,13.65
X$2660 243 11 244 644 645 cell_1rw
* cell instance $2661 r0 *1 63.45,13.65
X$2661 245 11 246 644 645 cell_1rw
* cell instance $2662 r0 *1 64.155,13.65
X$2662 247 11 248 644 645 cell_1rw
* cell instance $2663 r0 *1 64.86,13.65
X$2663 249 11 250 644 645 cell_1rw
* cell instance $2664 r0 *1 65.565,13.65
X$2664 251 11 252 644 645 cell_1rw
* cell instance $2665 r0 *1 66.27,13.65
X$2665 253 11 254 644 645 cell_1rw
* cell instance $2666 r0 *1 66.975,13.65
X$2666 255 11 256 644 645 cell_1rw
* cell instance $2667 r0 *1 67.68,13.65
X$2667 257 11 258 644 645 cell_1rw
* cell instance $2668 r0 *1 68.385,13.65
X$2668 259 11 260 644 645 cell_1rw
* cell instance $2669 r0 *1 69.09,13.65
X$2669 261 11 262 644 645 cell_1rw
* cell instance $2670 r0 *1 69.795,13.65
X$2670 263 11 264 644 645 cell_1rw
* cell instance $2671 r0 *1 70.5,13.65
X$2671 265 11 266 644 645 cell_1rw
* cell instance $2672 r0 *1 71.205,13.65
X$2672 267 11 268 644 645 cell_1rw
* cell instance $2673 r0 *1 71.91,13.65
X$2673 269 11 270 644 645 cell_1rw
* cell instance $2674 r0 *1 72.615,13.65
X$2674 271 11 272 644 645 cell_1rw
* cell instance $2675 r0 *1 73.32,13.65
X$2675 273 11 274 644 645 cell_1rw
* cell instance $2676 r0 *1 74.025,13.65
X$2676 275 11 276 644 645 cell_1rw
* cell instance $2677 r0 *1 74.73,13.65
X$2677 277 11 278 644 645 cell_1rw
* cell instance $2678 r0 *1 75.435,13.65
X$2678 279 11 280 644 645 cell_1rw
* cell instance $2679 r0 *1 76.14,13.65
X$2679 281 11 282 644 645 cell_1rw
* cell instance $2680 r0 *1 76.845,13.65
X$2680 283 11 284 644 645 cell_1rw
* cell instance $2681 r0 *1 77.55,13.65
X$2681 285 11 286 644 645 cell_1rw
* cell instance $2682 r0 *1 78.255,13.65
X$2682 287 11 288 644 645 cell_1rw
* cell instance $2683 r0 *1 78.96,13.65
X$2683 289 11 290 644 645 cell_1rw
* cell instance $2684 r0 *1 79.665,13.65
X$2684 291 11 292 644 645 cell_1rw
* cell instance $2685 r0 *1 80.37,13.65
X$2685 293 11 294 644 645 cell_1rw
* cell instance $2686 r0 *1 81.075,13.65
X$2686 295 11 296 644 645 cell_1rw
* cell instance $2687 r0 *1 81.78,13.65
X$2687 297 11 298 644 645 cell_1rw
* cell instance $2688 r0 *1 82.485,13.65
X$2688 299 11 300 644 645 cell_1rw
* cell instance $2689 r0 *1 83.19,13.65
X$2689 301 11 302 644 645 cell_1rw
* cell instance $2690 r0 *1 83.895,13.65
X$2690 303 11 304 644 645 cell_1rw
* cell instance $2691 r0 *1 84.6,13.65
X$2691 305 11 306 644 645 cell_1rw
* cell instance $2692 r0 *1 85.305,13.65
X$2692 307 11 308 644 645 cell_1rw
* cell instance $2693 r0 *1 86.01,13.65
X$2693 309 11 310 644 645 cell_1rw
* cell instance $2694 r0 *1 86.715,13.65
X$2694 311 11 312 644 645 cell_1rw
* cell instance $2695 r0 *1 87.42,13.65
X$2695 313 11 314 644 645 cell_1rw
* cell instance $2696 r0 *1 88.125,13.65
X$2696 315 11 316 644 645 cell_1rw
* cell instance $2697 r0 *1 88.83,13.65
X$2697 317 11 318 644 645 cell_1rw
* cell instance $2698 r0 *1 89.535,13.65
X$2698 319 11 320 644 645 cell_1rw
* cell instance $2699 r0 *1 90.24,13.65
X$2699 321 11 323 644 645 cell_1rw
* cell instance $2700 r0 *1 90.945,13.65
X$2700 324 11 325 644 645 cell_1rw
* cell instance $2701 r0 *1 91.65,13.65
X$2701 326 11 327 644 645 cell_1rw
* cell instance $2702 r0 *1 92.355,13.65
X$2702 328 11 329 644 645 cell_1rw
* cell instance $2703 r0 *1 93.06,13.65
X$2703 330 11 331 644 645 cell_1rw
* cell instance $2704 r0 *1 93.765,13.65
X$2704 332 11 333 644 645 cell_1rw
* cell instance $2705 r0 *1 94.47,13.65
X$2705 334 11 335 644 645 cell_1rw
* cell instance $2706 r0 *1 95.175,13.65
X$2706 336 11 337 644 645 cell_1rw
* cell instance $2707 r0 *1 95.88,13.65
X$2707 338 11 339 644 645 cell_1rw
* cell instance $2708 r0 *1 96.585,13.65
X$2708 340 11 341 644 645 cell_1rw
* cell instance $2709 r0 *1 97.29,13.65
X$2709 342 11 343 644 645 cell_1rw
* cell instance $2710 r0 *1 97.995,13.65
X$2710 344 11 345 644 645 cell_1rw
* cell instance $2711 r0 *1 98.7,13.65
X$2711 346 11 347 644 645 cell_1rw
* cell instance $2712 r0 *1 99.405,13.65
X$2712 348 11 349 644 645 cell_1rw
* cell instance $2713 r0 *1 100.11,13.65
X$2713 350 11 351 644 645 cell_1rw
* cell instance $2714 r0 *1 100.815,13.65
X$2714 352 11 353 644 645 cell_1rw
* cell instance $2715 r0 *1 101.52,13.65
X$2715 354 11 355 644 645 cell_1rw
* cell instance $2716 r0 *1 102.225,13.65
X$2716 356 11 357 644 645 cell_1rw
* cell instance $2717 r0 *1 102.93,13.65
X$2717 358 11 359 644 645 cell_1rw
* cell instance $2718 r0 *1 103.635,13.65
X$2718 360 11 361 644 645 cell_1rw
* cell instance $2719 r0 *1 104.34,13.65
X$2719 362 11 363 644 645 cell_1rw
* cell instance $2720 r0 *1 105.045,13.65
X$2720 364 11 365 644 645 cell_1rw
* cell instance $2721 r0 *1 105.75,13.65
X$2721 366 11 367 644 645 cell_1rw
* cell instance $2722 r0 *1 106.455,13.65
X$2722 368 11 369 644 645 cell_1rw
* cell instance $2723 r0 *1 107.16,13.65
X$2723 370 11 371 644 645 cell_1rw
* cell instance $2724 r0 *1 107.865,13.65
X$2724 372 11 373 644 645 cell_1rw
* cell instance $2725 r0 *1 108.57,13.65
X$2725 374 11 375 644 645 cell_1rw
* cell instance $2726 r0 *1 109.275,13.65
X$2726 376 11 377 644 645 cell_1rw
* cell instance $2727 r0 *1 109.98,13.65
X$2727 378 11 379 644 645 cell_1rw
* cell instance $2728 r0 *1 110.685,13.65
X$2728 380 11 381 644 645 cell_1rw
* cell instance $2729 r0 *1 111.39,13.65
X$2729 382 11 383 644 645 cell_1rw
* cell instance $2730 r0 *1 112.095,13.65
X$2730 384 11 385 644 645 cell_1rw
* cell instance $2731 r0 *1 112.8,13.65
X$2731 386 11 387 644 645 cell_1rw
* cell instance $2732 r0 *1 113.505,13.65
X$2732 388 11 389 644 645 cell_1rw
* cell instance $2733 r0 *1 114.21,13.65
X$2733 390 11 391 644 645 cell_1rw
* cell instance $2734 r0 *1 114.915,13.65
X$2734 392 11 393 644 645 cell_1rw
* cell instance $2735 r0 *1 115.62,13.65
X$2735 394 11 395 644 645 cell_1rw
* cell instance $2736 r0 *1 116.325,13.65
X$2736 396 11 397 644 645 cell_1rw
* cell instance $2737 r0 *1 117.03,13.65
X$2737 398 11 399 644 645 cell_1rw
* cell instance $2738 r0 *1 117.735,13.65
X$2738 400 11 401 644 645 cell_1rw
* cell instance $2739 r0 *1 118.44,13.65
X$2739 402 11 403 644 645 cell_1rw
* cell instance $2740 r0 *1 119.145,13.65
X$2740 404 11 405 644 645 cell_1rw
* cell instance $2741 r0 *1 119.85,13.65
X$2741 406 11 407 644 645 cell_1rw
* cell instance $2742 r0 *1 120.555,13.65
X$2742 408 11 409 644 645 cell_1rw
* cell instance $2743 r0 *1 121.26,13.65
X$2743 410 11 411 644 645 cell_1rw
* cell instance $2744 r0 *1 121.965,13.65
X$2744 412 11 413 644 645 cell_1rw
* cell instance $2745 r0 *1 122.67,13.65
X$2745 414 11 415 644 645 cell_1rw
* cell instance $2746 r0 *1 123.375,13.65
X$2746 416 11 417 644 645 cell_1rw
* cell instance $2747 r0 *1 124.08,13.65
X$2747 418 11 419 644 645 cell_1rw
* cell instance $2748 r0 *1 124.785,13.65
X$2748 420 11 421 644 645 cell_1rw
* cell instance $2749 r0 *1 125.49,13.65
X$2749 422 11 423 644 645 cell_1rw
* cell instance $2750 r0 *1 126.195,13.65
X$2750 424 11 425 644 645 cell_1rw
* cell instance $2751 r0 *1 126.9,13.65
X$2751 426 11 427 644 645 cell_1rw
* cell instance $2752 r0 *1 127.605,13.65
X$2752 428 11 429 644 645 cell_1rw
* cell instance $2753 r0 *1 128.31,13.65
X$2753 430 11 431 644 645 cell_1rw
* cell instance $2754 r0 *1 129.015,13.65
X$2754 432 11 433 644 645 cell_1rw
* cell instance $2755 r0 *1 129.72,13.65
X$2755 434 11 435 644 645 cell_1rw
* cell instance $2756 r0 *1 130.425,13.65
X$2756 436 11 437 644 645 cell_1rw
* cell instance $2757 r0 *1 131.13,13.65
X$2757 438 11 439 644 645 cell_1rw
* cell instance $2758 r0 *1 131.835,13.65
X$2758 440 11 441 644 645 cell_1rw
* cell instance $2759 r0 *1 132.54,13.65
X$2759 442 11 443 644 645 cell_1rw
* cell instance $2760 r0 *1 133.245,13.65
X$2760 444 11 445 644 645 cell_1rw
* cell instance $2761 r0 *1 133.95,13.65
X$2761 446 11 447 644 645 cell_1rw
* cell instance $2762 r0 *1 134.655,13.65
X$2762 448 11 449 644 645 cell_1rw
* cell instance $2763 r0 *1 135.36,13.65
X$2763 450 11 451 644 645 cell_1rw
* cell instance $2764 r0 *1 136.065,13.65
X$2764 452 11 453 644 645 cell_1rw
* cell instance $2765 r0 *1 136.77,13.65
X$2765 454 11 455 644 645 cell_1rw
* cell instance $2766 r0 *1 137.475,13.65
X$2766 456 11 457 644 645 cell_1rw
* cell instance $2767 r0 *1 138.18,13.65
X$2767 458 11 459 644 645 cell_1rw
* cell instance $2768 r0 *1 138.885,13.65
X$2768 460 11 461 644 645 cell_1rw
* cell instance $2769 r0 *1 139.59,13.65
X$2769 462 11 463 644 645 cell_1rw
* cell instance $2770 r0 *1 140.295,13.65
X$2770 464 11 465 644 645 cell_1rw
* cell instance $2771 r0 *1 141,13.65
X$2771 466 11 467 644 645 cell_1rw
* cell instance $2772 r0 *1 141.705,13.65
X$2772 468 11 469 644 645 cell_1rw
* cell instance $2773 r0 *1 142.41,13.65
X$2773 470 11 471 644 645 cell_1rw
* cell instance $2774 r0 *1 143.115,13.65
X$2774 472 11 473 644 645 cell_1rw
* cell instance $2775 r0 *1 143.82,13.65
X$2775 474 11 475 644 645 cell_1rw
* cell instance $2776 r0 *1 144.525,13.65
X$2776 476 11 477 644 645 cell_1rw
* cell instance $2777 r0 *1 145.23,13.65
X$2777 478 11 479 644 645 cell_1rw
* cell instance $2778 r0 *1 145.935,13.65
X$2778 480 11 481 644 645 cell_1rw
* cell instance $2779 r0 *1 146.64,13.65
X$2779 482 11 483 644 645 cell_1rw
* cell instance $2780 r0 *1 147.345,13.65
X$2780 484 11 485 644 645 cell_1rw
* cell instance $2781 r0 *1 148.05,13.65
X$2781 486 11 487 644 645 cell_1rw
* cell instance $2782 r0 *1 148.755,13.65
X$2782 488 11 489 644 645 cell_1rw
* cell instance $2783 r0 *1 149.46,13.65
X$2783 490 11 491 644 645 cell_1rw
* cell instance $2784 r0 *1 150.165,13.65
X$2784 492 11 493 644 645 cell_1rw
* cell instance $2785 r0 *1 150.87,13.65
X$2785 494 11 495 644 645 cell_1rw
* cell instance $2786 r0 *1 151.575,13.65
X$2786 496 11 497 644 645 cell_1rw
* cell instance $2787 r0 *1 152.28,13.65
X$2787 498 11 499 644 645 cell_1rw
* cell instance $2788 r0 *1 152.985,13.65
X$2788 500 11 501 644 645 cell_1rw
* cell instance $2789 r0 *1 153.69,13.65
X$2789 502 11 503 644 645 cell_1rw
* cell instance $2790 r0 *1 154.395,13.65
X$2790 504 11 505 644 645 cell_1rw
* cell instance $2791 r0 *1 155.1,13.65
X$2791 506 11 507 644 645 cell_1rw
* cell instance $2792 r0 *1 155.805,13.65
X$2792 508 11 509 644 645 cell_1rw
* cell instance $2793 r0 *1 156.51,13.65
X$2793 510 11 511 644 645 cell_1rw
* cell instance $2794 r0 *1 157.215,13.65
X$2794 512 11 513 644 645 cell_1rw
* cell instance $2795 r0 *1 157.92,13.65
X$2795 514 11 515 644 645 cell_1rw
* cell instance $2796 r0 *1 158.625,13.65
X$2796 516 11 517 644 645 cell_1rw
* cell instance $2797 r0 *1 159.33,13.65
X$2797 518 11 519 644 645 cell_1rw
* cell instance $2798 r0 *1 160.035,13.65
X$2798 520 11 521 644 645 cell_1rw
* cell instance $2799 r0 *1 160.74,13.65
X$2799 522 11 523 644 645 cell_1rw
* cell instance $2800 r0 *1 161.445,13.65
X$2800 524 11 525 644 645 cell_1rw
* cell instance $2801 r0 *1 162.15,13.65
X$2801 526 11 527 644 645 cell_1rw
* cell instance $2802 r0 *1 162.855,13.65
X$2802 528 11 529 644 645 cell_1rw
* cell instance $2803 r0 *1 163.56,13.65
X$2803 530 11 531 644 645 cell_1rw
* cell instance $2804 r0 *1 164.265,13.65
X$2804 532 11 533 644 645 cell_1rw
* cell instance $2805 r0 *1 164.97,13.65
X$2805 534 11 535 644 645 cell_1rw
* cell instance $2806 r0 *1 165.675,13.65
X$2806 536 11 537 644 645 cell_1rw
* cell instance $2807 r0 *1 166.38,13.65
X$2807 538 11 539 644 645 cell_1rw
* cell instance $2808 r0 *1 167.085,13.65
X$2808 540 11 541 644 645 cell_1rw
* cell instance $2809 r0 *1 167.79,13.65
X$2809 542 11 543 644 645 cell_1rw
* cell instance $2810 r0 *1 168.495,13.65
X$2810 544 11 545 644 645 cell_1rw
* cell instance $2811 r0 *1 169.2,13.65
X$2811 546 11 547 644 645 cell_1rw
* cell instance $2812 r0 *1 169.905,13.65
X$2812 548 11 549 644 645 cell_1rw
* cell instance $2813 r0 *1 170.61,13.65
X$2813 550 11 551 644 645 cell_1rw
* cell instance $2814 r0 *1 171.315,13.65
X$2814 552 11 553 644 645 cell_1rw
* cell instance $2815 r0 *1 172.02,13.65
X$2815 554 11 555 644 645 cell_1rw
* cell instance $2816 r0 *1 172.725,13.65
X$2816 556 11 557 644 645 cell_1rw
* cell instance $2817 r0 *1 173.43,13.65
X$2817 558 11 559 644 645 cell_1rw
* cell instance $2818 r0 *1 174.135,13.65
X$2818 560 11 561 644 645 cell_1rw
* cell instance $2819 r0 *1 174.84,13.65
X$2819 562 11 563 644 645 cell_1rw
* cell instance $2820 r0 *1 175.545,13.65
X$2820 564 11 565 644 645 cell_1rw
* cell instance $2821 r0 *1 176.25,13.65
X$2821 566 11 567 644 645 cell_1rw
* cell instance $2822 r0 *1 176.955,13.65
X$2822 568 11 569 644 645 cell_1rw
* cell instance $2823 r0 *1 177.66,13.65
X$2823 570 11 571 644 645 cell_1rw
* cell instance $2824 r0 *1 178.365,13.65
X$2824 572 11 573 644 645 cell_1rw
* cell instance $2825 r0 *1 179.07,13.65
X$2825 574 11 575 644 645 cell_1rw
* cell instance $2826 r0 *1 179.775,13.65
X$2826 576 11 577 644 645 cell_1rw
* cell instance $2827 r0 *1 180.48,13.65
X$2827 578 11 579 644 645 cell_1rw
* cell instance $2828 m0 *1 0.705,16.38
X$2828 67 12 68 644 645 cell_1rw
* cell instance $2829 m0 *1 0,16.38
X$2829 65 12 66 644 645 cell_1rw
* cell instance $2830 m0 *1 1.41,16.38
X$2830 69 12 70 644 645 cell_1rw
* cell instance $2831 m0 *1 2.115,16.38
X$2831 71 12 72 644 645 cell_1rw
* cell instance $2832 m0 *1 2.82,16.38
X$2832 73 12 74 644 645 cell_1rw
* cell instance $2833 m0 *1 3.525,16.38
X$2833 75 12 76 644 645 cell_1rw
* cell instance $2834 m0 *1 4.23,16.38
X$2834 77 12 78 644 645 cell_1rw
* cell instance $2835 m0 *1 4.935,16.38
X$2835 79 12 80 644 645 cell_1rw
* cell instance $2836 m0 *1 5.64,16.38
X$2836 81 12 82 644 645 cell_1rw
* cell instance $2837 m0 *1 6.345,16.38
X$2837 83 12 84 644 645 cell_1rw
* cell instance $2838 m0 *1 7.05,16.38
X$2838 85 12 86 644 645 cell_1rw
* cell instance $2839 m0 *1 7.755,16.38
X$2839 87 12 88 644 645 cell_1rw
* cell instance $2840 m0 *1 8.46,16.38
X$2840 89 12 90 644 645 cell_1rw
* cell instance $2841 m0 *1 9.165,16.38
X$2841 91 12 92 644 645 cell_1rw
* cell instance $2842 m0 *1 9.87,16.38
X$2842 93 12 94 644 645 cell_1rw
* cell instance $2843 m0 *1 10.575,16.38
X$2843 95 12 96 644 645 cell_1rw
* cell instance $2844 m0 *1 11.28,16.38
X$2844 97 12 98 644 645 cell_1rw
* cell instance $2845 m0 *1 11.985,16.38
X$2845 99 12 100 644 645 cell_1rw
* cell instance $2846 m0 *1 12.69,16.38
X$2846 101 12 102 644 645 cell_1rw
* cell instance $2847 m0 *1 13.395,16.38
X$2847 103 12 104 644 645 cell_1rw
* cell instance $2848 m0 *1 14.1,16.38
X$2848 105 12 106 644 645 cell_1rw
* cell instance $2849 m0 *1 14.805,16.38
X$2849 107 12 108 644 645 cell_1rw
* cell instance $2850 m0 *1 15.51,16.38
X$2850 109 12 110 644 645 cell_1rw
* cell instance $2851 m0 *1 16.215,16.38
X$2851 111 12 112 644 645 cell_1rw
* cell instance $2852 m0 *1 16.92,16.38
X$2852 113 12 114 644 645 cell_1rw
* cell instance $2853 m0 *1 17.625,16.38
X$2853 115 12 116 644 645 cell_1rw
* cell instance $2854 m0 *1 18.33,16.38
X$2854 117 12 118 644 645 cell_1rw
* cell instance $2855 m0 *1 19.035,16.38
X$2855 119 12 120 644 645 cell_1rw
* cell instance $2856 m0 *1 19.74,16.38
X$2856 121 12 122 644 645 cell_1rw
* cell instance $2857 m0 *1 20.445,16.38
X$2857 123 12 124 644 645 cell_1rw
* cell instance $2858 m0 *1 21.15,16.38
X$2858 125 12 126 644 645 cell_1rw
* cell instance $2859 m0 *1 21.855,16.38
X$2859 127 12 128 644 645 cell_1rw
* cell instance $2860 m0 *1 22.56,16.38
X$2860 129 12 130 644 645 cell_1rw
* cell instance $2861 m0 *1 23.265,16.38
X$2861 131 12 132 644 645 cell_1rw
* cell instance $2862 m0 *1 23.97,16.38
X$2862 133 12 134 644 645 cell_1rw
* cell instance $2863 m0 *1 24.675,16.38
X$2863 135 12 136 644 645 cell_1rw
* cell instance $2864 m0 *1 25.38,16.38
X$2864 137 12 138 644 645 cell_1rw
* cell instance $2865 m0 *1 26.085,16.38
X$2865 139 12 140 644 645 cell_1rw
* cell instance $2866 m0 *1 26.79,16.38
X$2866 141 12 142 644 645 cell_1rw
* cell instance $2867 m0 *1 27.495,16.38
X$2867 143 12 144 644 645 cell_1rw
* cell instance $2868 m0 *1 28.2,16.38
X$2868 145 12 146 644 645 cell_1rw
* cell instance $2869 m0 *1 28.905,16.38
X$2869 147 12 148 644 645 cell_1rw
* cell instance $2870 m0 *1 29.61,16.38
X$2870 149 12 150 644 645 cell_1rw
* cell instance $2871 m0 *1 30.315,16.38
X$2871 151 12 152 644 645 cell_1rw
* cell instance $2872 m0 *1 31.02,16.38
X$2872 153 12 154 644 645 cell_1rw
* cell instance $2873 m0 *1 31.725,16.38
X$2873 155 12 156 644 645 cell_1rw
* cell instance $2874 m0 *1 32.43,16.38
X$2874 157 12 158 644 645 cell_1rw
* cell instance $2875 m0 *1 33.135,16.38
X$2875 159 12 160 644 645 cell_1rw
* cell instance $2876 m0 *1 33.84,16.38
X$2876 161 12 162 644 645 cell_1rw
* cell instance $2877 m0 *1 34.545,16.38
X$2877 163 12 164 644 645 cell_1rw
* cell instance $2878 m0 *1 35.25,16.38
X$2878 165 12 166 644 645 cell_1rw
* cell instance $2879 m0 *1 35.955,16.38
X$2879 167 12 168 644 645 cell_1rw
* cell instance $2880 m0 *1 36.66,16.38
X$2880 169 12 170 644 645 cell_1rw
* cell instance $2881 m0 *1 37.365,16.38
X$2881 171 12 172 644 645 cell_1rw
* cell instance $2882 m0 *1 38.07,16.38
X$2882 173 12 174 644 645 cell_1rw
* cell instance $2883 m0 *1 38.775,16.38
X$2883 175 12 176 644 645 cell_1rw
* cell instance $2884 m0 *1 39.48,16.38
X$2884 177 12 178 644 645 cell_1rw
* cell instance $2885 m0 *1 40.185,16.38
X$2885 179 12 180 644 645 cell_1rw
* cell instance $2886 m0 *1 40.89,16.38
X$2886 181 12 182 644 645 cell_1rw
* cell instance $2887 m0 *1 41.595,16.38
X$2887 183 12 184 644 645 cell_1rw
* cell instance $2888 m0 *1 42.3,16.38
X$2888 185 12 186 644 645 cell_1rw
* cell instance $2889 m0 *1 43.005,16.38
X$2889 187 12 188 644 645 cell_1rw
* cell instance $2890 m0 *1 43.71,16.38
X$2890 189 12 190 644 645 cell_1rw
* cell instance $2891 m0 *1 44.415,16.38
X$2891 191 12 192 644 645 cell_1rw
* cell instance $2892 m0 *1 45.12,16.38
X$2892 193 12 194 644 645 cell_1rw
* cell instance $2893 m0 *1 45.825,16.38
X$2893 195 12 196 644 645 cell_1rw
* cell instance $2894 m0 *1 46.53,16.38
X$2894 197 12 198 644 645 cell_1rw
* cell instance $2895 m0 *1 47.235,16.38
X$2895 199 12 200 644 645 cell_1rw
* cell instance $2896 m0 *1 47.94,16.38
X$2896 201 12 202 644 645 cell_1rw
* cell instance $2897 m0 *1 48.645,16.38
X$2897 203 12 204 644 645 cell_1rw
* cell instance $2898 m0 *1 49.35,16.38
X$2898 205 12 206 644 645 cell_1rw
* cell instance $2899 m0 *1 50.055,16.38
X$2899 207 12 208 644 645 cell_1rw
* cell instance $2900 m0 *1 50.76,16.38
X$2900 209 12 210 644 645 cell_1rw
* cell instance $2901 m0 *1 51.465,16.38
X$2901 211 12 212 644 645 cell_1rw
* cell instance $2902 m0 *1 52.17,16.38
X$2902 213 12 214 644 645 cell_1rw
* cell instance $2903 m0 *1 52.875,16.38
X$2903 215 12 216 644 645 cell_1rw
* cell instance $2904 m0 *1 53.58,16.38
X$2904 217 12 218 644 645 cell_1rw
* cell instance $2905 m0 *1 54.285,16.38
X$2905 219 12 220 644 645 cell_1rw
* cell instance $2906 m0 *1 54.99,16.38
X$2906 221 12 222 644 645 cell_1rw
* cell instance $2907 m0 *1 55.695,16.38
X$2907 223 12 224 644 645 cell_1rw
* cell instance $2908 m0 *1 56.4,16.38
X$2908 225 12 226 644 645 cell_1rw
* cell instance $2909 m0 *1 57.105,16.38
X$2909 227 12 228 644 645 cell_1rw
* cell instance $2910 m0 *1 57.81,16.38
X$2910 229 12 230 644 645 cell_1rw
* cell instance $2911 m0 *1 58.515,16.38
X$2911 231 12 232 644 645 cell_1rw
* cell instance $2912 m0 *1 59.22,16.38
X$2912 233 12 234 644 645 cell_1rw
* cell instance $2913 m0 *1 59.925,16.38
X$2913 235 12 236 644 645 cell_1rw
* cell instance $2914 m0 *1 60.63,16.38
X$2914 237 12 238 644 645 cell_1rw
* cell instance $2915 m0 *1 61.335,16.38
X$2915 239 12 240 644 645 cell_1rw
* cell instance $2916 m0 *1 62.04,16.38
X$2916 241 12 242 644 645 cell_1rw
* cell instance $2917 m0 *1 62.745,16.38
X$2917 243 12 244 644 645 cell_1rw
* cell instance $2918 m0 *1 63.45,16.38
X$2918 245 12 246 644 645 cell_1rw
* cell instance $2919 m0 *1 64.155,16.38
X$2919 247 12 248 644 645 cell_1rw
* cell instance $2920 m0 *1 64.86,16.38
X$2920 249 12 250 644 645 cell_1rw
* cell instance $2921 m0 *1 65.565,16.38
X$2921 251 12 252 644 645 cell_1rw
* cell instance $2922 m0 *1 66.27,16.38
X$2922 253 12 254 644 645 cell_1rw
* cell instance $2923 m0 *1 66.975,16.38
X$2923 255 12 256 644 645 cell_1rw
* cell instance $2924 m0 *1 67.68,16.38
X$2924 257 12 258 644 645 cell_1rw
* cell instance $2925 m0 *1 68.385,16.38
X$2925 259 12 260 644 645 cell_1rw
* cell instance $2926 m0 *1 69.09,16.38
X$2926 261 12 262 644 645 cell_1rw
* cell instance $2927 m0 *1 69.795,16.38
X$2927 263 12 264 644 645 cell_1rw
* cell instance $2928 m0 *1 70.5,16.38
X$2928 265 12 266 644 645 cell_1rw
* cell instance $2929 m0 *1 71.205,16.38
X$2929 267 12 268 644 645 cell_1rw
* cell instance $2930 m0 *1 71.91,16.38
X$2930 269 12 270 644 645 cell_1rw
* cell instance $2931 m0 *1 72.615,16.38
X$2931 271 12 272 644 645 cell_1rw
* cell instance $2932 m0 *1 73.32,16.38
X$2932 273 12 274 644 645 cell_1rw
* cell instance $2933 m0 *1 74.025,16.38
X$2933 275 12 276 644 645 cell_1rw
* cell instance $2934 m0 *1 74.73,16.38
X$2934 277 12 278 644 645 cell_1rw
* cell instance $2935 m0 *1 75.435,16.38
X$2935 279 12 280 644 645 cell_1rw
* cell instance $2936 m0 *1 76.14,16.38
X$2936 281 12 282 644 645 cell_1rw
* cell instance $2937 m0 *1 76.845,16.38
X$2937 283 12 284 644 645 cell_1rw
* cell instance $2938 m0 *1 77.55,16.38
X$2938 285 12 286 644 645 cell_1rw
* cell instance $2939 m0 *1 78.255,16.38
X$2939 287 12 288 644 645 cell_1rw
* cell instance $2940 m0 *1 78.96,16.38
X$2940 289 12 290 644 645 cell_1rw
* cell instance $2941 m0 *1 79.665,16.38
X$2941 291 12 292 644 645 cell_1rw
* cell instance $2942 m0 *1 80.37,16.38
X$2942 293 12 294 644 645 cell_1rw
* cell instance $2943 m0 *1 81.075,16.38
X$2943 295 12 296 644 645 cell_1rw
* cell instance $2944 m0 *1 81.78,16.38
X$2944 297 12 298 644 645 cell_1rw
* cell instance $2945 m0 *1 82.485,16.38
X$2945 299 12 300 644 645 cell_1rw
* cell instance $2946 m0 *1 83.19,16.38
X$2946 301 12 302 644 645 cell_1rw
* cell instance $2947 m0 *1 83.895,16.38
X$2947 303 12 304 644 645 cell_1rw
* cell instance $2948 m0 *1 84.6,16.38
X$2948 305 12 306 644 645 cell_1rw
* cell instance $2949 m0 *1 85.305,16.38
X$2949 307 12 308 644 645 cell_1rw
* cell instance $2950 m0 *1 86.01,16.38
X$2950 309 12 310 644 645 cell_1rw
* cell instance $2951 m0 *1 86.715,16.38
X$2951 311 12 312 644 645 cell_1rw
* cell instance $2952 m0 *1 87.42,16.38
X$2952 313 12 314 644 645 cell_1rw
* cell instance $2953 m0 *1 88.125,16.38
X$2953 315 12 316 644 645 cell_1rw
* cell instance $2954 m0 *1 88.83,16.38
X$2954 317 12 318 644 645 cell_1rw
* cell instance $2955 m0 *1 89.535,16.38
X$2955 319 12 320 644 645 cell_1rw
* cell instance $2956 m0 *1 90.24,16.38
X$2956 321 12 323 644 645 cell_1rw
* cell instance $2957 m0 *1 90.945,16.38
X$2957 324 12 325 644 645 cell_1rw
* cell instance $2958 m0 *1 91.65,16.38
X$2958 326 12 327 644 645 cell_1rw
* cell instance $2959 m0 *1 92.355,16.38
X$2959 328 12 329 644 645 cell_1rw
* cell instance $2960 m0 *1 93.06,16.38
X$2960 330 12 331 644 645 cell_1rw
* cell instance $2961 m0 *1 93.765,16.38
X$2961 332 12 333 644 645 cell_1rw
* cell instance $2962 m0 *1 94.47,16.38
X$2962 334 12 335 644 645 cell_1rw
* cell instance $2963 m0 *1 95.175,16.38
X$2963 336 12 337 644 645 cell_1rw
* cell instance $2964 m0 *1 95.88,16.38
X$2964 338 12 339 644 645 cell_1rw
* cell instance $2965 m0 *1 96.585,16.38
X$2965 340 12 341 644 645 cell_1rw
* cell instance $2966 m0 *1 97.29,16.38
X$2966 342 12 343 644 645 cell_1rw
* cell instance $2967 m0 *1 97.995,16.38
X$2967 344 12 345 644 645 cell_1rw
* cell instance $2968 m0 *1 98.7,16.38
X$2968 346 12 347 644 645 cell_1rw
* cell instance $2969 m0 *1 99.405,16.38
X$2969 348 12 349 644 645 cell_1rw
* cell instance $2970 m0 *1 100.11,16.38
X$2970 350 12 351 644 645 cell_1rw
* cell instance $2971 m0 *1 100.815,16.38
X$2971 352 12 353 644 645 cell_1rw
* cell instance $2972 m0 *1 101.52,16.38
X$2972 354 12 355 644 645 cell_1rw
* cell instance $2973 m0 *1 102.225,16.38
X$2973 356 12 357 644 645 cell_1rw
* cell instance $2974 m0 *1 102.93,16.38
X$2974 358 12 359 644 645 cell_1rw
* cell instance $2975 m0 *1 103.635,16.38
X$2975 360 12 361 644 645 cell_1rw
* cell instance $2976 m0 *1 104.34,16.38
X$2976 362 12 363 644 645 cell_1rw
* cell instance $2977 m0 *1 105.045,16.38
X$2977 364 12 365 644 645 cell_1rw
* cell instance $2978 m0 *1 105.75,16.38
X$2978 366 12 367 644 645 cell_1rw
* cell instance $2979 m0 *1 106.455,16.38
X$2979 368 12 369 644 645 cell_1rw
* cell instance $2980 m0 *1 107.16,16.38
X$2980 370 12 371 644 645 cell_1rw
* cell instance $2981 m0 *1 107.865,16.38
X$2981 372 12 373 644 645 cell_1rw
* cell instance $2982 m0 *1 108.57,16.38
X$2982 374 12 375 644 645 cell_1rw
* cell instance $2983 m0 *1 109.275,16.38
X$2983 376 12 377 644 645 cell_1rw
* cell instance $2984 m0 *1 109.98,16.38
X$2984 378 12 379 644 645 cell_1rw
* cell instance $2985 m0 *1 110.685,16.38
X$2985 380 12 381 644 645 cell_1rw
* cell instance $2986 m0 *1 111.39,16.38
X$2986 382 12 383 644 645 cell_1rw
* cell instance $2987 m0 *1 112.095,16.38
X$2987 384 12 385 644 645 cell_1rw
* cell instance $2988 m0 *1 112.8,16.38
X$2988 386 12 387 644 645 cell_1rw
* cell instance $2989 m0 *1 113.505,16.38
X$2989 388 12 389 644 645 cell_1rw
* cell instance $2990 m0 *1 114.21,16.38
X$2990 390 12 391 644 645 cell_1rw
* cell instance $2991 m0 *1 114.915,16.38
X$2991 392 12 393 644 645 cell_1rw
* cell instance $2992 m0 *1 115.62,16.38
X$2992 394 12 395 644 645 cell_1rw
* cell instance $2993 m0 *1 116.325,16.38
X$2993 396 12 397 644 645 cell_1rw
* cell instance $2994 m0 *1 117.03,16.38
X$2994 398 12 399 644 645 cell_1rw
* cell instance $2995 m0 *1 117.735,16.38
X$2995 400 12 401 644 645 cell_1rw
* cell instance $2996 m0 *1 118.44,16.38
X$2996 402 12 403 644 645 cell_1rw
* cell instance $2997 m0 *1 119.145,16.38
X$2997 404 12 405 644 645 cell_1rw
* cell instance $2998 m0 *1 119.85,16.38
X$2998 406 12 407 644 645 cell_1rw
* cell instance $2999 m0 *1 120.555,16.38
X$2999 408 12 409 644 645 cell_1rw
* cell instance $3000 m0 *1 121.26,16.38
X$3000 410 12 411 644 645 cell_1rw
* cell instance $3001 m0 *1 121.965,16.38
X$3001 412 12 413 644 645 cell_1rw
* cell instance $3002 m0 *1 122.67,16.38
X$3002 414 12 415 644 645 cell_1rw
* cell instance $3003 m0 *1 123.375,16.38
X$3003 416 12 417 644 645 cell_1rw
* cell instance $3004 m0 *1 124.08,16.38
X$3004 418 12 419 644 645 cell_1rw
* cell instance $3005 m0 *1 124.785,16.38
X$3005 420 12 421 644 645 cell_1rw
* cell instance $3006 m0 *1 125.49,16.38
X$3006 422 12 423 644 645 cell_1rw
* cell instance $3007 m0 *1 126.195,16.38
X$3007 424 12 425 644 645 cell_1rw
* cell instance $3008 m0 *1 126.9,16.38
X$3008 426 12 427 644 645 cell_1rw
* cell instance $3009 m0 *1 127.605,16.38
X$3009 428 12 429 644 645 cell_1rw
* cell instance $3010 m0 *1 128.31,16.38
X$3010 430 12 431 644 645 cell_1rw
* cell instance $3011 m0 *1 129.015,16.38
X$3011 432 12 433 644 645 cell_1rw
* cell instance $3012 m0 *1 129.72,16.38
X$3012 434 12 435 644 645 cell_1rw
* cell instance $3013 m0 *1 130.425,16.38
X$3013 436 12 437 644 645 cell_1rw
* cell instance $3014 m0 *1 131.13,16.38
X$3014 438 12 439 644 645 cell_1rw
* cell instance $3015 m0 *1 131.835,16.38
X$3015 440 12 441 644 645 cell_1rw
* cell instance $3016 m0 *1 132.54,16.38
X$3016 442 12 443 644 645 cell_1rw
* cell instance $3017 m0 *1 133.245,16.38
X$3017 444 12 445 644 645 cell_1rw
* cell instance $3018 m0 *1 133.95,16.38
X$3018 446 12 447 644 645 cell_1rw
* cell instance $3019 m0 *1 134.655,16.38
X$3019 448 12 449 644 645 cell_1rw
* cell instance $3020 m0 *1 135.36,16.38
X$3020 450 12 451 644 645 cell_1rw
* cell instance $3021 m0 *1 136.065,16.38
X$3021 452 12 453 644 645 cell_1rw
* cell instance $3022 m0 *1 136.77,16.38
X$3022 454 12 455 644 645 cell_1rw
* cell instance $3023 m0 *1 137.475,16.38
X$3023 456 12 457 644 645 cell_1rw
* cell instance $3024 m0 *1 138.18,16.38
X$3024 458 12 459 644 645 cell_1rw
* cell instance $3025 m0 *1 138.885,16.38
X$3025 460 12 461 644 645 cell_1rw
* cell instance $3026 m0 *1 139.59,16.38
X$3026 462 12 463 644 645 cell_1rw
* cell instance $3027 m0 *1 140.295,16.38
X$3027 464 12 465 644 645 cell_1rw
* cell instance $3028 m0 *1 141,16.38
X$3028 466 12 467 644 645 cell_1rw
* cell instance $3029 m0 *1 141.705,16.38
X$3029 468 12 469 644 645 cell_1rw
* cell instance $3030 m0 *1 142.41,16.38
X$3030 470 12 471 644 645 cell_1rw
* cell instance $3031 m0 *1 143.115,16.38
X$3031 472 12 473 644 645 cell_1rw
* cell instance $3032 m0 *1 143.82,16.38
X$3032 474 12 475 644 645 cell_1rw
* cell instance $3033 m0 *1 144.525,16.38
X$3033 476 12 477 644 645 cell_1rw
* cell instance $3034 m0 *1 145.23,16.38
X$3034 478 12 479 644 645 cell_1rw
* cell instance $3035 m0 *1 145.935,16.38
X$3035 480 12 481 644 645 cell_1rw
* cell instance $3036 m0 *1 146.64,16.38
X$3036 482 12 483 644 645 cell_1rw
* cell instance $3037 m0 *1 147.345,16.38
X$3037 484 12 485 644 645 cell_1rw
* cell instance $3038 m0 *1 148.05,16.38
X$3038 486 12 487 644 645 cell_1rw
* cell instance $3039 m0 *1 148.755,16.38
X$3039 488 12 489 644 645 cell_1rw
* cell instance $3040 m0 *1 149.46,16.38
X$3040 490 12 491 644 645 cell_1rw
* cell instance $3041 m0 *1 150.165,16.38
X$3041 492 12 493 644 645 cell_1rw
* cell instance $3042 m0 *1 150.87,16.38
X$3042 494 12 495 644 645 cell_1rw
* cell instance $3043 m0 *1 151.575,16.38
X$3043 496 12 497 644 645 cell_1rw
* cell instance $3044 m0 *1 152.28,16.38
X$3044 498 12 499 644 645 cell_1rw
* cell instance $3045 m0 *1 152.985,16.38
X$3045 500 12 501 644 645 cell_1rw
* cell instance $3046 m0 *1 153.69,16.38
X$3046 502 12 503 644 645 cell_1rw
* cell instance $3047 m0 *1 154.395,16.38
X$3047 504 12 505 644 645 cell_1rw
* cell instance $3048 m0 *1 155.1,16.38
X$3048 506 12 507 644 645 cell_1rw
* cell instance $3049 m0 *1 155.805,16.38
X$3049 508 12 509 644 645 cell_1rw
* cell instance $3050 m0 *1 156.51,16.38
X$3050 510 12 511 644 645 cell_1rw
* cell instance $3051 m0 *1 157.215,16.38
X$3051 512 12 513 644 645 cell_1rw
* cell instance $3052 m0 *1 157.92,16.38
X$3052 514 12 515 644 645 cell_1rw
* cell instance $3053 m0 *1 158.625,16.38
X$3053 516 12 517 644 645 cell_1rw
* cell instance $3054 m0 *1 159.33,16.38
X$3054 518 12 519 644 645 cell_1rw
* cell instance $3055 m0 *1 160.035,16.38
X$3055 520 12 521 644 645 cell_1rw
* cell instance $3056 m0 *1 160.74,16.38
X$3056 522 12 523 644 645 cell_1rw
* cell instance $3057 m0 *1 161.445,16.38
X$3057 524 12 525 644 645 cell_1rw
* cell instance $3058 m0 *1 162.15,16.38
X$3058 526 12 527 644 645 cell_1rw
* cell instance $3059 m0 *1 162.855,16.38
X$3059 528 12 529 644 645 cell_1rw
* cell instance $3060 m0 *1 163.56,16.38
X$3060 530 12 531 644 645 cell_1rw
* cell instance $3061 m0 *1 164.265,16.38
X$3061 532 12 533 644 645 cell_1rw
* cell instance $3062 m0 *1 164.97,16.38
X$3062 534 12 535 644 645 cell_1rw
* cell instance $3063 m0 *1 165.675,16.38
X$3063 536 12 537 644 645 cell_1rw
* cell instance $3064 m0 *1 166.38,16.38
X$3064 538 12 539 644 645 cell_1rw
* cell instance $3065 m0 *1 167.085,16.38
X$3065 540 12 541 644 645 cell_1rw
* cell instance $3066 m0 *1 167.79,16.38
X$3066 542 12 543 644 645 cell_1rw
* cell instance $3067 m0 *1 168.495,16.38
X$3067 544 12 545 644 645 cell_1rw
* cell instance $3068 m0 *1 169.2,16.38
X$3068 546 12 547 644 645 cell_1rw
* cell instance $3069 m0 *1 169.905,16.38
X$3069 548 12 549 644 645 cell_1rw
* cell instance $3070 m0 *1 170.61,16.38
X$3070 550 12 551 644 645 cell_1rw
* cell instance $3071 m0 *1 171.315,16.38
X$3071 552 12 553 644 645 cell_1rw
* cell instance $3072 m0 *1 172.02,16.38
X$3072 554 12 555 644 645 cell_1rw
* cell instance $3073 m0 *1 172.725,16.38
X$3073 556 12 557 644 645 cell_1rw
* cell instance $3074 m0 *1 173.43,16.38
X$3074 558 12 559 644 645 cell_1rw
* cell instance $3075 m0 *1 174.135,16.38
X$3075 560 12 561 644 645 cell_1rw
* cell instance $3076 m0 *1 174.84,16.38
X$3076 562 12 563 644 645 cell_1rw
* cell instance $3077 m0 *1 175.545,16.38
X$3077 564 12 565 644 645 cell_1rw
* cell instance $3078 m0 *1 176.25,16.38
X$3078 566 12 567 644 645 cell_1rw
* cell instance $3079 m0 *1 176.955,16.38
X$3079 568 12 569 644 645 cell_1rw
* cell instance $3080 m0 *1 177.66,16.38
X$3080 570 12 571 644 645 cell_1rw
* cell instance $3081 m0 *1 178.365,16.38
X$3081 572 12 573 644 645 cell_1rw
* cell instance $3082 m0 *1 179.07,16.38
X$3082 574 12 575 644 645 cell_1rw
* cell instance $3083 m0 *1 179.775,16.38
X$3083 576 12 577 644 645 cell_1rw
* cell instance $3084 m0 *1 180.48,16.38
X$3084 578 12 579 644 645 cell_1rw
* cell instance $3085 r0 *1 0.705,16.38
X$3085 67 13 68 644 645 cell_1rw
* cell instance $3086 r0 *1 0,16.38
X$3086 65 13 66 644 645 cell_1rw
* cell instance $3087 r0 *1 1.41,16.38
X$3087 69 13 70 644 645 cell_1rw
* cell instance $3088 r0 *1 2.115,16.38
X$3088 71 13 72 644 645 cell_1rw
* cell instance $3089 r0 *1 2.82,16.38
X$3089 73 13 74 644 645 cell_1rw
* cell instance $3090 r0 *1 3.525,16.38
X$3090 75 13 76 644 645 cell_1rw
* cell instance $3091 r0 *1 4.23,16.38
X$3091 77 13 78 644 645 cell_1rw
* cell instance $3092 r0 *1 4.935,16.38
X$3092 79 13 80 644 645 cell_1rw
* cell instance $3093 r0 *1 5.64,16.38
X$3093 81 13 82 644 645 cell_1rw
* cell instance $3094 r0 *1 6.345,16.38
X$3094 83 13 84 644 645 cell_1rw
* cell instance $3095 r0 *1 7.05,16.38
X$3095 85 13 86 644 645 cell_1rw
* cell instance $3096 r0 *1 7.755,16.38
X$3096 87 13 88 644 645 cell_1rw
* cell instance $3097 r0 *1 8.46,16.38
X$3097 89 13 90 644 645 cell_1rw
* cell instance $3098 r0 *1 9.165,16.38
X$3098 91 13 92 644 645 cell_1rw
* cell instance $3099 r0 *1 9.87,16.38
X$3099 93 13 94 644 645 cell_1rw
* cell instance $3100 r0 *1 10.575,16.38
X$3100 95 13 96 644 645 cell_1rw
* cell instance $3101 r0 *1 11.28,16.38
X$3101 97 13 98 644 645 cell_1rw
* cell instance $3102 r0 *1 11.985,16.38
X$3102 99 13 100 644 645 cell_1rw
* cell instance $3103 r0 *1 12.69,16.38
X$3103 101 13 102 644 645 cell_1rw
* cell instance $3104 r0 *1 13.395,16.38
X$3104 103 13 104 644 645 cell_1rw
* cell instance $3105 r0 *1 14.1,16.38
X$3105 105 13 106 644 645 cell_1rw
* cell instance $3106 r0 *1 14.805,16.38
X$3106 107 13 108 644 645 cell_1rw
* cell instance $3107 r0 *1 15.51,16.38
X$3107 109 13 110 644 645 cell_1rw
* cell instance $3108 r0 *1 16.215,16.38
X$3108 111 13 112 644 645 cell_1rw
* cell instance $3109 r0 *1 16.92,16.38
X$3109 113 13 114 644 645 cell_1rw
* cell instance $3110 r0 *1 17.625,16.38
X$3110 115 13 116 644 645 cell_1rw
* cell instance $3111 r0 *1 18.33,16.38
X$3111 117 13 118 644 645 cell_1rw
* cell instance $3112 r0 *1 19.035,16.38
X$3112 119 13 120 644 645 cell_1rw
* cell instance $3113 r0 *1 19.74,16.38
X$3113 121 13 122 644 645 cell_1rw
* cell instance $3114 r0 *1 20.445,16.38
X$3114 123 13 124 644 645 cell_1rw
* cell instance $3115 r0 *1 21.15,16.38
X$3115 125 13 126 644 645 cell_1rw
* cell instance $3116 r0 *1 21.855,16.38
X$3116 127 13 128 644 645 cell_1rw
* cell instance $3117 r0 *1 22.56,16.38
X$3117 129 13 130 644 645 cell_1rw
* cell instance $3118 r0 *1 23.265,16.38
X$3118 131 13 132 644 645 cell_1rw
* cell instance $3119 r0 *1 23.97,16.38
X$3119 133 13 134 644 645 cell_1rw
* cell instance $3120 r0 *1 24.675,16.38
X$3120 135 13 136 644 645 cell_1rw
* cell instance $3121 r0 *1 25.38,16.38
X$3121 137 13 138 644 645 cell_1rw
* cell instance $3122 r0 *1 26.085,16.38
X$3122 139 13 140 644 645 cell_1rw
* cell instance $3123 r0 *1 26.79,16.38
X$3123 141 13 142 644 645 cell_1rw
* cell instance $3124 r0 *1 27.495,16.38
X$3124 143 13 144 644 645 cell_1rw
* cell instance $3125 r0 *1 28.2,16.38
X$3125 145 13 146 644 645 cell_1rw
* cell instance $3126 r0 *1 28.905,16.38
X$3126 147 13 148 644 645 cell_1rw
* cell instance $3127 r0 *1 29.61,16.38
X$3127 149 13 150 644 645 cell_1rw
* cell instance $3128 r0 *1 30.315,16.38
X$3128 151 13 152 644 645 cell_1rw
* cell instance $3129 r0 *1 31.02,16.38
X$3129 153 13 154 644 645 cell_1rw
* cell instance $3130 r0 *1 31.725,16.38
X$3130 155 13 156 644 645 cell_1rw
* cell instance $3131 r0 *1 32.43,16.38
X$3131 157 13 158 644 645 cell_1rw
* cell instance $3132 r0 *1 33.135,16.38
X$3132 159 13 160 644 645 cell_1rw
* cell instance $3133 r0 *1 33.84,16.38
X$3133 161 13 162 644 645 cell_1rw
* cell instance $3134 r0 *1 34.545,16.38
X$3134 163 13 164 644 645 cell_1rw
* cell instance $3135 r0 *1 35.25,16.38
X$3135 165 13 166 644 645 cell_1rw
* cell instance $3136 r0 *1 35.955,16.38
X$3136 167 13 168 644 645 cell_1rw
* cell instance $3137 r0 *1 36.66,16.38
X$3137 169 13 170 644 645 cell_1rw
* cell instance $3138 r0 *1 37.365,16.38
X$3138 171 13 172 644 645 cell_1rw
* cell instance $3139 r0 *1 38.07,16.38
X$3139 173 13 174 644 645 cell_1rw
* cell instance $3140 r0 *1 38.775,16.38
X$3140 175 13 176 644 645 cell_1rw
* cell instance $3141 r0 *1 39.48,16.38
X$3141 177 13 178 644 645 cell_1rw
* cell instance $3142 r0 *1 40.185,16.38
X$3142 179 13 180 644 645 cell_1rw
* cell instance $3143 r0 *1 40.89,16.38
X$3143 181 13 182 644 645 cell_1rw
* cell instance $3144 r0 *1 41.595,16.38
X$3144 183 13 184 644 645 cell_1rw
* cell instance $3145 r0 *1 42.3,16.38
X$3145 185 13 186 644 645 cell_1rw
* cell instance $3146 r0 *1 43.005,16.38
X$3146 187 13 188 644 645 cell_1rw
* cell instance $3147 r0 *1 43.71,16.38
X$3147 189 13 190 644 645 cell_1rw
* cell instance $3148 r0 *1 44.415,16.38
X$3148 191 13 192 644 645 cell_1rw
* cell instance $3149 r0 *1 45.12,16.38
X$3149 193 13 194 644 645 cell_1rw
* cell instance $3150 r0 *1 45.825,16.38
X$3150 195 13 196 644 645 cell_1rw
* cell instance $3151 r0 *1 46.53,16.38
X$3151 197 13 198 644 645 cell_1rw
* cell instance $3152 r0 *1 47.235,16.38
X$3152 199 13 200 644 645 cell_1rw
* cell instance $3153 r0 *1 47.94,16.38
X$3153 201 13 202 644 645 cell_1rw
* cell instance $3154 r0 *1 48.645,16.38
X$3154 203 13 204 644 645 cell_1rw
* cell instance $3155 r0 *1 49.35,16.38
X$3155 205 13 206 644 645 cell_1rw
* cell instance $3156 r0 *1 50.055,16.38
X$3156 207 13 208 644 645 cell_1rw
* cell instance $3157 r0 *1 50.76,16.38
X$3157 209 13 210 644 645 cell_1rw
* cell instance $3158 r0 *1 51.465,16.38
X$3158 211 13 212 644 645 cell_1rw
* cell instance $3159 r0 *1 52.17,16.38
X$3159 213 13 214 644 645 cell_1rw
* cell instance $3160 r0 *1 52.875,16.38
X$3160 215 13 216 644 645 cell_1rw
* cell instance $3161 r0 *1 53.58,16.38
X$3161 217 13 218 644 645 cell_1rw
* cell instance $3162 r0 *1 54.285,16.38
X$3162 219 13 220 644 645 cell_1rw
* cell instance $3163 r0 *1 54.99,16.38
X$3163 221 13 222 644 645 cell_1rw
* cell instance $3164 r0 *1 55.695,16.38
X$3164 223 13 224 644 645 cell_1rw
* cell instance $3165 r0 *1 56.4,16.38
X$3165 225 13 226 644 645 cell_1rw
* cell instance $3166 r0 *1 57.105,16.38
X$3166 227 13 228 644 645 cell_1rw
* cell instance $3167 r0 *1 57.81,16.38
X$3167 229 13 230 644 645 cell_1rw
* cell instance $3168 r0 *1 58.515,16.38
X$3168 231 13 232 644 645 cell_1rw
* cell instance $3169 r0 *1 59.22,16.38
X$3169 233 13 234 644 645 cell_1rw
* cell instance $3170 r0 *1 59.925,16.38
X$3170 235 13 236 644 645 cell_1rw
* cell instance $3171 r0 *1 60.63,16.38
X$3171 237 13 238 644 645 cell_1rw
* cell instance $3172 r0 *1 61.335,16.38
X$3172 239 13 240 644 645 cell_1rw
* cell instance $3173 r0 *1 62.04,16.38
X$3173 241 13 242 644 645 cell_1rw
* cell instance $3174 r0 *1 62.745,16.38
X$3174 243 13 244 644 645 cell_1rw
* cell instance $3175 r0 *1 63.45,16.38
X$3175 245 13 246 644 645 cell_1rw
* cell instance $3176 r0 *1 64.155,16.38
X$3176 247 13 248 644 645 cell_1rw
* cell instance $3177 r0 *1 64.86,16.38
X$3177 249 13 250 644 645 cell_1rw
* cell instance $3178 r0 *1 65.565,16.38
X$3178 251 13 252 644 645 cell_1rw
* cell instance $3179 r0 *1 66.27,16.38
X$3179 253 13 254 644 645 cell_1rw
* cell instance $3180 r0 *1 66.975,16.38
X$3180 255 13 256 644 645 cell_1rw
* cell instance $3181 r0 *1 67.68,16.38
X$3181 257 13 258 644 645 cell_1rw
* cell instance $3182 r0 *1 68.385,16.38
X$3182 259 13 260 644 645 cell_1rw
* cell instance $3183 r0 *1 69.09,16.38
X$3183 261 13 262 644 645 cell_1rw
* cell instance $3184 r0 *1 69.795,16.38
X$3184 263 13 264 644 645 cell_1rw
* cell instance $3185 r0 *1 70.5,16.38
X$3185 265 13 266 644 645 cell_1rw
* cell instance $3186 r0 *1 71.205,16.38
X$3186 267 13 268 644 645 cell_1rw
* cell instance $3187 r0 *1 71.91,16.38
X$3187 269 13 270 644 645 cell_1rw
* cell instance $3188 r0 *1 72.615,16.38
X$3188 271 13 272 644 645 cell_1rw
* cell instance $3189 r0 *1 73.32,16.38
X$3189 273 13 274 644 645 cell_1rw
* cell instance $3190 r0 *1 74.025,16.38
X$3190 275 13 276 644 645 cell_1rw
* cell instance $3191 r0 *1 74.73,16.38
X$3191 277 13 278 644 645 cell_1rw
* cell instance $3192 r0 *1 75.435,16.38
X$3192 279 13 280 644 645 cell_1rw
* cell instance $3193 r0 *1 76.14,16.38
X$3193 281 13 282 644 645 cell_1rw
* cell instance $3194 r0 *1 76.845,16.38
X$3194 283 13 284 644 645 cell_1rw
* cell instance $3195 r0 *1 77.55,16.38
X$3195 285 13 286 644 645 cell_1rw
* cell instance $3196 r0 *1 78.255,16.38
X$3196 287 13 288 644 645 cell_1rw
* cell instance $3197 r0 *1 78.96,16.38
X$3197 289 13 290 644 645 cell_1rw
* cell instance $3198 r0 *1 79.665,16.38
X$3198 291 13 292 644 645 cell_1rw
* cell instance $3199 r0 *1 80.37,16.38
X$3199 293 13 294 644 645 cell_1rw
* cell instance $3200 r0 *1 81.075,16.38
X$3200 295 13 296 644 645 cell_1rw
* cell instance $3201 r0 *1 81.78,16.38
X$3201 297 13 298 644 645 cell_1rw
* cell instance $3202 r0 *1 82.485,16.38
X$3202 299 13 300 644 645 cell_1rw
* cell instance $3203 r0 *1 83.19,16.38
X$3203 301 13 302 644 645 cell_1rw
* cell instance $3204 r0 *1 83.895,16.38
X$3204 303 13 304 644 645 cell_1rw
* cell instance $3205 r0 *1 84.6,16.38
X$3205 305 13 306 644 645 cell_1rw
* cell instance $3206 r0 *1 85.305,16.38
X$3206 307 13 308 644 645 cell_1rw
* cell instance $3207 r0 *1 86.01,16.38
X$3207 309 13 310 644 645 cell_1rw
* cell instance $3208 r0 *1 86.715,16.38
X$3208 311 13 312 644 645 cell_1rw
* cell instance $3209 r0 *1 87.42,16.38
X$3209 313 13 314 644 645 cell_1rw
* cell instance $3210 r0 *1 88.125,16.38
X$3210 315 13 316 644 645 cell_1rw
* cell instance $3211 r0 *1 88.83,16.38
X$3211 317 13 318 644 645 cell_1rw
* cell instance $3212 r0 *1 89.535,16.38
X$3212 319 13 320 644 645 cell_1rw
* cell instance $3213 r0 *1 90.24,16.38
X$3213 321 13 323 644 645 cell_1rw
* cell instance $3214 r0 *1 90.945,16.38
X$3214 324 13 325 644 645 cell_1rw
* cell instance $3215 r0 *1 91.65,16.38
X$3215 326 13 327 644 645 cell_1rw
* cell instance $3216 r0 *1 92.355,16.38
X$3216 328 13 329 644 645 cell_1rw
* cell instance $3217 r0 *1 93.06,16.38
X$3217 330 13 331 644 645 cell_1rw
* cell instance $3218 r0 *1 93.765,16.38
X$3218 332 13 333 644 645 cell_1rw
* cell instance $3219 r0 *1 94.47,16.38
X$3219 334 13 335 644 645 cell_1rw
* cell instance $3220 r0 *1 95.175,16.38
X$3220 336 13 337 644 645 cell_1rw
* cell instance $3221 r0 *1 95.88,16.38
X$3221 338 13 339 644 645 cell_1rw
* cell instance $3222 r0 *1 96.585,16.38
X$3222 340 13 341 644 645 cell_1rw
* cell instance $3223 r0 *1 97.29,16.38
X$3223 342 13 343 644 645 cell_1rw
* cell instance $3224 r0 *1 97.995,16.38
X$3224 344 13 345 644 645 cell_1rw
* cell instance $3225 r0 *1 98.7,16.38
X$3225 346 13 347 644 645 cell_1rw
* cell instance $3226 r0 *1 99.405,16.38
X$3226 348 13 349 644 645 cell_1rw
* cell instance $3227 r0 *1 100.11,16.38
X$3227 350 13 351 644 645 cell_1rw
* cell instance $3228 r0 *1 100.815,16.38
X$3228 352 13 353 644 645 cell_1rw
* cell instance $3229 r0 *1 101.52,16.38
X$3229 354 13 355 644 645 cell_1rw
* cell instance $3230 r0 *1 102.225,16.38
X$3230 356 13 357 644 645 cell_1rw
* cell instance $3231 r0 *1 102.93,16.38
X$3231 358 13 359 644 645 cell_1rw
* cell instance $3232 r0 *1 103.635,16.38
X$3232 360 13 361 644 645 cell_1rw
* cell instance $3233 r0 *1 104.34,16.38
X$3233 362 13 363 644 645 cell_1rw
* cell instance $3234 r0 *1 105.045,16.38
X$3234 364 13 365 644 645 cell_1rw
* cell instance $3235 r0 *1 105.75,16.38
X$3235 366 13 367 644 645 cell_1rw
* cell instance $3236 r0 *1 106.455,16.38
X$3236 368 13 369 644 645 cell_1rw
* cell instance $3237 r0 *1 107.16,16.38
X$3237 370 13 371 644 645 cell_1rw
* cell instance $3238 r0 *1 107.865,16.38
X$3238 372 13 373 644 645 cell_1rw
* cell instance $3239 r0 *1 108.57,16.38
X$3239 374 13 375 644 645 cell_1rw
* cell instance $3240 r0 *1 109.275,16.38
X$3240 376 13 377 644 645 cell_1rw
* cell instance $3241 r0 *1 109.98,16.38
X$3241 378 13 379 644 645 cell_1rw
* cell instance $3242 r0 *1 110.685,16.38
X$3242 380 13 381 644 645 cell_1rw
* cell instance $3243 r0 *1 111.39,16.38
X$3243 382 13 383 644 645 cell_1rw
* cell instance $3244 r0 *1 112.095,16.38
X$3244 384 13 385 644 645 cell_1rw
* cell instance $3245 r0 *1 112.8,16.38
X$3245 386 13 387 644 645 cell_1rw
* cell instance $3246 r0 *1 113.505,16.38
X$3246 388 13 389 644 645 cell_1rw
* cell instance $3247 r0 *1 114.21,16.38
X$3247 390 13 391 644 645 cell_1rw
* cell instance $3248 r0 *1 114.915,16.38
X$3248 392 13 393 644 645 cell_1rw
* cell instance $3249 r0 *1 115.62,16.38
X$3249 394 13 395 644 645 cell_1rw
* cell instance $3250 r0 *1 116.325,16.38
X$3250 396 13 397 644 645 cell_1rw
* cell instance $3251 r0 *1 117.03,16.38
X$3251 398 13 399 644 645 cell_1rw
* cell instance $3252 r0 *1 117.735,16.38
X$3252 400 13 401 644 645 cell_1rw
* cell instance $3253 r0 *1 118.44,16.38
X$3253 402 13 403 644 645 cell_1rw
* cell instance $3254 r0 *1 119.145,16.38
X$3254 404 13 405 644 645 cell_1rw
* cell instance $3255 r0 *1 119.85,16.38
X$3255 406 13 407 644 645 cell_1rw
* cell instance $3256 r0 *1 120.555,16.38
X$3256 408 13 409 644 645 cell_1rw
* cell instance $3257 r0 *1 121.26,16.38
X$3257 410 13 411 644 645 cell_1rw
* cell instance $3258 r0 *1 121.965,16.38
X$3258 412 13 413 644 645 cell_1rw
* cell instance $3259 r0 *1 122.67,16.38
X$3259 414 13 415 644 645 cell_1rw
* cell instance $3260 r0 *1 123.375,16.38
X$3260 416 13 417 644 645 cell_1rw
* cell instance $3261 r0 *1 124.08,16.38
X$3261 418 13 419 644 645 cell_1rw
* cell instance $3262 r0 *1 124.785,16.38
X$3262 420 13 421 644 645 cell_1rw
* cell instance $3263 r0 *1 125.49,16.38
X$3263 422 13 423 644 645 cell_1rw
* cell instance $3264 r0 *1 126.195,16.38
X$3264 424 13 425 644 645 cell_1rw
* cell instance $3265 r0 *1 126.9,16.38
X$3265 426 13 427 644 645 cell_1rw
* cell instance $3266 r0 *1 127.605,16.38
X$3266 428 13 429 644 645 cell_1rw
* cell instance $3267 r0 *1 128.31,16.38
X$3267 430 13 431 644 645 cell_1rw
* cell instance $3268 r0 *1 129.015,16.38
X$3268 432 13 433 644 645 cell_1rw
* cell instance $3269 r0 *1 129.72,16.38
X$3269 434 13 435 644 645 cell_1rw
* cell instance $3270 r0 *1 130.425,16.38
X$3270 436 13 437 644 645 cell_1rw
* cell instance $3271 r0 *1 131.13,16.38
X$3271 438 13 439 644 645 cell_1rw
* cell instance $3272 r0 *1 131.835,16.38
X$3272 440 13 441 644 645 cell_1rw
* cell instance $3273 r0 *1 132.54,16.38
X$3273 442 13 443 644 645 cell_1rw
* cell instance $3274 r0 *1 133.245,16.38
X$3274 444 13 445 644 645 cell_1rw
* cell instance $3275 r0 *1 133.95,16.38
X$3275 446 13 447 644 645 cell_1rw
* cell instance $3276 r0 *1 134.655,16.38
X$3276 448 13 449 644 645 cell_1rw
* cell instance $3277 r0 *1 135.36,16.38
X$3277 450 13 451 644 645 cell_1rw
* cell instance $3278 r0 *1 136.065,16.38
X$3278 452 13 453 644 645 cell_1rw
* cell instance $3279 r0 *1 136.77,16.38
X$3279 454 13 455 644 645 cell_1rw
* cell instance $3280 r0 *1 137.475,16.38
X$3280 456 13 457 644 645 cell_1rw
* cell instance $3281 r0 *1 138.18,16.38
X$3281 458 13 459 644 645 cell_1rw
* cell instance $3282 r0 *1 138.885,16.38
X$3282 460 13 461 644 645 cell_1rw
* cell instance $3283 r0 *1 139.59,16.38
X$3283 462 13 463 644 645 cell_1rw
* cell instance $3284 r0 *1 140.295,16.38
X$3284 464 13 465 644 645 cell_1rw
* cell instance $3285 r0 *1 141,16.38
X$3285 466 13 467 644 645 cell_1rw
* cell instance $3286 r0 *1 141.705,16.38
X$3286 468 13 469 644 645 cell_1rw
* cell instance $3287 r0 *1 142.41,16.38
X$3287 470 13 471 644 645 cell_1rw
* cell instance $3288 r0 *1 143.115,16.38
X$3288 472 13 473 644 645 cell_1rw
* cell instance $3289 r0 *1 143.82,16.38
X$3289 474 13 475 644 645 cell_1rw
* cell instance $3290 r0 *1 144.525,16.38
X$3290 476 13 477 644 645 cell_1rw
* cell instance $3291 r0 *1 145.23,16.38
X$3291 478 13 479 644 645 cell_1rw
* cell instance $3292 r0 *1 145.935,16.38
X$3292 480 13 481 644 645 cell_1rw
* cell instance $3293 r0 *1 146.64,16.38
X$3293 482 13 483 644 645 cell_1rw
* cell instance $3294 r0 *1 147.345,16.38
X$3294 484 13 485 644 645 cell_1rw
* cell instance $3295 r0 *1 148.05,16.38
X$3295 486 13 487 644 645 cell_1rw
* cell instance $3296 r0 *1 148.755,16.38
X$3296 488 13 489 644 645 cell_1rw
* cell instance $3297 r0 *1 149.46,16.38
X$3297 490 13 491 644 645 cell_1rw
* cell instance $3298 r0 *1 150.165,16.38
X$3298 492 13 493 644 645 cell_1rw
* cell instance $3299 r0 *1 150.87,16.38
X$3299 494 13 495 644 645 cell_1rw
* cell instance $3300 r0 *1 151.575,16.38
X$3300 496 13 497 644 645 cell_1rw
* cell instance $3301 r0 *1 152.28,16.38
X$3301 498 13 499 644 645 cell_1rw
* cell instance $3302 r0 *1 152.985,16.38
X$3302 500 13 501 644 645 cell_1rw
* cell instance $3303 r0 *1 153.69,16.38
X$3303 502 13 503 644 645 cell_1rw
* cell instance $3304 r0 *1 154.395,16.38
X$3304 504 13 505 644 645 cell_1rw
* cell instance $3305 r0 *1 155.1,16.38
X$3305 506 13 507 644 645 cell_1rw
* cell instance $3306 r0 *1 155.805,16.38
X$3306 508 13 509 644 645 cell_1rw
* cell instance $3307 r0 *1 156.51,16.38
X$3307 510 13 511 644 645 cell_1rw
* cell instance $3308 r0 *1 157.215,16.38
X$3308 512 13 513 644 645 cell_1rw
* cell instance $3309 r0 *1 157.92,16.38
X$3309 514 13 515 644 645 cell_1rw
* cell instance $3310 r0 *1 158.625,16.38
X$3310 516 13 517 644 645 cell_1rw
* cell instance $3311 r0 *1 159.33,16.38
X$3311 518 13 519 644 645 cell_1rw
* cell instance $3312 r0 *1 160.035,16.38
X$3312 520 13 521 644 645 cell_1rw
* cell instance $3313 r0 *1 160.74,16.38
X$3313 522 13 523 644 645 cell_1rw
* cell instance $3314 r0 *1 161.445,16.38
X$3314 524 13 525 644 645 cell_1rw
* cell instance $3315 r0 *1 162.15,16.38
X$3315 526 13 527 644 645 cell_1rw
* cell instance $3316 r0 *1 162.855,16.38
X$3316 528 13 529 644 645 cell_1rw
* cell instance $3317 r0 *1 163.56,16.38
X$3317 530 13 531 644 645 cell_1rw
* cell instance $3318 r0 *1 164.265,16.38
X$3318 532 13 533 644 645 cell_1rw
* cell instance $3319 r0 *1 164.97,16.38
X$3319 534 13 535 644 645 cell_1rw
* cell instance $3320 r0 *1 165.675,16.38
X$3320 536 13 537 644 645 cell_1rw
* cell instance $3321 r0 *1 166.38,16.38
X$3321 538 13 539 644 645 cell_1rw
* cell instance $3322 r0 *1 167.085,16.38
X$3322 540 13 541 644 645 cell_1rw
* cell instance $3323 r0 *1 167.79,16.38
X$3323 542 13 543 644 645 cell_1rw
* cell instance $3324 r0 *1 168.495,16.38
X$3324 544 13 545 644 645 cell_1rw
* cell instance $3325 r0 *1 169.2,16.38
X$3325 546 13 547 644 645 cell_1rw
* cell instance $3326 r0 *1 169.905,16.38
X$3326 548 13 549 644 645 cell_1rw
* cell instance $3327 r0 *1 170.61,16.38
X$3327 550 13 551 644 645 cell_1rw
* cell instance $3328 r0 *1 171.315,16.38
X$3328 552 13 553 644 645 cell_1rw
* cell instance $3329 r0 *1 172.02,16.38
X$3329 554 13 555 644 645 cell_1rw
* cell instance $3330 r0 *1 172.725,16.38
X$3330 556 13 557 644 645 cell_1rw
* cell instance $3331 r0 *1 173.43,16.38
X$3331 558 13 559 644 645 cell_1rw
* cell instance $3332 r0 *1 174.135,16.38
X$3332 560 13 561 644 645 cell_1rw
* cell instance $3333 r0 *1 174.84,16.38
X$3333 562 13 563 644 645 cell_1rw
* cell instance $3334 r0 *1 175.545,16.38
X$3334 564 13 565 644 645 cell_1rw
* cell instance $3335 r0 *1 176.25,16.38
X$3335 566 13 567 644 645 cell_1rw
* cell instance $3336 r0 *1 176.955,16.38
X$3336 568 13 569 644 645 cell_1rw
* cell instance $3337 r0 *1 177.66,16.38
X$3337 570 13 571 644 645 cell_1rw
* cell instance $3338 r0 *1 178.365,16.38
X$3338 572 13 573 644 645 cell_1rw
* cell instance $3339 r0 *1 179.07,16.38
X$3339 574 13 575 644 645 cell_1rw
* cell instance $3340 r0 *1 179.775,16.38
X$3340 576 13 577 644 645 cell_1rw
* cell instance $3341 r0 *1 180.48,16.38
X$3341 578 13 579 644 645 cell_1rw
* cell instance $3342 m0 *1 0.705,19.11
X$3342 67 14 68 644 645 cell_1rw
* cell instance $3343 m0 *1 0,19.11
X$3343 65 14 66 644 645 cell_1rw
* cell instance $3344 m0 *1 1.41,19.11
X$3344 69 14 70 644 645 cell_1rw
* cell instance $3345 m0 *1 2.115,19.11
X$3345 71 14 72 644 645 cell_1rw
* cell instance $3346 m0 *1 2.82,19.11
X$3346 73 14 74 644 645 cell_1rw
* cell instance $3347 m0 *1 3.525,19.11
X$3347 75 14 76 644 645 cell_1rw
* cell instance $3348 m0 *1 4.23,19.11
X$3348 77 14 78 644 645 cell_1rw
* cell instance $3349 m0 *1 4.935,19.11
X$3349 79 14 80 644 645 cell_1rw
* cell instance $3350 m0 *1 5.64,19.11
X$3350 81 14 82 644 645 cell_1rw
* cell instance $3351 m0 *1 6.345,19.11
X$3351 83 14 84 644 645 cell_1rw
* cell instance $3352 m0 *1 7.05,19.11
X$3352 85 14 86 644 645 cell_1rw
* cell instance $3353 m0 *1 7.755,19.11
X$3353 87 14 88 644 645 cell_1rw
* cell instance $3354 m0 *1 8.46,19.11
X$3354 89 14 90 644 645 cell_1rw
* cell instance $3355 m0 *1 9.165,19.11
X$3355 91 14 92 644 645 cell_1rw
* cell instance $3356 m0 *1 9.87,19.11
X$3356 93 14 94 644 645 cell_1rw
* cell instance $3357 m0 *1 10.575,19.11
X$3357 95 14 96 644 645 cell_1rw
* cell instance $3358 m0 *1 11.28,19.11
X$3358 97 14 98 644 645 cell_1rw
* cell instance $3359 m0 *1 11.985,19.11
X$3359 99 14 100 644 645 cell_1rw
* cell instance $3360 m0 *1 12.69,19.11
X$3360 101 14 102 644 645 cell_1rw
* cell instance $3361 m0 *1 13.395,19.11
X$3361 103 14 104 644 645 cell_1rw
* cell instance $3362 m0 *1 14.1,19.11
X$3362 105 14 106 644 645 cell_1rw
* cell instance $3363 m0 *1 14.805,19.11
X$3363 107 14 108 644 645 cell_1rw
* cell instance $3364 m0 *1 15.51,19.11
X$3364 109 14 110 644 645 cell_1rw
* cell instance $3365 m0 *1 16.215,19.11
X$3365 111 14 112 644 645 cell_1rw
* cell instance $3366 m0 *1 16.92,19.11
X$3366 113 14 114 644 645 cell_1rw
* cell instance $3367 m0 *1 17.625,19.11
X$3367 115 14 116 644 645 cell_1rw
* cell instance $3368 m0 *1 18.33,19.11
X$3368 117 14 118 644 645 cell_1rw
* cell instance $3369 m0 *1 19.035,19.11
X$3369 119 14 120 644 645 cell_1rw
* cell instance $3370 m0 *1 19.74,19.11
X$3370 121 14 122 644 645 cell_1rw
* cell instance $3371 m0 *1 20.445,19.11
X$3371 123 14 124 644 645 cell_1rw
* cell instance $3372 m0 *1 21.15,19.11
X$3372 125 14 126 644 645 cell_1rw
* cell instance $3373 m0 *1 21.855,19.11
X$3373 127 14 128 644 645 cell_1rw
* cell instance $3374 m0 *1 22.56,19.11
X$3374 129 14 130 644 645 cell_1rw
* cell instance $3375 m0 *1 23.265,19.11
X$3375 131 14 132 644 645 cell_1rw
* cell instance $3376 m0 *1 23.97,19.11
X$3376 133 14 134 644 645 cell_1rw
* cell instance $3377 m0 *1 24.675,19.11
X$3377 135 14 136 644 645 cell_1rw
* cell instance $3378 m0 *1 25.38,19.11
X$3378 137 14 138 644 645 cell_1rw
* cell instance $3379 m0 *1 26.085,19.11
X$3379 139 14 140 644 645 cell_1rw
* cell instance $3380 m0 *1 26.79,19.11
X$3380 141 14 142 644 645 cell_1rw
* cell instance $3381 m0 *1 27.495,19.11
X$3381 143 14 144 644 645 cell_1rw
* cell instance $3382 m0 *1 28.2,19.11
X$3382 145 14 146 644 645 cell_1rw
* cell instance $3383 m0 *1 28.905,19.11
X$3383 147 14 148 644 645 cell_1rw
* cell instance $3384 m0 *1 29.61,19.11
X$3384 149 14 150 644 645 cell_1rw
* cell instance $3385 m0 *1 30.315,19.11
X$3385 151 14 152 644 645 cell_1rw
* cell instance $3386 m0 *1 31.02,19.11
X$3386 153 14 154 644 645 cell_1rw
* cell instance $3387 m0 *1 31.725,19.11
X$3387 155 14 156 644 645 cell_1rw
* cell instance $3388 m0 *1 32.43,19.11
X$3388 157 14 158 644 645 cell_1rw
* cell instance $3389 m0 *1 33.135,19.11
X$3389 159 14 160 644 645 cell_1rw
* cell instance $3390 m0 *1 33.84,19.11
X$3390 161 14 162 644 645 cell_1rw
* cell instance $3391 m0 *1 34.545,19.11
X$3391 163 14 164 644 645 cell_1rw
* cell instance $3392 m0 *1 35.25,19.11
X$3392 165 14 166 644 645 cell_1rw
* cell instance $3393 m0 *1 35.955,19.11
X$3393 167 14 168 644 645 cell_1rw
* cell instance $3394 m0 *1 36.66,19.11
X$3394 169 14 170 644 645 cell_1rw
* cell instance $3395 m0 *1 37.365,19.11
X$3395 171 14 172 644 645 cell_1rw
* cell instance $3396 m0 *1 38.07,19.11
X$3396 173 14 174 644 645 cell_1rw
* cell instance $3397 m0 *1 38.775,19.11
X$3397 175 14 176 644 645 cell_1rw
* cell instance $3398 m0 *1 39.48,19.11
X$3398 177 14 178 644 645 cell_1rw
* cell instance $3399 m0 *1 40.185,19.11
X$3399 179 14 180 644 645 cell_1rw
* cell instance $3400 m0 *1 40.89,19.11
X$3400 181 14 182 644 645 cell_1rw
* cell instance $3401 m0 *1 41.595,19.11
X$3401 183 14 184 644 645 cell_1rw
* cell instance $3402 m0 *1 42.3,19.11
X$3402 185 14 186 644 645 cell_1rw
* cell instance $3403 m0 *1 43.005,19.11
X$3403 187 14 188 644 645 cell_1rw
* cell instance $3404 m0 *1 43.71,19.11
X$3404 189 14 190 644 645 cell_1rw
* cell instance $3405 m0 *1 44.415,19.11
X$3405 191 14 192 644 645 cell_1rw
* cell instance $3406 m0 *1 45.12,19.11
X$3406 193 14 194 644 645 cell_1rw
* cell instance $3407 m0 *1 45.825,19.11
X$3407 195 14 196 644 645 cell_1rw
* cell instance $3408 m0 *1 46.53,19.11
X$3408 197 14 198 644 645 cell_1rw
* cell instance $3409 m0 *1 47.235,19.11
X$3409 199 14 200 644 645 cell_1rw
* cell instance $3410 m0 *1 47.94,19.11
X$3410 201 14 202 644 645 cell_1rw
* cell instance $3411 m0 *1 48.645,19.11
X$3411 203 14 204 644 645 cell_1rw
* cell instance $3412 m0 *1 49.35,19.11
X$3412 205 14 206 644 645 cell_1rw
* cell instance $3413 m0 *1 50.055,19.11
X$3413 207 14 208 644 645 cell_1rw
* cell instance $3414 m0 *1 50.76,19.11
X$3414 209 14 210 644 645 cell_1rw
* cell instance $3415 m0 *1 51.465,19.11
X$3415 211 14 212 644 645 cell_1rw
* cell instance $3416 m0 *1 52.17,19.11
X$3416 213 14 214 644 645 cell_1rw
* cell instance $3417 m0 *1 52.875,19.11
X$3417 215 14 216 644 645 cell_1rw
* cell instance $3418 m0 *1 53.58,19.11
X$3418 217 14 218 644 645 cell_1rw
* cell instance $3419 m0 *1 54.285,19.11
X$3419 219 14 220 644 645 cell_1rw
* cell instance $3420 m0 *1 54.99,19.11
X$3420 221 14 222 644 645 cell_1rw
* cell instance $3421 m0 *1 55.695,19.11
X$3421 223 14 224 644 645 cell_1rw
* cell instance $3422 m0 *1 56.4,19.11
X$3422 225 14 226 644 645 cell_1rw
* cell instance $3423 m0 *1 57.105,19.11
X$3423 227 14 228 644 645 cell_1rw
* cell instance $3424 m0 *1 57.81,19.11
X$3424 229 14 230 644 645 cell_1rw
* cell instance $3425 m0 *1 58.515,19.11
X$3425 231 14 232 644 645 cell_1rw
* cell instance $3426 m0 *1 59.22,19.11
X$3426 233 14 234 644 645 cell_1rw
* cell instance $3427 m0 *1 59.925,19.11
X$3427 235 14 236 644 645 cell_1rw
* cell instance $3428 m0 *1 60.63,19.11
X$3428 237 14 238 644 645 cell_1rw
* cell instance $3429 m0 *1 61.335,19.11
X$3429 239 14 240 644 645 cell_1rw
* cell instance $3430 m0 *1 62.04,19.11
X$3430 241 14 242 644 645 cell_1rw
* cell instance $3431 m0 *1 62.745,19.11
X$3431 243 14 244 644 645 cell_1rw
* cell instance $3432 m0 *1 63.45,19.11
X$3432 245 14 246 644 645 cell_1rw
* cell instance $3433 m0 *1 64.155,19.11
X$3433 247 14 248 644 645 cell_1rw
* cell instance $3434 m0 *1 64.86,19.11
X$3434 249 14 250 644 645 cell_1rw
* cell instance $3435 m0 *1 65.565,19.11
X$3435 251 14 252 644 645 cell_1rw
* cell instance $3436 m0 *1 66.27,19.11
X$3436 253 14 254 644 645 cell_1rw
* cell instance $3437 m0 *1 66.975,19.11
X$3437 255 14 256 644 645 cell_1rw
* cell instance $3438 m0 *1 67.68,19.11
X$3438 257 14 258 644 645 cell_1rw
* cell instance $3439 m0 *1 68.385,19.11
X$3439 259 14 260 644 645 cell_1rw
* cell instance $3440 m0 *1 69.09,19.11
X$3440 261 14 262 644 645 cell_1rw
* cell instance $3441 m0 *1 69.795,19.11
X$3441 263 14 264 644 645 cell_1rw
* cell instance $3442 m0 *1 70.5,19.11
X$3442 265 14 266 644 645 cell_1rw
* cell instance $3443 m0 *1 71.205,19.11
X$3443 267 14 268 644 645 cell_1rw
* cell instance $3444 m0 *1 71.91,19.11
X$3444 269 14 270 644 645 cell_1rw
* cell instance $3445 m0 *1 72.615,19.11
X$3445 271 14 272 644 645 cell_1rw
* cell instance $3446 m0 *1 73.32,19.11
X$3446 273 14 274 644 645 cell_1rw
* cell instance $3447 m0 *1 74.025,19.11
X$3447 275 14 276 644 645 cell_1rw
* cell instance $3448 m0 *1 74.73,19.11
X$3448 277 14 278 644 645 cell_1rw
* cell instance $3449 m0 *1 75.435,19.11
X$3449 279 14 280 644 645 cell_1rw
* cell instance $3450 m0 *1 76.14,19.11
X$3450 281 14 282 644 645 cell_1rw
* cell instance $3451 m0 *1 76.845,19.11
X$3451 283 14 284 644 645 cell_1rw
* cell instance $3452 m0 *1 77.55,19.11
X$3452 285 14 286 644 645 cell_1rw
* cell instance $3453 m0 *1 78.255,19.11
X$3453 287 14 288 644 645 cell_1rw
* cell instance $3454 m0 *1 78.96,19.11
X$3454 289 14 290 644 645 cell_1rw
* cell instance $3455 m0 *1 79.665,19.11
X$3455 291 14 292 644 645 cell_1rw
* cell instance $3456 m0 *1 80.37,19.11
X$3456 293 14 294 644 645 cell_1rw
* cell instance $3457 m0 *1 81.075,19.11
X$3457 295 14 296 644 645 cell_1rw
* cell instance $3458 m0 *1 81.78,19.11
X$3458 297 14 298 644 645 cell_1rw
* cell instance $3459 m0 *1 82.485,19.11
X$3459 299 14 300 644 645 cell_1rw
* cell instance $3460 m0 *1 83.19,19.11
X$3460 301 14 302 644 645 cell_1rw
* cell instance $3461 m0 *1 83.895,19.11
X$3461 303 14 304 644 645 cell_1rw
* cell instance $3462 m0 *1 84.6,19.11
X$3462 305 14 306 644 645 cell_1rw
* cell instance $3463 m0 *1 85.305,19.11
X$3463 307 14 308 644 645 cell_1rw
* cell instance $3464 m0 *1 86.01,19.11
X$3464 309 14 310 644 645 cell_1rw
* cell instance $3465 m0 *1 86.715,19.11
X$3465 311 14 312 644 645 cell_1rw
* cell instance $3466 m0 *1 87.42,19.11
X$3466 313 14 314 644 645 cell_1rw
* cell instance $3467 m0 *1 88.125,19.11
X$3467 315 14 316 644 645 cell_1rw
* cell instance $3468 m0 *1 88.83,19.11
X$3468 317 14 318 644 645 cell_1rw
* cell instance $3469 m0 *1 89.535,19.11
X$3469 319 14 320 644 645 cell_1rw
* cell instance $3470 m0 *1 90.24,19.11
X$3470 321 14 323 644 645 cell_1rw
* cell instance $3471 m0 *1 90.945,19.11
X$3471 324 14 325 644 645 cell_1rw
* cell instance $3472 m0 *1 91.65,19.11
X$3472 326 14 327 644 645 cell_1rw
* cell instance $3473 m0 *1 92.355,19.11
X$3473 328 14 329 644 645 cell_1rw
* cell instance $3474 m0 *1 93.06,19.11
X$3474 330 14 331 644 645 cell_1rw
* cell instance $3475 m0 *1 93.765,19.11
X$3475 332 14 333 644 645 cell_1rw
* cell instance $3476 m0 *1 94.47,19.11
X$3476 334 14 335 644 645 cell_1rw
* cell instance $3477 m0 *1 95.175,19.11
X$3477 336 14 337 644 645 cell_1rw
* cell instance $3478 m0 *1 95.88,19.11
X$3478 338 14 339 644 645 cell_1rw
* cell instance $3479 m0 *1 96.585,19.11
X$3479 340 14 341 644 645 cell_1rw
* cell instance $3480 m0 *1 97.29,19.11
X$3480 342 14 343 644 645 cell_1rw
* cell instance $3481 m0 *1 97.995,19.11
X$3481 344 14 345 644 645 cell_1rw
* cell instance $3482 m0 *1 98.7,19.11
X$3482 346 14 347 644 645 cell_1rw
* cell instance $3483 m0 *1 99.405,19.11
X$3483 348 14 349 644 645 cell_1rw
* cell instance $3484 m0 *1 100.11,19.11
X$3484 350 14 351 644 645 cell_1rw
* cell instance $3485 m0 *1 100.815,19.11
X$3485 352 14 353 644 645 cell_1rw
* cell instance $3486 m0 *1 101.52,19.11
X$3486 354 14 355 644 645 cell_1rw
* cell instance $3487 m0 *1 102.225,19.11
X$3487 356 14 357 644 645 cell_1rw
* cell instance $3488 m0 *1 102.93,19.11
X$3488 358 14 359 644 645 cell_1rw
* cell instance $3489 m0 *1 103.635,19.11
X$3489 360 14 361 644 645 cell_1rw
* cell instance $3490 m0 *1 104.34,19.11
X$3490 362 14 363 644 645 cell_1rw
* cell instance $3491 m0 *1 105.045,19.11
X$3491 364 14 365 644 645 cell_1rw
* cell instance $3492 m0 *1 105.75,19.11
X$3492 366 14 367 644 645 cell_1rw
* cell instance $3493 m0 *1 106.455,19.11
X$3493 368 14 369 644 645 cell_1rw
* cell instance $3494 m0 *1 107.16,19.11
X$3494 370 14 371 644 645 cell_1rw
* cell instance $3495 m0 *1 107.865,19.11
X$3495 372 14 373 644 645 cell_1rw
* cell instance $3496 m0 *1 108.57,19.11
X$3496 374 14 375 644 645 cell_1rw
* cell instance $3497 m0 *1 109.275,19.11
X$3497 376 14 377 644 645 cell_1rw
* cell instance $3498 m0 *1 109.98,19.11
X$3498 378 14 379 644 645 cell_1rw
* cell instance $3499 m0 *1 110.685,19.11
X$3499 380 14 381 644 645 cell_1rw
* cell instance $3500 m0 *1 111.39,19.11
X$3500 382 14 383 644 645 cell_1rw
* cell instance $3501 m0 *1 112.095,19.11
X$3501 384 14 385 644 645 cell_1rw
* cell instance $3502 m0 *1 112.8,19.11
X$3502 386 14 387 644 645 cell_1rw
* cell instance $3503 m0 *1 113.505,19.11
X$3503 388 14 389 644 645 cell_1rw
* cell instance $3504 m0 *1 114.21,19.11
X$3504 390 14 391 644 645 cell_1rw
* cell instance $3505 m0 *1 114.915,19.11
X$3505 392 14 393 644 645 cell_1rw
* cell instance $3506 m0 *1 115.62,19.11
X$3506 394 14 395 644 645 cell_1rw
* cell instance $3507 m0 *1 116.325,19.11
X$3507 396 14 397 644 645 cell_1rw
* cell instance $3508 m0 *1 117.03,19.11
X$3508 398 14 399 644 645 cell_1rw
* cell instance $3509 m0 *1 117.735,19.11
X$3509 400 14 401 644 645 cell_1rw
* cell instance $3510 m0 *1 118.44,19.11
X$3510 402 14 403 644 645 cell_1rw
* cell instance $3511 m0 *1 119.145,19.11
X$3511 404 14 405 644 645 cell_1rw
* cell instance $3512 m0 *1 119.85,19.11
X$3512 406 14 407 644 645 cell_1rw
* cell instance $3513 m0 *1 120.555,19.11
X$3513 408 14 409 644 645 cell_1rw
* cell instance $3514 m0 *1 121.26,19.11
X$3514 410 14 411 644 645 cell_1rw
* cell instance $3515 m0 *1 121.965,19.11
X$3515 412 14 413 644 645 cell_1rw
* cell instance $3516 m0 *1 122.67,19.11
X$3516 414 14 415 644 645 cell_1rw
* cell instance $3517 m0 *1 123.375,19.11
X$3517 416 14 417 644 645 cell_1rw
* cell instance $3518 m0 *1 124.08,19.11
X$3518 418 14 419 644 645 cell_1rw
* cell instance $3519 m0 *1 124.785,19.11
X$3519 420 14 421 644 645 cell_1rw
* cell instance $3520 m0 *1 125.49,19.11
X$3520 422 14 423 644 645 cell_1rw
* cell instance $3521 m0 *1 126.195,19.11
X$3521 424 14 425 644 645 cell_1rw
* cell instance $3522 m0 *1 126.9,19.11
X$3522 426 14 427 644 645 cell_1rw
* cell instance $3523 m0 *1 127.605,19.11
X$3523 428 14 429 644 645 cell_1rw
* cell instance $3524 m0 *1 128.31,19.11
X$3524 430 14 431 644 645 cell_1rw
* cell instance $3525 m0 *1 129.015,19.11
X$3525 432 14 433 644 645 cell_1rw
* cell instance $3526 m0 *1 129.72,19.11
X$3526 434 14 435 644 645 cell_1rw
* cell instance $3527 m0 *1 130.425,19.11
X$3527 436 14 437 644 645 cell_1rw
* cell instance $3528 m0 *1 131.13,19.11
X$3528 438 14 439 644 645 cell_1rw
* cell instance $3529 m0 *1 131.835,19.11
X$3529 440 14 441 644 645 cell_1rw
* cell instance $3530 m0 *1 132.54,19.11
X$3530 442 14 443 644 645 cell_1rw
* cell instance $3531 m0 *1 133.245,19.11
X$3531 444 14 445 644 645 cell_1rw
* cell instance $3532 m0 *1 133.95,19.11
X$3532 446 14 447 644 645 cell_1rw
* cell instance $3533 m0 *1 134.655,19.11
X$3533 448 14 449 644 645 cell_1rw
* cell instance $3534 m0 *1 135.36,19.11
X$3534 450 14 451 644 645 cell_1rw
* cell instance $3535 m0 *1 136.065,19.11
X$3535 452 14 453 644 645 cell_1rw
* cell instance $3536 m0 *1 136.77,19.11
X$3536 454 14 455 644 645 cell_1rw
* cell instance $3537 m0 *1 137.475,19.11
X$3537 456 14 457 644 645 cell_1rw
* cell instance $3538 m0 *1 138.18,19.11
X$3538 458 14 459 644 645 cell_1rw
* cell instance $3539 m0 *1 138.885,19.11
X$3539 460 14 461 644 645 cell_1rw
* cell instance $3540 m0 *1 139.59,19.11
X$3540 462 14 463 644 645 cell_1rw
* cell instance $3541 m0 *1 140.295,19.11
X$3541 464 14 465 644 645 cell_1rw
* cell instance $3542 m0 *1 141,19.11
X$3542 466 14 467 644 645 cell_1rw
* cell instance $3543 m0 *1 141.705,19.11
X$3543 468 14 469 644 645 cell_1rw
* cell instance $3544 m0 *1 142.41,19.11
X$3544 470 14 471 644 645 cell_1rw
* cell instance $3545 m0 *1 143.115,19.11
X$3545 472 14 473 644 645 cell_1rw
* cell instance $3546 m0 *1 143.82,19.11
X$3546 474 14 475 644 645 cell_1rw
* cell instance $3547 m0 *1 144.525,19.11
X$3547 476 14 477 644 645 cell_1rw
* cell instance $3548 m0 *1 145.23,19.11
X$3548 478 14 479 644 645 cell_1rw
* cell instance $3549 m0 *1 145.935,19.11
X$3549 480 14 481 644 645 cell_1rw
* cell instance $3550 m0 *1 146.64,19.11
X$3550 482 14 483 644 645 cell_1rw
* cell instance $3551 m0 *1 147.345,19.11
X$3551 484 14 485 644 645 cell_1rw
* cell instance $3552 m0 *1 148.05,19.11
X$3552 486 14 487 644 645 cell_1rw
* cell instance $3553 m0 *1 148.755,19.11
X$3553 488 14 489 644 645 cell_1rw
* cell instance $3554 m0 *1 149.46,19.11
X$3554 490 14 491 644 645 cell_1rw
* cell instance $3555 m0 *1 150.165,19.11
X$3555 492 14 493 644 645 cell_1rw
* cell instance $3556 m0 *1 150.87,19.11
X$3556 494 14 495 644 645 cell_1rw
* cell instance $3557 m0 *1 151.575,19.11
X$3557 496 14 497 644 645 cell_1rw
* cell instance $3558 m0 *1 152.28,19.11
X$3558 498 14 499 644 645 cell_1rw
* cell instance $3559 m0 *1 152.985,19.11
X$3559 500 14 501 644 645 cell_1rw
* cell instance $3560 m0 *1 153.69,19.11
X$3560 502 14 503 644 645 cell_1rw
* cell instance $3561 m0 *1 154.395,19.11
X$3561 504 14 505 644 645 cell_1rw
* cell instance $3562 m0 *1 155.1,19.11
X$3562 506 14 507 644 645 cell_1rw
* cell instance $3563 m0 *1 155.805,19.11
X$3563 508 14 509 644 645 cell_1rw
* cell instance $3564 m0 *1 156.51,19.11
X$3564 510 14 511 644 645 cell_1rw
* cell instance $3565 m0 *1 157.215,19.11
X$3565 512 14 513 644 645 cell_1rw
* cell instance $3566 m0 *1 157.92,19.11
X$3566 514 14 515 644 645 cell_1rw
* cell instance $3567 m0 *1 158.625,19.11
X$3567 516 14 517 644 645 cell_1rw
* cell instance $3568 m0 *1 159.33,19.11
X$3568 518 14 519 644 645 cell_1rw
* cell instance $3569 m0 *1 160.035,19.11
X$3569 520 14 521 644 645 cell_1rw
* cell instance $3570 m0 *1 160.74,19.11
X$3570 522 14 523 644 645 cell_1rw
* cell instance $3571 m0 *1 161.445,19.11
X$3571 524 14 525 644 645 cell_1rw
* cell instance $3572 m0 *1 162.15,19.11
X$3572 526 14 527 644 645 cell_1rw
* cell instance $3573 m0 *1 162.855,19.11
X$3573 528 14 529 644 645 cell_1rw
* cell instance $3574 m0 *1 163.56,19.11
X$3574 530 14 531 644 645 cell_1rw
* cell instance $3575 m0 *1 164.265,19.11
X$3575 532 14 533 644 645 cell_1rw
* cell instance $3576 m0 *1 164.97,19.11
X$3576 534 14 535 644 645 cell_1rw
* cell instance $3577 m0 *1 165.675,19.11
X$3577 536 14 537 644 645 cell_1rw
* cell instance $3578 m0 *1 166.38,19.11
X$3578 538 14 539 644 645 cell_1rw
* cell instance $3579 m0 *1 167.085,19.11
X$3579 540 14 541 644 645 cell_1rw
* cell instance $3580 m0 *1 167.79,19.11
X$3580 542 14 543 644 645 cell_1rw
* cell instance $3581 m0 *1 168.495,19.11
X$3581 544 14 545 644 645 cell_1rw
* cell instance $3582 m0 *1 169.2,19.11
X$3582 546 14 547 644 645 cell_1rw
* cell instance $3583 m0 *1 169.905,19.11
X$3583 548 14 549 644 645 cell_1rw
* cell instance $3584 m0 *1 170.61,19.11
X$3584 550 14 551 644 645 cell_1rw
* cell instance $3585 m0 *1 171.315,19.11
X$3585 552 14 553 644 645 cell_1rw
* cell instance $3586 m0 *1 172.02,19.11
X$3586 554 14 555 644 645 cell_1rw
* cell instance $3587 m0 *1 172.725,19.11
X$3587 556 14 557 644 645 cell_1rw
* cell instance $3588 m0 *1 173.43,19.11
X$3588 558 14 559 644 645 cell_1rw
* cell instance $3589 m0 *1 174.135,19.11
X$3589 560 14 561 644 645 cell_1rw
* cell instance $3590 m0 *1 174.84,19.11
X$3590 562 14 563 644 645 cell_1rw
* cell instance $3591 m0 *1 175.545,19.11
X$3591 564 14 565 644 645 cell_1rw
* cell instance $3592 m0 *1 176.25,19.11
X$3592 566 14 567 644 645 cell_1rw
* cell instance $3593 m0 *1 176.955,19.11
X$3593 568 14 569 644 645 cell_1rw
* cell instance $3594 m0 *1 177.66,19.11
X$3594 570 14 571 644 645 cell_1rw
* cell instance $3595 m0 *1 178.365,19.11
X$3595 572 14 573 644 645 cell_1rw
* cell instance $3596 m0 *1 179.07,19.11
X$3596 574 14 575 644 645 cell_1rw
* cell instance $3597 m0 *1 179.775,19.11
X$3597 576 14 577 644 645 cell_1rw
* cell instance $3598 m0 *1 180.48,19.11
X$3598 578 14 579 644 645 cell_1rw
* cell instance $3599 r0 *1 0.705,19.11
X$3599 67 15 68 644 645 cell_1rw
* cell instance $3600 r0 *1 0,19.11
X$3600 65 15 66 644 645 cell_1rw
* cell instance $3601 r0 *1 1.41,19.11
X$3601 69 15 70 644 645 cell_1rw
* cell instance $3602 r0 *1 2.115,19.11
X$3602 71 15 72 644 645 cell_1rw
* cell instance $3603 r0 *1 2.82,19.11
X$3603 73 15 74 644 645 cell_1rw
* cell instance $3604 r0 *1 3.525,19.11
X$3604 75 15 76 644 645 cell_1rw
* cell instance $3605 r0 *1 4.23,19.11
X$3605 77 15 78 644 645 cell_1rw
* cell instance $3606 r0 *1 4.935,19.11
X$3606 79 15 80 644 645 cell_1rw
* cell instance $3607 r0 *1 5.64,19.11
X$3607 81 15 82 644 645 cell_1rw
* cell instance $3608 r0 *1 6.345,19.11
X$3608 83 15 84 644 645 cell_1rw
* cell instance $3609 r0 *1 7.05,19.11
X$3609 85 15 86 644 645 cell_1rw
* cell instance $3610 r0 *1 7.755,19.11
X$3610 87 15 88 644 645 cell_1rw
* cell instance $3611 r0 *1 8.46,19.11
X$3611 89 15 90 644 645 cell_1rw
* cell instance $3612 r0 *1 9.165,19.11
X$3612 91 15 92 644 645 cell_1rw
* cell instance $3613 r0 *1 9.87,19.11
X$3613 93 15 94 644 645 cell_1rw
* cell instance $3614 r0 *1 10.575,19.11
X$3614 95 15 96 644 645 cell_1rw
* cell instance $3615 r0 *1 11.28,19.11
X$3615 97 15 98 644 645 cell_1rw
* cell instance $3616 r0 *1 11.985,19.11
X$3616 99 15 100 644 645 cell_1rw
* cell instance $3617 r0 *1 12.69,19.11
X$3617 101 15 102 644 645 cell_1rw
* cell instance $3618 r0 *1 13.395,19.11
X$3618 103 15 104 644 645 cell_1rw
* cell instance $3619 r0 *1 14.1,19.11
X$3619 105 15 106 644 645 cell_1rw
* cell instance $3620 r0 *1 14.805,19.11
X$3620 107 15 108 644 645 cell_1rw
* cell instance $3621 r0 *1 15.51,19.11
X$3621 109 15 110 644 645 cell_1rw
* cell instance $3622 r0 *1 16.215,19.11
X$3622 111 15 112 644 645 cell_1rw
* cell instance $3623 r0 *1 16.92,19.11
X$3623 113 15 114 644 645 cell_1rw
* cell instance $3624 r0 *1 17.625,19.11
X$3624 115 15 116 644 645 cell_1rw
* cell instance $3625 r0 *1 18.33,19.11
X$3625 117 15 118 644 645 cell_1rw
* cell instance $3626 r0 *1 19.035,19.11
X$3626 119 15 120 644 645 cell_1rw
* cell instance $3627 r0 *1 19.74,19.11
X$3627 121 15 122 644 645 cell_1rw
* cell instance $3628 r0 *1 20.445,19.11
X$3628 123 15 124 644 645 cell_1rw
* cell instance $3629 r0 *1 21.15,19.11
X$3629 125 15 126 644 645 cell_1rw
* cell instance $3630 r0 *1 21.855,19.11
X$3630 127 15 128 644 645 cell_1rw
* cell instance $3631 r0 *1 22.56,19.11
X$3631 129 15 130 644 645 cell_1rw
* cell instance $3632 r0 *1 23.265,19.11
X$3632 131 15 132 644 645 cell_1rw
* cell instance $3633 r0 *1 23.97,19.11
X$3633 133 15 134 644 645 cell_1rw
* cell instance $3634 r0 *1 24.675,19.11
X$3634 135 15 136 644 645 cell_1rw
* cell instance $3635 r0 *1 25.38,19.11
X$3635 137 15 138 644 645 cell_1rw
* cell instance $3636 r0 *1 26.085,19.11
X$3636 139 15 140 644 645 cell_1rw
* cell instance $3637 r0 *1 26.79,19.11
X$3637 141 15 142 644 645 cell_1rw
* cell instance $3638 r0 *1 27.495,19.11
X$3638 143 15 144 644 645 cell_1rw
* cell instance $3639 r0 *1 28.2,19.11
X$3639 145 15 146 644 645 cell_1rw
* cell instance $3640 r0 *1 28.905,19.11
X$3640 147 15 148 644 645 cell_1rw
* cell instance $3641 r0 *1 29.61,19.11
X$3641 149 15 150 644 645 cell_1rw
* cell instance $3642 r0 *1 30.315,19.11
X$3642 151 15 152 644 645 cell_1rw
* cell instance $3643 r0 *1 31.02,19.11
X$3643 153 15 154 644 645 cell_1rw
* cell instance $3644 r0 *1 31.725,19.11
X$3644 155 15 156 644 645 cell_1rw
* cell instance $3645 r0 *1 32.43,19.11
X$3645 157 15 158 644 645 cell_1rw
* cell instance $3646 r0 *1 33.135,19.11
X$3646 159 15 160 644 645 cell_1rw
* cell instance $3647 r0 *1 33.84,19.11
X$3647 161 15 162 644 645 cell_1rw
* cell instance $3648 r0 *1 34.545,19.11
X$3648 163 15 164 644 645 cell_1rw
* cell instance $3649 r0 *1 35.25,19.11
X$3649 165 15 166 644 645 cell_1rw
* cell instance $3650 r0 *1 35.955,19.11
X$3650 167 15 168 644 645 cell_1rw
* cell instance $3651 r0 *1 36.66,19.11
X$3651 169 15 170 644 645 cell_1rw
* cell instance $3652 r0 *1 37.365,19.11
X$3652 171 15 172 644 645 cell_1rw
* cell instance $3653 r0 *1 38.07,19.11
X$3653 173 15 174 644 645 cell_1rw
* cell instance $3654 r0 *1 38.775,19.11
X$3654 175 15 176 644 645 cell_1rw
* cell instance $3655 r0 *1 39.48,19.11
X$3655 177 15 178 644 645 cell_1rw
* cell instance $3656 r0 *1 40.185,19.11
X$3656 179 15 180 644 645 cell_1rw
* cell instance $3657 r0 *1 40.89,19.11
X$3657 181 15 182 644 645 cell_1rw
* cell instance $3658 r0 *1 41.595,19.11
X$3658 183 15 184 644 645 cell_1rw
* cell instance $3659 r0 *1 42.3,19.11
X$3659 185 15 186 644 645 cell_1rw
* cell instance $3660 r0 *1 43.005,19.11
X$3660 187 15 188 644 645 cell_1rw
* cell instance $3661 r0 *1 43.71,19.11
X$3661 189 15 190 644 645 cell_1rw
* cell instance $3662 r0 *1 44.415,19.11
X$3662 191 15 192 644 645 cell_1rw
* cell instance $3663 r0 *1 45.12,19.11
X$3663 193 15 194 644 645 cell_1rw
* cell instance $3664 r0 *1 45.825,19.11
X$3664 195 15 196 644 645 cell_1rw
* cell instance $3665 r0 *1 46.53,19.11
X$3665 197 15 198 644 645 cell_1rw
* cell instance $3666 r0 *1 47.235,19.11
X$3666 199 15 200 644 645 cell_1rw
* cell instance $3667 r0 *1 47.94,19.11
X$3667 201 15 202 644 645 cell_1rw
* cell instance $3668 r0 *1 48.645,19.11
X$3668 203 15 204 644 645 cell_1rw
* cell instance $3669 r0 *1 49.35,19.11
X$3669 205 15 206 644 645 cell_1rw
* cell instance $3670 r0 *1 50.055,19.11
X$3670 207 15 208 644 645 cell_1rw
* cell instance $3671 r0 *1 50.76,19.11
X$3671 209 15 210 644 645 cell_1rw
* cell instance $3672 r0 *1 51.465,19.11
X$3672 211 15 212 644 645 cell_1rw
* cell instance $3673 r0 *1 52.17,19.11
X$3673 213 15 214 644 645 cell_1rw
* cell instance $3674 r0 *1 52.875,19.11
X$3674 215 15 216 644 645 cell_1rw
* cell instance $3675 r0 *1 53.58,19.11
X$3675 217 15 218 644 645 cell_1rw
* cell instance $3676 r0 *1 54.285,19.11
X$3676 219 15 220 644 645 cell_1rw
* cell instance $3677 r0 *1 54.99,19.11
X$3677 221 15 222 644 645 cell_1rw
* cell instance $3678 r0 *1 55.695,19.11
X$3678 223 15 224 644 645 cell_1rw
* cell instance $3679 r0 *1 56.4,19.11
X$3679 225 15 226 644 645 cell_1rw
* cell instance $3680 r0 *1 57.105,19.11
X$3680 227 15 228 644 645 cell_1rw
* cell instance $3681 r0 *1 57.81,19.11
X$3681 229 15 230 644 645 cell_1rw
* cell instance $3682 r0 *1 58.515,19.11
X$3682 231 15 232 644 645 cell_1rw
* cell instance $3683 r0 *1 59.22,19.11
X$3683 233 15 234 644 645 cell_1rw
* cell instance $3684 r0 *1 59.925,19.11
X$3684 235 15 236 644 645 cell_1rw
* cell instance $3685 r0 *1 60.63,19.11
X$3685 237 15 238 644 645 cell_1rw
* cell instance $3686 r0 *1 61.335,19.11
X$3686 239 15 240 644 645 cell_1rw
* cell instance $3687 r0 *1 62.04,19.11
X$3687 241 15 242 644 645 cell_1rw
* cell instance $3688 r0 *1 62.745,19.11
X$3688 243 15 244 644 645 cell_1rw
* cell instance $3689 r0 *1 63.45,19.11
X$3689 245 15 246 644 645 cell_1rw
* cell instance $3690 r0 *1 64.155,19.11
X$3690 247 15 248 644 645 cell_1rw
* cell instance $3691 r0 *1 64.86,19.11
X$3691 249 15 250 644 645 cell_1rw
* cell instance $3692 r0 *1 65.565,19.11
X$3692 251 15 252 644 645 cell_1rw
* cell instance $3693 r0 *1 66.27,19.11
X$3693 253 15 254 644 645 cell_1rw
* cell instance $3694 r0 *1 66.975,19.11
X$3694 255 15 256 644 645 cell_1rw
* cell instance $3695 r0 *1 67.68,19.11
X$3695 257 15 258 644 645 cell_1rw
* cell instance $3696 r0 *1 68.385,19.11
X$3696 259 15 260 644 645 cell_1rw
* cell instance $3697 r0 *1 69.09,19.11
X$3697 261 15 262 644 645 cell_1rw
* cell instance $3698 r0 *1 69.795,19.11
X$3698 263 15 264 644 645 cell_1rw
* cell instance $3699 r0 *1 70.5,19.11
X$3699 265 15 266 644 645 cell_1rw
* cell instance $3700 r0 *1 71.205,19.11
X$3700 267 15 268 644 645 cell_1rw
* cell instance $3701 r0 *1 71.91,19.11
X$3701 269 15 270 644 645 cell_1rw
* cell instance $3702 r0 *1 72.615,19.11
X$3702 271 15 272 644 645 cell_1rw
* cell instance $3703 r0 *1 73.32,19.11
X$3703 273 15 274 644 645 cell_1rw
* cell instance $3704 r0 *1 74.025,19.11
X$3704 275 15 276 644 645 cell_1rw
* cell instance $3705 r0 *1 74.73,19.11
X$3705 277 15 278 644 645 cell_1rw
* cell instance $3706 r0 *1 75.435,19.11
X$3706 279 15 280 644 645 cell_1rw
* cell instance $3707 r0 *1 76.14,19.11
X$3707 281 15 282 644 645 cell_1rw
* cell instance $3708 r0 *1 76.845,19.11
X$3708 283 15 284 644 645 cell_1rw
* cell instance $3709 r0 *1 77.55,19.11
X$3709 285 15 286 644 645 cell_1rw
* cell instance $3710 r0 *1 78.255,19.11
X$3710 287 15 288 644 645 cell_1rw
* cell instance $3711 r0 *1 78.96,19.11
X$3711 289 15 290 644 645 cell_1rw
* cell instance $3712 r0 *1 79.665,19.11
X$3712 291 15 292 644 645 cell_1rw
* cell instance $3713 r0 *1 80.37,19.11
X$3713 293 15 294 644 645 cell_1rw
* cell instance $3714 r0 *1 81.075,19.11
X$3714 295 15 296 644 645 cell_1rw
* cell instance $3715 r0 *1 81.78,19.11
X$3715 297 15 298 644 645 cell_1rw
* cell instance $3716 r0 *1 82.485,19.11
X$3716 299 15 300 644 645 cell_1rw
* cell instance $3717 r0 *1 83.19,19.11
X$3717 301 15 302 644 645 cell_1rw
* cell instance $3718 r0 *1 83.895,19.11
X$3718 303 15 304 644 645 cell_1rw
* cell instance $3719 r0 *1 84.6,19.11
X$3719 305 15 306 644 645 cell_1rw
* cell instance $3720 r0 *1 85.305,19.11
X$3720 307 15 308 644 645 cell_1rw
* cell instance $3721 r0 *1 86.01,19.11
X$3721 309 15 310 644 645 cell_1rw
* cell instance $3722 r0 *1 86.715,19.11
X$3722 311 15 312 644 645 cell_1rw
* cell instance $3723 r0 *1 87.42,19.11
X$3723 313 15 314 644 645 cell_1rw
* cell instance $3724 r0 *1 88.125,19.11
X$3724 315 15 316 644 645 cell_1rw
* cell instance $3725 r0 *1 88.83,19.11
X$3725 317 15 318 644 645 cell_1rw
* cell instance $3726 r0 *1 89.535,19.11
X$3726 319 15 320 644 645 cell_1rw
* cell instance $3727 r0 *1 90.24,19.11
X$3727 321 15 323 644 645 cell_1rw
* cell instance $3728 r0 *1 90.945,19.11
X$3728 324 15 325 644 645 cell_1rw
* cell instance $3729 r0 *1 91.65,19.11
X$3729 326 15 327 644 645 cell_1rw
* cell instance $3730 r0 *1 92.355,19.11
X$3730 328 15 329 644 645 cell_1rw
* cell instance $3731 r0 *1 93.06,19.11
X$3731 330 15 331 644 645 cell_1rw
* cell instance $3732 r0 *1 93.765,19.11
X$3732 332 15 333 644 645 cell_1rw
* cell instance $3733 r0 *1 94.47,19.11
X$3733 334 15 335 644 645 cell_1rw
* cell instance $3734 r0 *1 95.175,19.11
X$3734 336 15 337 644 645 cell_1rw
* cell instance $3735 r0 *1 95.88,19.11
X$3735 338 15 339 644 645 cell_1rw
* cell instance $3736 r0 *1 96.585,19.11
X$3736 340 15 341 644 645 cell_1rw
* cell instance $3737 r0 *1 97.29,19.11
X$3737 342 15 343 644 645 cell_1rw
* cell instance $3738 r0 *1 97.995,19.11
X$3738 344 15 345 644 645 cell_1rw
* cell instance $3739 r0 *1 98.7,19.11
X$3739 346 15 347 644 645 cell_1rw
* cell instance $3740 r0 *1 99.405,19.11
X$3740 348 15 349 644 645 cell_1rw
* cell instance $3741 r0 *1 100.11,19.11
X$3741 350 15 351 644 645 cell_1rw
* cell instance $3742 r0 *1 100.815,19.11
X$3742 352 15 353 644 645 cell_1rw
* cell instance $3743 r0 *1 101.52,19.11
X$3743 354 15 355 644 645 cell_1rw
* cell instance $3744 r0 *1 102.225,19.11
X$3744 356 15 357 644 645 cell_1rw
* cell instance $3745 r0 *1 102.93,19.11
X$3745 358 15 359 644 645 cell_1rw
* cell instance $3746 r0 *1 103.635,19.11
X$3746 360 15 361 644 645 cell_1rw
* cell instance $3747 r0 *1 104.34,19.11
X$3747 362 15 363 644 645 cell_1rw
* cell instance $3748 r0 *1 105.045,19.11
X$3748 364 15 365 644 645 cell_1rw
* cell instance $3749 r0 *1 105.75,19.11
X$3749 366 15 367 644 645 cell_1rw
* cell instance $3750 r0 *1 106.455,19.11
X$3750 368 15 369 644 645 cell_1rw
* cell instance $3751 r0 *1 107.16,19.11
X$3751 370 15 371 644 645 cell_1rw
* cell instance $3752 r0 *1 107.865,19.11
X$3752 372 15 373 644 645 cell_1rw
* cell instance $3753 r0 *1 108.57,19.11
X$3753 374 15 375 644 645 cell_1rw
* cell instance $3754 r0 *1 109.275,19.11
X$3754 376 15 377 644 645 cell_1rw
* cell instance $3755 r0 *1 109.98,19.11
X$3755 378 15 379 644 645 cell_1rw
* cell instance $3756 r0 *1 110.685,19.11
X$3756 380 15 381 644 645 cell_1rw
* cell instance $3757 r0 *1 111.39,19.11
X$3757 382 15 383 644 645 cell_1rw
* cell instance $3758 r0 *1 112.095,19.11
X$3758 384 15 385 644 645 cell_1rw
* cell instance $3759 r0 *1 112.8,19.11
X$3759 386 15 387 644 645 cell_1rw
* cell instance $3760 r0 *1 113.505,19.11
X$3760 388 15 389 644 645 cell_1rw
* cell instance $3761 r0 *1 114.21,19.11
X$3761 390 15 391 644 645 cell_1rw
* cell instance $3762 r0 *1 114.915,19.11
X$3762 392 15 393 644 645 cell_1rw
* cell instance $3763 r0 *1 115.62,19.11
X$3763 394 15 395 644 645 cell_1rw
* cell instance $3764 r0 *1 116.325,19.11
X$3764 396 15 397 644 645 cell_1rw
* cell instance $3765 r0 *1 117.03,19.11
X$3765 398 15 399 644 645 cell_1rw
* cell instance $3766 r0 *1 117.735,19.11
X$3766 400 15 401 644 645 cell_1rw
* cell instance $3767 r0 *1 118.44,19.11
X$3767 402 15 403 644 645 cell_1rw
* cell instance $3768 r0 *1 119.145,19.11
X$3768 404 15 405 644 645 cell_1rw
* cell instance $3769 r0 *1 119.85,19.11
X$3769 406 15 407 644 645 cell_1rw
* cell instance $3770 r0 *1 120.555,19.11
X$3770 408 15 409 644 645 cell_1rw
* cell instance $3771 r0 *1 121.26,19.11
X$3771 410 15 411 644 645 cell_1rw
* cell instance $3772 r0 *1 121.965,19.11
X$3772 412 15 413 644 645 cell_1rw
* cell instance $3773 r0 *1 122.67,19.11
X$3773 414 15 415 644 645 cell_1rw
* cell instance $3774 r0 *1 123.375,19.11
X$3774 416 15 417 644 645 cell_1rw
* cell instance $3775 r0 *1 124.08,19.11
X$3775 418 15 419 644 645 cell_1rw
* cell instance $3776 r0 *1 124.785,19.11
X$3776 420 15 421 644 645 cell_1rw
* cell instance $3777 r0 *1 125.49,19.11
X$3777 422 15 423 644 645 cell_1rw
* cell instance $3778 r0 *1 126.195,19.11
X$3778 424 15 425 644 645 cell_1rw
* cell instance $3779 r0 *1 126.9,19.11
X$3779 426 15 427 644 645 cell_1rw
* cell instance $3780 r0 *1 127.605,19.11
X$3780 428 15 429 644 645 cell_1rw
* cell instance $3781 r0 *1 128.31,19.11
X$3781 430 15 431 644 645 cell_1rw
* cell instance $3782 r0 *1 129.015,19.11
X$3782 432 15 433 644 645 cell_1rw
* cell instance $3783 r0 *1 129.72,19.11
X$3783 434 15 435 644 645 cell_1rw
* cell instance $3784 r0 *1 130.425,19.11
X$3784 436 15 437 644 645 cell_1rw
* cell instance $3785 r0 *1 131.13,19.11
X$3785 438 15 439 644 645 cell_1rw
* cell instance $3786 r0 *1 131.835,19.11
X$3786 440 15 441 644 645 cell_1rw
* cell instance $3787 r0 *1 132.54,19.11
X$3787 442 15 443 644 645 cell_1rw
* cell instance $3788 r0 *1 133.245,19.11
X$3788 444 15 445 644 645 cell_1rw
* cell instance $3789 r0 *1 133.95,19.11
X$3789 446 15 447 644 645 cell_1rw
* cell instance $3790 r0 *1 134.655,19.11
X$3790 448 15 449 644 645 cell_1rw
* cell instance $3791 r0 *1 135.36,19.11
X$3791 450 15 451 644 645 cell_1rw
* cell instance $3792 r0 *1 136.065,19.11
X$3792 452 15 453 644 645 cell_1rw
* cell instance $3793 r0 *1 136.77,19.11
X$3793 454 15 455 644 645 cell_1rw
* cell instance $3794 r0 *1 137.475,19.11
X$3794 456 15 457 644 645 cell_1rw
* cell instance $3795 r0 *1 138.18,19.11
X$3795 458 15 459 644 645 cell_1rw
* cell instance $3796 r0 *1 138.885,19.11
X$3796 460 15 461 644 645 cell_1rw
* cell instance $3797 r0 *1 139.59,19.11
X$3797 462 15 463 644 645 cell_1rw
* cell instance $3798 r0 *1 140.295,19.11
X$3798 464 15 465 644 645 cell_1rw
* cell instance $3799 r0 *1 141,19.11
X$3799 466 15 467 644 645 cell_1rw
* cell instance $3800 r0 *1 141.705,19.11
X$3800 468 15 469 644 645 cell_1rw
* cell instance $3801 r0 *1 142.41,19.11
X$3801 470 15 471 644 645 cell_1rw
* cell instance $3802 r0 *1 143.115,19.11
X$3802 472 15 473 644 645 cell_1rw
* cell instance $3803 r0 *1 143.82,19.11
X$3803 474 15 475 644 645 cell_1rw
* cell instance $3804 r0 *1 144.525,19.11
X$3804 476 15 477 644 645 cell_1rw
* cell instance $3805 r0 *1 145.23,19.11
X$3805 478 15 479 644 645 cell_1rw
* cell instance $3806 r0 *1 145.935,19.11
X$3806 480 15 481 644 645 cell_1rw
* cell instance $3807 r0 *1 146.64,19.11
X$3807 482 15 483 644 645 cell_1rw
* cell instance $3808 r0 *1 147.345,19.11
X$3808 484 15 485 644 645 cell_1rw
* cell instance $3809 r0 *1 148.05,19.11
X$3809 486 15 487 644 645 cell_1rw
* cell instance $3810 r0 *1 148.755,19.11
X$3810 488 15 489 644 645 cell_1rw
* cell instance $3811 r0 *1 149.46,19.11
X$3811 490 15 491 644 645 cell_1rw
* cell instance $3812 r0 *1 150.165,19.11
X$3812 492 15 493 644 645 cell_1rw
* cell instance $3813 r0 *1 150.87,19.11
X$3813 494 15 495 644 645 cell_1rw
* cell instance $3814 r0 *1 151.575,19.11
X$3814 496 15 497 644 645 cell_1rw
* cell instance $3815 r0 *1 152.28,19.11
X$3815 498 15 499 644 645 cell_1rw
* cell instance $3816 r0 *1 152.985,19.11
X$3816 500 15 501 644 645 cell_1rw
* cell instance $3817 r0 *1 153.69,19.11
X$3817 502 15 503 644 645 cell_1rw
* cell instance $3818 r0 *1 154.395,19.11
X$3818 504 15 505 644 645 cell_1rw
* cell instance $3819 r0 *1 155.1,19.11
X$3819 506 15 507 644 645 cell_1rw
* cell instance $3820 r0 *1 155.805,19.11
X$3820 508 15 509 644 645 cell_1rw
* cell instance $3821 r0 *1 156.51,19.11
X$3821 510 15 511 644 645 cell_1rw
* cell instance $3822 r0 *1 157.215,19.11
X$3822 512 15 513 644 645 cell_1rw
* cell instance $3823 r0 *1 157.92,19.11
X$3823 514 15 515 644 645 cell_1rw
* cell instance $3824 r0 *1 158.625,19.11
X$3824 516 15 517 644 645 cell_1rw
* cell instance $3825 r0 *1 159.33,19.11
X$3825 518 15 519 644 645 cell_1rw
* cell instance $3826 r0 *1 160.035,19.11
X$3826 520 15 521 644 645 cell_1rw
* cell instance $3827 r0 *1 160.74,19.11
X$3827 522 15 523 644 645 cell_1rw
* cell instance $3828 r0 *1 161.445,19.11
X$3828 524 15 525 644 645 cell_1rw
* cell instance $3829 r0 *1 162.15,19.11
X$3829 526 15 527 644 645 cell_1rw
* cell instance $3830 r0 *1 162.855,19.11
X$3830 528 15 529 644 645 cell_1rw
* cell instance $3831 r0 *1 163.56,19.11
X$3831 530 15 531 644 645 cell_1rw
* cell instance $3832 r0 *1 164.265,19.11
X$3832 532 15 533 644 645 cell_1rw
* cell instance $3833 r0 *1 164.97,19.11
X$3833 534 15 535 644 645 cell_1rw
* cell instance $3834 r0 *1 165.675,19.11
X$3834 536 15 537 644 645 cell_1rw
* cell instance $3835 r0 *1 166.38,19.11
X$3835 538 15 539 644 645 cell_1rw
* cell instance $3836 r0 *1 167.085,19.11
X$3836 540 15 541 644 645 cell_1rw
* cell instance $3837 r0 *1 167.79,19.11
X$3837 542 15 543 644 645 cell_1rw
* cell instance $3838 r0 *1 168.495,19.11
X$3838 544 15 545 644 645 cell_1rw
* cell instance $3839 r0 *1 169.2,19.11
X$3839 546 15 547 644 645 cell_1rw
* cell instance $3840 r0 *1 169.905,19.11
X$3840 548 15 549 644 645 cell_1rw
* cell instance $3841 r0 *1 170.61,19.11
X$3841 550 15 551 644 645 cell_1rw
* cell instance $3842 r0 *1 171.315,19.11
X$3842 552 15 553 644 645 cell_1rw
* cell instance $3843 r0 *1 172.02,19.11
X$3843 554 15 555 644 645 cell_1rw
* cell instance $3844 r0 *1 172.725,19.11
X$3844 556 15 557 644 645 cell_1rw
* cell instance $3845 r0 *1 173.43,19.11
X$3845 558 15 559 644 645 cell_1rw
* cell instance $3846 r0 *1 174.135,19.11
X$3846 560 15 561 644 645 cell_1rw
* cell instance $3847 r0 *1 174.84,19.11
X$3847 562 15 563 644 645 cell_1rw
* cell instance $3848 r0 *1 175.545,19.11
X$3848 564 15 565 644 645 cell_1rw
* cell instance $3849 r0 *1 176.25,19.11
X$3849 566 15 567 644 645 cell_1rw
* cell instance $3850 r0 *1 176.955,19.11
X$3850 568 15 569 644 645 cell_1rw
* cell instance $3851 r0 *1 177.66,19.11
X$3851 570 15 571 644 645 cell_1rw
* cell instance $3852 r0 *1 178.365,19.11
X$3852 572 15 573 644 645 cell_1rw
* cell instance $3853 r0 *1 179.07,19.11
X$3853 574 15 575 644 645 cell_1rw
* cell instance $3854 r0 *1 179.775,19.11
X$3854 576 15 577 644 645 cell_1rw
* cell instance $3855 r0 *1 180.48,19.11
X$3855 578 15 579 644 645 cell_1rw
* cell instance $3856 m0 *1 0.705,21.84
X$3856 67 16 68 644 645 cell_1rw
* cell instance $3857 m0 *1 0,21.84
X$3857 65 16 66 644 645 cell_1rw
* cell instance $3858 m0 *1 1.41,21.84
X$3858 69 16 70 644 645 cell_1rw
* cell instance $3859 m0 *1 2.115,21.84
X$3859 71 16 72 644 645 cell_1rw
* cell instance $3860 m0 *1 2.82,21.84
X$3860 73 16 74 644 645 cell_1rw
* cell instance $3861 m0 *1 3.525,21.84
X$3861 75 16 76 644 645 cell_1rw
* cell instance $3862 m0 *1 4.23,21.84
X$3862 77 16 78 644 645 cell_1rw
* cell instance $3863 m0 *1 4.935,21.84
X$3863 79 16 80 644 645 cell_1rw
* cell instance $3864 m0 *1 5.64,21.84
X$3864 81 16 82 644 645 cell_1rw
* cell instance $3865 m0 *1 6.345,21.84
X$3865 83 16 84 644 645 cell_1rw
* cell instance $3866 m0 *1 7.05,21.84
X$3866 85 16 86 644 645 cell_1rw
* cell instance $3867 m0 *1 7.755,21.84
X$3867 87 16 88 644 645 cell_1rw
* cell instance $3868 m0 *1 8.46,21.84
X$3868 89 16 90 644 645 cell_1rw
* cell instance $3869 m0 *1 9.165,21.84
X$3869 91 16 92 644 645 cell_1rw
* cell instance $3870 m0 *1 9.87,21.84
X$3870 93 16 94 644 645 cell_1rw
* cell instance $3871 m0 *1 10.575,21.84
X$3871 95 16 96 644 645 cell_1rw
* cell instance $3872 m0 *1 11.28,21.84
X$3872 97 16 98 644 645 cell_1rw
* cell instance $3873 m0 *1 11.985,21.84
X$3873 99 16 100 644 645 cell_1rw
* cell instance $3874 m0 *1 12.69,21.84
X$3874 101 16 102 644 645 cell_1rw
* cell instance $3875 m0 *1 13.395,21.84
X$3875 103 16 104 644 645 cell_1rw
* cell instance $3876 m0 *1 14.1,21.84
X$3876 105 16 106 644 645 cell_1rw
* cell instance $3877 m0 *1 14.805,21.84
X$3877 107 16 108 644 645 cell_1rw
* cell instance $3878 m0 *1 15.51,21.84
X$3878 109 16 110 644 645 cell_1rw
* cell instance $3879 m0 *1 16.215,21.84
X$3879 111 16 112 644 645 cell_1rw
* cell instance $3880 m0 *1 16.92,21.84
X$3880 113 16 114 644 645 cell_1rw
* cell instance $3881 m0 *1 17.625,21.84
X$3881 115 16 116 644 645 cell_1rw
* cell instance $3882 m0 *1 18.33,21.84
X$3882 117 16 118 644 645 cell_1rw
* cell instance $3883 m0 *1 19.035,21.84
X$3883 119 16 120 644 645 cell_1rw
* cell instance $3884 m0 *1 19.74,21.84
X$3884 121 16 122 644 645 cell_1rw
* cell instance $3885 m0 *1 20.445,21.84
X$3885 123 16 124 644 645 cell_1rw
* cell instance $3886 m0 *1 21.15,21.84
X$3886 125 16 126 644 645 cell_1rw
* cell instance $3887 m0 *1 21.855,21.84
X$3887 127 16 128 644 645 cell_1rw
* cell instance $3888 m0 *1 22.56,21.84
X$3888 129 16 130 644 645 cell_1rw
* cell instance $3889 m0 *1 23.265,21.84
X$3889 131 16 132 644 645 cell_1rw
* cell instance $3890 m0 *1 23.97,21.84
X$3890 133 16 134 644 645 cell_1rw
* cell instance $3891 m0 *1 24.675,21.84
X$3891 135 16 136 644 645 cell_1rw
* cell instance $3892 m0 *1 25.38,21.84
X$3892 137 16 138 644 645 cell_1rw
* cell instance $3893 m0 *1 26.085,21.84
X$3893 139 16 140 644 645 cell_1rw
* cell instance $3894 m0 *1 26.79,21.84
X$3894 141 16 142 644 645 cell_1rw
* cell instance $3895 m0 *1 27.495,21.84
X$3895 143 16 144 644 645 cell_1rw
* cell instance $3896 m0 *1 28.2,21.84
X$3896 145 16 146 644 645 cell_1rw
* cell instance $3897 m0 *1 28.905,21.84
X$3897 147 16 148 644 645 cell_1rw
* cell instance $3898 m0 *1 29.61,21.84
X$3898 149 16 150 644 645 cell_1rw
* cell instance $3899 m0 *1 30.315,21.84
X$3899 151 16 152 644 645 cell_1rw
* cell instance $3900 m0 *1 31.02,21.84
X$3900 153 16 154 644 645 cell_1rw
* cell instance $3901 m0 *1 31.725,21.84
X$3901 155 16 156 644 645 cell_1rw
* cell instance $3902 m0 *1 32.43,21.84
X$3902 157 16 158 644 645 cell_1rw
* cell instance $3903 m0 *1 33.135,21.84
X$3903 159 16 160 644 645 cell_1rw
* cell instance $3904 m0 *1 33.84,21.84
X$3904 161 16 162 644 645 cell_1rw
* cell instance $3905 m0 *1 34.545,21.84
X$3905 163 16 164 644 645 cell_1rw
* cell instance $3906 m0 *1 35.25,21.84
X$3906 165 16 166 644 645 cell_1rw
* cell instance $3907 m0 *1 35.955,21.84
X$3907 167 16 168 644 645 cell_1rw
* cell instance $3908 m0 *1 36.66,21.84
X$3908 169 16 170 644 645 cell_1rw
* cell instance $3909 m0 *1 37.365,21.84
X$3909 171 16 172 644 645 cell_1rw
* cell instance $3910 m0 *1 38.07,21.84
X$3910 173 16 174 644 645 cell_1rw
* cell instance $3911 m0 *1 38.775,21.84
X$3911 175 16 176 644 645 cell_1rw
* cell instance $3912 m0 *1 39.48,21.84
X$3912 177 16 178 644 645 cell_1rw
* cell instance $3913 m0 *1 40.185,21.84
X$3913 179 16 180 644 645 cell_1rw
* cell instance $3914 m0 *1 40.89,21.84
X$3914 181 16 182 644 645 cell_1rw
* cell instance $3915 m0 *1 41.595,21.84
X$3915 183 16 184 644 645 cell_1rw
* cell instance $3916 m0 *1 42.3,21.84
X$3916 185 16 186 644 645 cell_1rw
* cell instance $3917 m0 *1 43.005,21.84
X$3917 187 16 188 644 645 cell_1rw
* cell instance $3918 m0 *1 43.71,21.84
X$3918 189 16 190 644 645 cell_1rw
* cell instance $3919 m0 *1 44.415,21.84
X$3919 191 16 192 644 645 cell_1rw
* cell instance $3920 m0 *1 45.12,21.84
X$3920 193 16 194 644 645 cell_1rw
* cell instance $3921 m0 *1 45.825,21.84
X$3921 195 16 196 644 645 cell_1rw
* cell instance $3922 m0 *1 46.53,21.84
X$3922 197 16 198 644 645 cell_1rw
* cell instance $3923 m0 *1 47.235,21.84
X$3923 199 16 200 644 645 cell_1rw
* cell instance $3924 m0 *1 47.94,21.84
X$3924 201 16 202 644 645 cell_1rw
* cell instance $3925 m0 *1 48.645,21.84
X$3925 203 16 204 644 645 cell_1rw
* cell instance $3926 m0 *1 49.35,21.84
X$3926 205 16 206 644 645 cell_1rw
* cell instance $3927 m0 *1 50.055,21.84
X$3927 207 16 208 644 645 cell_1rw
* cell instance $3928 m0 *1 50.76,21.84
X$3928 209 16 210 644 645 cell_1rw
* cell instance $3929 m0 *1 51.465,21.84
X$3929 211 16 212 644 645 cell_1rw
* cell instance $3930 m0 *1 52.17,21.84
X$3930 213 16 214 644 645 cell_1rw
* cell instance $3931 m0 *1 52.875,21.84
X$3931 215 16 216 644 645 cell_1rw
* cell instance $3932 m0 *1 53.58,21.84
X$3932 217 16 218 644 645 cell_1rw
* cell instance $3933 m0 *1 54.285,21.84
X$3933 219 16 220 644 645 cell_1rw
* cell instance $3934 m0 *1 54.99,21.84
X$3934 221 16 222 644 645 cell_1rw
* cell instance $3935 m0 *1 55.695,21.84
X$3935 223 16 224 644 645 cell_1rw
* cell instance $3936 m0 *1 56.4,21.84
X$3936 225 16 226 644 645 cell_1rw
* cell instance $3937 m0 *1 57.105,21.84
X$3937 227 16 228 644 645 cell_1rw
* cell instance $3938 m0 *1 57.81,21.84
X$3938 229 16 230 644 645 cell_1rw
* cell instance $3939 m0 *1 58.515,21.84
X$3939 231 16 232 644 645 cell_1rw
* cell instance $3940 m0 *1 59.22,21.84
X$3940 233 16 234 644 645 cell_1rw
* cell instance $3941 m0 *1 59.925,21.84
X$3941 235 16 236 644 645 cell_1rw
* cell instance $3942 m0 *1 60.63,21.84
X$3942 237 16 238 644 645 cell_1rw
* cell instance $3943 m0 *1 61.335,21.84
X$3943 239 16 240 644 645 cell_1rw
* cell instance $3944 m0 *1 62.04,21.84
X$3944 241 16 242 644 645 cell_1rw
* cell instance $3945 m0 *1 62.745,21.84
X$3945 243 16 244 644 645 cell_1rw
* cell instance $3946 m0 *1 63.45,21.84
X$3946 245 16 246 644 645 cell_1rw
* cell instance $3947 m0 *1 64.155,21.84
X$3947 247 16 248 644 645 cell_1rw
* cell instance $3948 m0 *1 64.86,21.84
X$3948 249 16 250 644 645 cell_1rw
* cell instance $3949 m0 *1 65.565,21.84
X$3949 251 16 252 644 645 cell_1rw
* cell instance $3950 m0 *1 66.27,21.84
X$3950 253 16 254 644 645 cell_1rw
* cell instance $3951 m0 *1 66.975,21.84
X$3951 255 16 256 644 645 cell_1rw
* cell instance $3952 m0 *1 67.68,21.84
X$3952 257 16 258 644 645 cell_1rw
* cell instance $3953 m0 *1 68.385,21.84
X$3953 259 16 260 644 645 cell_1rw
* cell instance $3954 m0 *1 69.09,21.84
X$3954 261 16 262 644 645 cell_1rw
* cell instance $3955 m0 *1 69.795,21.84
X$3955 263 16 264 644 645 cell_1rw
* cell instance $3956 m0 *1 70.5,21.84
X$3956 265 16 266 644 645 cell_1rw
* cell instance $3957 m0 *1 71.205,21.84
X$3957 267 16 268 644 645 cell_1rw
* cell instance $3958 m0 *1 71.91,21.84
X$3958 269 16 270 644 645 cell_1rw
* cell instance $3959 m0 *1 72.615,21.84
X$3959 271 16 272 644 645 cell_1rw
* cell instance $3960 m0 *1 73.32,21.84
X$3960 273 16 274 644 645 cell_1rw
* cell instance $3961 m0 *1 74.025,21.84
X$3961 275 16 276 644 645 cell_1rw
* cell instance $3962 m0 *1 74.73,21.84
X$3962 277 16 278 644 645 cell_1rw
* cell instance $3963 m0 *1 75.435,21.84
X$3963 279 16 280 644 645 cell_1rw
* cell instance $3964 m0 *1 76.14,21.84
X$3964 281 16 282 644 645 cell_1rw
* cell instance $3965 m0 *1 76.845,21.84
X$3965 283 16 284 644 645 cell_1rw
* cell instance $3966 m0 *1 77.55,21.84
X$3966 285 16 286 644 645 cell_1rw
* cell instance $3967 m0 *1 78.255,21.84
X$3967 287 16 288 644 645 cell_1rw
* cell instance $3968 m0 *1 78.96,21.84
X$3968 289 16 290 644 645 cell_1rw
* cell instance $3969 m0 *1 79.665,21.84
X$3969 291 16 292 644 645 cell_1rw
* cell instance $3970 m0 *1 80.37,21.84
X$3970 293 16 294 644 645 cell_1rw
* cell instance $3971 m0 *1 81.075,21.84
X$3971 295 16 296 644 645 cell_1rw
* cell instance $3972 m0 *1 81.78,21.84
X$3972 297 16 298 644 645 cell_1rw
* cell instance $3973 m0 *1 82.485,21.84
X$3973 299 16 300 644 645 cell_1rw
* cell instance $3974 m0 *1 83.19,21.84
X$3974 301 16 302 644 645 cell_1rw
* cell instance $3975 m0 *1 83.895,21.84
X$3975 303 16 304 644 645 cell_1rw
* cell instance $3976 m0 *1 84.6,21.84
X$3976 305 16 306 644 645 cell_1rw
* cell instance $3977 m0 *1 85.305,21.84
X$3977 307 16 308 644 645 cell_1rw
* cell instance $3978 m0 *1 86.01,21.84
X$3978 309 16 310 644 645 cell_1rw
* cell instance $3979 m0 *1 86.715,21.84
X$3979 311 16 312 644 645 cell_1rw
* cell instance $3980 m0 *1 87.42,21.84
X$3980 313 16 314 644 645 cell_1rw
* cell instance $3981 m0 *1 88.125,21.84
X$3981 315 16 316 644 645 cell_1rw
* cell instance $3982 m0 *1 88.83,21.84
X$3982 317 16 318 644 645 cell_1rw
* cell instance $3983 m0 *1 89.535,21.84
X$3983 319 16 320 644 645 cell_1rw
* cell instance $3984 m0 *1 90.24,21.84
X$3984 321 16 323 644 645 cell_1rw
* cell instance $3985 m0 *1 90.945,21.84
X$3985 324 16 325 644 645 cell_1rw
* cell instance $3986 m0 *1 91.65,21.84
X$3986 326 16 327 644 645 cell_1rw
* cell instance $3987 m0 *1 92.355,21.84
X$3987 328 16 329 644 645 cell_1rw
* cell instance $3988 m0 *1 93.06,21.84
X$3988 330 16 331 644 645 cell_1rw
* cell instance $3989 m0 *1 93.765,21.84
X$3989 332 16 333 644 645 cell_1rw
* cell instance $3990 m0 *1 94.47,21.84
X$3990 334 16 335 644 645 cell_1rw
* cell instance $3991 m0 *1 95.175,21.84
X$3991 336 16 337 644 645 cell_1rw
* cell instance $3992 m0 *1 95.88,21.84
X$3992 338 16 339 644 645 cell_1rw
* cell instance $3993 m0 *1 96.585,21.84
X$3993 340 16 341 644 645 cell_1rw
* cell instance $3994 m0 *1 97.29,21.84
X$3994 342 16 343 644 645 cell_1rw
* cell instance $3995 m0 *1 97.995,21.84
X$3995 344 16 345 644 645 cell_1rw
* cell instance $3996 m0 *1 98.7,21.84
X$3996 346 16 347 644 645 cell_1rw
* cell instance $3997 m0 *1 99.405,21.84
X$3997 348 16 349 644 645 cell_1rw
* cell instance $3998 m0 *1 100.11,21.84
X$3998 350 16 351 644 645 cell_1rw
* cell instance $3999 m0 *1 100.815,21.84
X$3999 352 16 353 644 645 cell_1rw
* cell instance $4000 m0 *1 101.52,21.84
X$4000 354 16 355 644 645 cell_1rw
* cell instance $4001 m0 *1 102.225,21.84
X$4001 356 16 357 644 645 cell_1rw
* cell instance $4002 m0 *1 102.93,21.84
X$4002 358 16 359 644 645 cell_1rw
* cell instance $4003 m0 *1 103.635,21.84
X$4003 360 16 361 644 645 cell_1rw
* cell instance $4004 m0 *1 104.34,21.84
X$4004 362 16 363 644 645 cell_1rw
* cell instance $4005 m0 *1 105.045,21.84
X$4005 364 16 365 644 645 cell_1rw
* cell instance $4006 m0 *1 105.75,21.84
X$4006 366 16 367 644 645 cell_1rw
* cell instance $4007 m0 *1 106.455,21.84
X$4007 368 16 369 644 645 cell_1rw
* cell instance $4008 m0 *1 107.16,21.84
X$4008 370 16 371 644 645 cell_1rw
* cell instance $4009 m0 *1 107.865,21.84
X$4009 372 16 373 644 645 cell_1rw
* cell instance $4010 m0 *1 108.57,21.84
X$4010 374 16 375 644 645 cell_1rw
* cell instance $4011 m0 *1 109.275,21.84
X$4011 376 16 377 644 645 cell_1rw
* cell instance $4012 m0 *1 109.98,21.84
X$4012 378 16 379 644 645 cell_1rw
* cell instance $4013 m0 *1 110.685,21.84
X$4013 380 16 381 644 645 cell_1rw
* cell instance $4014 m0 *1 111.39,21.84
X$4014 382 16 383 644 645 cell_1rw
* cell instance $4015 m0 *1 112.095,21.84
X$4015 384 16 385 644 645 cell_1rw
* cell instance $4016 m0 *1 112.8,21.84
X$4016 386 16 387 644 645 cell_1rw
* cell instance $4017 m0 *1 113.505,21.84
X$4017 388 16 389 644 645 cell_1rw
* cell instance $4018 m0 *1 114.21,21.84
X$4018 390 16 391 644 645 cell_1rw
* cell instance $4019 m0 *1 114.915,21.84
X$4019 392 16 393 644 645 cell_1rw
* cell instance $4020 m0 *1 115.62,21.84
X$4020 394 16 395 644 645 cell_1rw
* cell instance $4021 m0 *1 116.325,21.84
X$4021 396 16 397 644 645 cell_1rw
* cell instance $4022 m0 *1 117.03,21.84
X$4022 398 16 399 644 645 cell_1rw
* cell instance $4023 m0 *1 117.735,21.84
X$4023 400 16 401 644 645 cell_1rw
* cell instance $4024 m0 *1 118.44,21.84
X$4024 402 16 403 644 645 cell_1rw
* cell instance $4025 m0 *1 119.145,21.84
X$4025 404 16 405 644 645 cell_1rw
* cell instance $4026 m0 *1 119.85,21.84
X$4026 406 16 407 644 645 cell_1rw
* cell instance $4027 m0 *1 120.555,21.84
X$4027 408 16 409 644 645 cell_1rw
* cell instance $4028 m0 *1 121.26,21.84
X$4028 410 16 411 644 645 cell_1rw
* cell instance $4029 m0 *1 121.965,21.84
X$4029 412 16 413 644 645 cell_1rw
* cell instance $4030 m0 *1 122.67,21.84
X$4030 414 16 415 644 645 cell_1rw
* cell instance $4031 m0 *1 123.375,21.84
X$4031 416 16 417 644 645 cell_1rw
* cell instance $4032 m0 *1 124.08,21.84
X$4032 418 16 419 644 645 cell_1rw
* cell instance $4033 m0 *1 124.785,21.84
X$4033 420 16 421 644 645 cell_1rw
* cell instance $4034 m0 *1 125.49,21.84
X$4034 422 16 423 644 645 cell_1rw
* cell instance $4035 m0 *1 126.195,21.84
X$4035 424 16 425 644 645 cell_1rw
* cell instance $4036 m0 *1 126.9,21.84
X$4036 426 16 427 644 645 cell_1rw
* cell instance $4037 m0 *1 127.605,21.84
X$4037 428 16 429 644 645 cell_1rw
* cell instance $4038 m0 *1 128.31,21.84
X$4038 430 16 431 644 645 cell_1rw
* cell instance $4039 m0 *1 129.015,21.84
X$4039 432 16 433 644 645 cell_1rw
* cell instance $4040 m0 *1 129.72,21.84
X$4040 434 16 435 644 645 cell_1rw
* cell instance $4041 m0 *1 130.425,21.84
X$4041 436 16 437 644 645 cell_1rw
* cell instance $4042 m0 *1 131.13,21.84
X$4042 438 16 439 644 645 cell_1rw
* cell instance $4043 m0 *1 131.835,21.84
X$4043 440 16 441 644 645 cell_1rw
* cell instance $4044 m0 *1 132.54,21.84
X$4044 442 16 443 644 645 cell_1rw
* cell instance $4045 m0 *1 133.245,21.84
X$4045 444 16 445 644 645 cell_1rw
* cell instance $4046 m0 *1 133.95,21.84
X$4046 446 16 447 644 645 cell_1rw
* cell instance $4047 m0 *1 134.655,21.84
X$4047 448 16 449 644 645 cell_1rw
* cell instance $4048 m0 *1 135.36,21.84
X$4048 450 16 451 644 645 cell_1rw
* cell instance $4049 m0 *1 136.065,21.84
X$4049 452 16 453 644 645 cell_1rw
* cell instance $4050 m0 *1 136.77,21.84
X$4050 454 16 455 644 645 cell_1rw
* cell instance $4051 m0 *1 137.475,21.84
X$4051 456 16 457 644 645 cell_1rw
* cell instance $4052 m0 *1 138.18,21.84
X$4052 458 16 459 644 645 cell_1rw
* cell instance $4053 m0 *1 138.885,21.84
X$4053 460 16 461 644 645 cell_1rw
* cell instance $4054 m0 *1 139.59,21.84
X$4054 462 16 463 644 645 cell_1rw
* cell instance $4055 m0 *1 140.295,21.84
X$4055 464 16 465 644 645 cell_1rw
* cell instance $4056 m0 *1 141,21.84
X$4056 466 16 467 644 645 cell_1rw
* cell instance $4057 m0 *1 141.705,21.84
X$4057 468 16 469 644 645 cell_1rw
* cell instance $4058 m0 *1 142.41,21.84
X$4058 470 16 471 644 645 cell_1rw
* cell instance $4059 m0 *1 143.115,21.84
X$4059 472 16 473 644 645 cell_1rw
* cell instance $4060 m0 *1 143.82,21.84
X$4060 474 16 475 644 645 cell_1rw
* cell instance $4061 m0 *1 144.525,21.84
X$4061 476 16 477 644 645 cell_1rw
* cell instance $4062 m0 *1 145.23,21.84
X$4062 478 16 479 644 645 cell_1rw
* cell instance $4063 m0 *1 145.935,21.84
X$4063 480 16 481 644 645 cell_1rw
* cell instance $4064 m0 *1 146.64,21.84
X$4064 482 16 483 644 645 cell_1rw
* cell instance $4065 m0 *1 147.345,21.84
X$4065 484 16 485 644 645 cell_1rw
* cell instance $4066 m0 *1 148.05,21.84
X$4066 486 16 487 644 645 cell_1rw
* cell instance $4067 m0 *1 148.755,21.84
X$4067 488 16 489 644 645 cell_1rw
* cell instance $4068 m0 *1 149.46,21.84
X$4068 490 16 491 644 645 cell_1rw
* cell instance $4069 m0 *1 150.165,21.84
X$4069 492 16 493 644 645 cell_1rw
* cell instance $4070 m0 *1 150.87,21.84
X$4070 494 16 495 644 645 cell_1rw
* cell instance $4071 m0 *1 151.575,21.84
X$4071 496 16 497 644 645 cell_1rw
* cell instance $4072 m0 *1 152.28,21.84
X$4072 498 16 499 644 645 cell_1rw
* cell instance $4073 m0 *1 152.985,21.84
X$4073 500 16 501 644 645 cell_1rw
* cell instance $4074 m0 *1 153.69,21.84
X$4074 502 16 503 644 645 cell_1rw
* cell instance $4075 m0 *1 154.395,21.84
X$4075 504 16 505 644 645 cell_1rw
* cell instance $4076 m0 *1 155.1,21.84
X$4076 506 16 507 644 645 cell_1rw
* cell instance $4077 m0 *1 155.805,21.84
X$4077 508 16 509 644 645 cell_1rw
* cell instance $4078 m0 *1 156.51,21.84
X$4078 510 16 511 644 645 cell_1rw
* cell instance $4079 m0 *1 157.215,21.84
X$4079 512 16 513 644 645 cell_1rw
* cell instance $4080 m0 *1 157.92,21.84
X$4080 514 16 515 644 645 cell_1rw
* cell instance $4081 m0 *1 158.625,21.84
X$4081 516 16 517 644 645 cell_1rw
* cell instance $4082 m0 *1 159.33,21.84
X$4082 518 16 519 644 645 cell_1rw
* cell instance $4083 m0 *1 160.035,21.84
X$4083 520 16 521 644 645 cell_1rw
* cell instance $4084 m0 *1 160.74,21.84
X$4084 522 16 523 644 645 cell_1rw
* cell instance $4085 m0 *1 161.445,21.84
X$4085 524 16 525 644 645 cell_1rw
* cell instance $4086 m0 *1 162.15,21.84
X$4086 526 16 527 644 645 cell_1rw
* cell instance $4087 m0 *1 162.855,21.84
X$4087 528 16 529 644 645 cell_1rw
* cell instance $4088 m0 *1 163.56,21.84
X$4088 530 16 531 644 645 cell_1rw
* cell instance $4089 m0 *1 164.265,21.84
X$4089 532 16 533 644 645 cell_1rw
* cell instance $4090 m0 *1 164.97,21.84
X$4090 534 16 535 644 645 cell_1rw
* cell instance $4091 m0 *1 165.675,21.84
X$4091 536 16 537 644 645 cell_1rw
* cell instance $4092 m0 *1 166.38,21.84
X$4092 538 16 539 644 645 cell_1rw
* cell instance $4093 m0 *1 167.085,21.84
X$4093 540 16 541 644 645 cell_1rw
* cell instance $4094 m0 *1 167.79,21.84
X$4094 542 16 543 644 645 cell_1rw
* cell instance $4095 m0 *1 168.495,21.84
X$4095 544 16 545 644 645 cell_1rw
* cell instance $4096 m0 *1 169.2,21.84
X$4096 546 16 547 644 645 cell_1rw
* cell instance $4097 m0 *1 169.905,21.84
X$4097 548 16 549 644 645 cell_1rw
* cell instance $4098 m0 *1 170.61,21.84
X$4098 550 16 551 644 645 cell_1rw
* cell instance $4099 m0 *1 171.315,21.84
X$4099 552 16 553 644 645 cell_1rw
* cell instance $4100 m0 *1 172.02,21.84
X$4100 554 16 555 644 645 cell_1rw
* cell instance $4101 m0 *1 172.725,21.84
X$4101 556 16 557 644 645 cell_1rw
* cell instance $4102 m0 *1 173.43,21.84
X$4102 558 16 559 644 645 cell_1rw
* cell instance $4103 m0 *1 174.135,21.84
X$4103 560 16 561 644 645 cell_1rw
* cell instance $4104 m0 *1 174.84,21.84
X$4104 562 16 563 644 645 cell_1rw
* cell instance $4105 m0 *1 175.545,21.84
X$4105 564 16 565 644 645 cell_1rw
* cell instance $4106 m0 *1 176.25,21.84
X$4106 566 16 567 644 645 cell_1rw
* cell instance $4107 m0 *1 176.955,21.84
X$4107 568 16 569 644 645 cell_1rw
* cell instance $4108 m0 *1 177.66,21.84
X$4108 570 16 571 644 645 cell_1rw
* cell instance $4109 m0 *1 178.365,21.84
X$4109 572 16 573 644 645 cell_1rw
* cell instance $4110 m0 *1 179.07,21.84
X$4110 574 16 575 644 645 cell_1rw
* cell instance $4111 m0 *1 179.775,21.84
X$4111 576 16 577 644 645 cell_1rw
* cell instance $4112 m0 *1 180.48,21.84
X$4112 578 16 579 644 645 cell_1rw
* cell instance $4113 r0 *1 0.705,21.84
X$4113 67 17 68 644 645 cell_1rw
* cell instance $4114 r0 *1 0,21.84
X$4114 65 17 66 644 645 cell_1rw
* cell instance $4115 r0 *1 1.41,21.84
X$4115 69 17 70 644 645 cell_1rw
* cell instance $4116 r0 *1 2.115,21.84
X$4116 71 17 72 644 645 cell_1rw
* cell instance $4117 r0 *1 2.82,21.84
X$4117 73 17 74 644 645 cell_1rw
* cell instance $4118 r0 *1 3.525,21.84
X$4118 75 17 76 644 645 cell_1rw
* cell instance $4119 r0 *1 4.23,21.84
X$4119 77 17 78 644 645 cell_1rw
* cell instance $4120 r0 *1 4.935,21.84
X$4120 79 17 80 644 645 cell_1rw
* cell instance $4121 r0 *1 5.64,21.84
X$4121 81 17 82 644 645 cell_1rw
* cell instance $4122 r0 *1 6.345,21.84
X$4122 83 17 84 644 645 cell_1rw
* cell instance $4123 r0 *1 7.05,21.84
X$4123 85 17 86 644 645 cell_1rw
* cell instance $4124 r0 *1 7.755,21.84
X$4124 87 17 88 644 645 cell_1rw
* cell instance $4125 r0 *1 8.46,21.84
X$4125 89 17 90 644 645 cell_1rw
* cell instance $4126 r0 *1 9.165,21.84
X$4126 91 17 92 644 645 cell_1rw
* cell instance $4127 r0 *1 9.87,21.84
X$4127 93 17 94 644 645 cell_1rw
* cell instance $4128 r0 *1 10.575,21.84
X$4128 95 17 96 644 645 cell_1rw
* cell instance $4129 r0 *1 11.28,21.84
X$4129 97 17 98 644 645 cell_1rw
* cell instance $4130 r0 *1 11.985,21.84
X$4130 99 17 100 644 645 cell_1rw
* cell instance $4131 r0 *1 12.69,21.84
X$4131 101 17 102 644 645 cell_1rw
* cell instance $4132 r0 *1 13.395,21.84
X$4132 103 17 104 644 645 cell_1rw
* cell instance $4133 r0 *1 14.1,21.84
X$4133 105 17 106 644 645 cell_1rw
* cell instance $4134 r0 *1 14.805,21.84
X$4134 107 17 108 644 645 cell_1rw
* cell instance $4135 r0 *1 15.51,21.84
X$4135 109 17 110 644 645 cell_1rw
* cell instance $4136 r0 *1 16.215,21.84
X$4136 111 17 112 644 645 cell_1rw
* cell instance $4137 r0 *1 16.92,21.84
X$4137 113 17 114 644 645 cell_1rw
* cell instance $4138 r0 *1 17.625,21.84
X$4138 115 17 116 644 645 cell_1rw
* cell instance $4139 r0 *1 18.33,21.84
X$4139 117 17 118 644 645 cell_1rw
* cell instance $4140 r0 *1 19.035,21.84
X$4140 119 17 120 644 645 cell_1rw
* cell instance $4141 r0 *1 19.74,21.84
X$4141 121 17 122 644 645 cell_1rw
* cell instance $4142 r0 *1 20.445,21.84
X$4142 123 17 124 644 645 cell_1rw
* cell instance $4143 r0 *1 21.15,21.84
X$4143 125 17 126 644 645 cell_1rw
* cell instance $4144 r0 *1 21.855,21.84
X$4144 127 17 128 644 645 cell_1rw
* cell instance $4145 r0 *1 22.56,21.84
X$4145 129 17 130 644 645 cell_1rw
* cell instance $4146 r0 *1 23.265,21.84
X$4146 131 17 132 644 645 cell_1rw
* cell instance $4147 r0 *1 23.97,21.84
X$4147 133 17 134 644 645 cell_1rw
* cell instance $4148 r0 *1 24.675,21.84
X$4148 135 17 136 644 645 cell_1rw
* cell instance $4149 r0 *1 25.38,21.84
X$4149 137 17 138 644 645 cell_1rw
* cell instance $4150 r0 *1 26.085,21.84
X$4150 139 17 140 644 645 cell_1rw
* cell instance $4151 r0 *1 26.79,21.84
X$4151 141 17 142 644 645 cell_1rw
* cell instance $4152 r0 *1 27.495,21.84
X$4152 143 17 144 644 645 cell_1rw
* cell instance $4153 r0 *1 28.2,21.84
X$4153 145 17 146 644 645 cell_1rw
* cell instance $4154 r0 *1 28.905,21.84
X$4154 147 17 148 644 645 cell_1rw
* cell instance $4155 r0 *1 29.61,21.84
X$4155 149 17 150 644 645 cell_1rw
* cell instance $4156 r0 *1 30.315,21.84
X$4156 151 17 152 644 645 cell_1rw
* cell instance $4157 r0 *1 31.02,21.84
X$4157 153 17 154 644 645 cell_1rw
* cell instance $4158 r0 *1 31.725,21.84
X$4158 155 17 156 644 645 cell_1rw
* cell instance $4159 r0 *1 32.43,21.84
X$4159 157 17 158 644 645 cell_1rw
* cell instance $4160 r0 *1 33.135,21.84
X$4160 159 17 160 644 645 cell_1rw
* cell instance $4161 r0 *1 33.84,21.84
X$4161 161 17 162 644 645 cell_1rw
* cell instance $4162 r0 *1 34.545,21.84
X$4162 163 17 164 644 645 cell_1rw
* cell instance $4163 r0 *1 35.25,21.84
X$4163 165 17 166 644 645 cell_1rw
* cell instance $4164 r0 *1 35.955,21.84
X$4164 167 17 168 644 645 cell_1rw
* cell instance $4165 r0 *1 36.66,21.84
X$4165 169 17 170 644 645 cell_1rw
* cell instance $4166 r0 *1 37.365,21.84
X$4166 171 17 172 644 645 cell_1rw
* cell instance $4167 r0 *1 38.07,21.84
X$4167 173 17 174 644 645 cell_1rw
* cell instance $4168 r0 *1 38.775,21.84
X$4168 175 17 176 644 645 cell_1rw
* cell instance $4169 r0 *1 39.48,21.84
X$4169 177 17 178 644 645 cell_1rw
* cell instance $4170 r0 *1 40.185,21.84
X$4170 179 17 180 644 645 cell_1rw
* cell instance $4171 r0 *1 40.89,21.84
X$4171 181 17 182 644 645 cell_1rw
* cell instance $4172 r0 *1 41.595,21.84
X$4172 183 17 184 644 645 cell_1rw
* cell instance $4173 r0 *1 42.3,21.84
X$4173 185 17 186 644 645 cell_1rw
* cell instance $4174 r0 *1 43.005,21.84
X$4174 187 17 188 644 645 cell_1rw
* cell instance $4175 r0 *1 43.71,21.84
X$4175 189 17 190 644 645 cell_1rw
* cell instance $4176 r0 *1 44.415,21.84
X$4176 191 17 192 644 645 cell_1rw
* cell instance $4177 r0 *1 45.12,21.84
X$4177 193 17 194 644 645 cell_1rw
* cell instance $4178 r0 *1 45.825,21.84
X$4178 195 17 196 644 645 cell_1rw
* cell instance $4179 r0 *1 46.53,21.84
X$4179 197 17 198 644 645 cell_1rw
* cell instance $4180 r0 *1 47.235,21.84
X$4180 199 17 200 644 645 cell_1rw
* cell instance $4181 r0 *1 47.94,21.84
X$4181 201 17 202 644 645 cell_1rw
* cell instance $4182 r0 *1 48.645,21.84
X$4182 203 17 204 644 645 cell_1rw
* cell instance $4183 r0 *1 49.35,21.84
X$4183 205 17 206 644 645 cell_1rw
* cell instance $4184 r0 *1 50.055,21.84
X$4184 207 17 208 644 645 cell_1rw
* cell instance $4185 r0 *1 50.76,21.84
X$4185 209 17 210 644 645 cell_1rw
* cell instance $4186 r0 *1 51.465,21.84
X$4186 211 17 212 644 645 cell_1rw
* cell instance $4187 r0 *1 52.17,21.84
X$4187 213 17 214 644 645 cell_1rw
* cell instance $4188 r0 *1 52.875,21.84
X$4188 215 17 216 644 645 cell_1rw
* cell instance $4189 r0 *1 53.58,21.84
X$4189 217 17 218 644 645 cell_1rw
* cell instance $4190 r0 *1 54.285,21.84
X$4190 219 17 220 644 645 cell_1rw
* cell instance $4191 r0 *1 54.99,21.84
X$4191 221 17 222 644 645 cell_1rw
* cell instance $4192 r0 *1 55.695,21.84
X$4192 223 17 224 644 645 cell_1rw
* cell instance $4193 r0 *1 56.4,21.84
X$4193 225 17 226 644 645 cell_1rw
* cell instance $4194 r0 *1 57.105,21.84
X$4194 227 17 228 644 645 cell_1rw
* cell instance $4195 r0 *1 57.81,21.84
X$4195 229 17 230 644 645 cell_1rw
* cell instance $4196 r0 *1 58.515,21.84
X$4196 231 17 232 644 645 cell_1rw
* cell instance $4197 r0 *1 59.22,21.84
X$4197 233 17 234 644 645 cell_1rw
* cell instance $4198 r0 *1 59.925,21.84
X$4198 235 17 236 644 645 cell_1rw
* cell instance $4199 r0 *1 60.63,21.84
X$4199 237 17 238 644 645 cell_1rw
* cell instance $4200 r0 *1 61.335,21.84
X$4200 239 17 240 644 645 cell_1rw
* cell instance $4201 r0 *1 62.04,21.84
X$4201 241 17 242 644 645 cell_1rw
* cell instance $4202 r0 *1 62.745,21.84
X$4202 243 17 244 644 645 cell_1rw
* cell instance $4203 r0 *1 63.45,21.84
X$4203 245 17 246 644 645 cell_1rw
* cell instance $4204 r0 *1 64.155,21.84
X$4204 247 17 248 644 645 cell_1rw
* cell instance $4205 r0 *1 64.86,21.84
X$4205 249 17 250 644 645 cell_1rw
* cell instance $4206 r0 *1 65.565,21.84
X$4206 251 17 252 644 645 cell_1rw
* cell instance $4207 r0 *1 66.27,21.84
X$4207 253 17 254 644 645 cell_1rw
* cell instance $4208 r0 *1 66.975,21.84
X$4208 255 17 256 644 645 cell_1rw
* cell instance $4209 r0 *1 67.68,21.84
X$4209 257 17 258 644 645 cell_1rw
* cell instance $4210 r0 *1 68.385,21.84
X$4210 259 17 260 644 645 cell_1rw
* cell instance $4211 r0 *1 69.09,21.84
X$4211 261 17 262 644 645 cell_1rw
* cell instance $4212 r0 *1 69.795,21.84
X$4212 263 17 264 644 645 cell_1rw
* cell instance $4213 r0 *1 70.5,21.84
X$4213 265 17 266 644 645 cell_1rw
* cell instance $4214 r0 *1 71.205,21.84
X$4214 267 17 268 644 645 cell_1rw
* cell instance $4215 r0 *1 71.91,21.84
X$4215 269 17 270 644 645 cell_1rw
* cell instance $4216 r0 *1 72.615,21.84
X$4216 271 17 272 644 645 cell_1rw
* cell instance $4217 r0 *1 73.32,21.84
X$4217 273 17 274 644 645 cell_1rw
* cell instance $4218 r0 *1 74.025,21.84
X$4218 275 17 276 644 645 cell_1rw
* cell instance $4219 r0 *1 74.73,21.84
X$4219 277 17 278 644 645 cell_1rw
* cell instance $4220 r0 *1 75.435,21.84
X$4220 279 17 280 644 645 cell_1rw
* cell instance $4221 r0 *1 76.14,21.84
X$4221 281 17 282 644 645 cell_1rw
* cell instance $4222 r0 *1 76.845,21.84
X$4222 283 17 284 644 645 cell_1rw
* cell instance $4223 r0 *1 77.55,21.84
X$4223 285 17 286 644 645 cell_1rw
* cell instance $4224 r0 *1 78.255,21.84
X$4224 287 17 288 644 645 cell_1rw
* cell instance $4225 r0 *1 78.96,21.84
X$4225 289 17 290 644 645 cell_1rw
* cell instance $4226 r0 *1 79.665,21.84
X$4226 291 17 292 644 645 cell_1rw
* cell instance $4227 r0 *1 80.37,21.84
X$4227 293 17 294 644 645 cell_1rw
* cell instance $4228 r0 *1 81.075,21.84
X$4228 295 17 296 644 645 cell_1rw
* cell instance $4229 r0 *1 81.78,21.84
X$4229 297 17 298 644 645 cell_1rw
* cell instance $4230 r0 *1 82.485,21.84
X$4230 299 17 300 644 645 cell_1rw
* cell instance $4231 r0 *1 83.19,21.84
X$4231 301 17 302 644 645 cell_1rw
* cell instance $4232 r0 *1 83.895,21.84
X$4232 303 17 304 644 645 cell_1rw
* cell instance $4233 r0 *1 84.6,21.84
X$4233 305 17 306 644 645 cell_1rw
* cell instance $4234 r0 *1 85.305,21.84
X$4234 307 17 308 644 645 cell_1rw
* cell instance $4235 r0 *1 86.01,21.84
X$4235 309 17 310 644 645 cell_1rw
* cell instance $4236 r0 *1 86.715,21.84
X$4236 311 17 312 644 645 cell_1rw
* cell instance $4237 r0 *1 87.42,21.84
X$4237 313 17 314 644 645 cell_1rw
* cell instance $4238 r0 *1 88.125,21.84
X$4238 315 17 316 644 645 cell_1rw
* cell instance $4239 r0 *1 88.83,21.84
X$4239 317 17 318 644 645 cell_1rw
* cell instance $4240 r0 *1 89.535,21.84
X$4240 319 17 320 644 645 cell_1rw
* cell instance $4241 r0 *1 90.24,21.84
X$4241 321 17 323 644 645 cell_1rw
* cell instance $4242 r0 *1 90.945,21.84
X$4242 324 17 325 644 645 cell_1rw
* cell instance $4243 r0 *1 91.65,21.84
X$4243 326 17 327 644 645 cell_1rw
* cell instance $4244 r0 *1 92.355,21.84
X$4244 328 17 329 644 645 cell_1rw
* cell instance $4245 r0 *1 93.06,21.84
X$4245 330 17 331 644 645 cell_1rw
* cell instance $4246 r0 *1 93.765,21.84
X$4246 332 17 333 644 645 cell_1rw
* cell instance $4247 r0 *1 94.47,21.84
X$4247 334 17 335 644 645 cell_1rw
* cell instance $4248 r0 *1 95.175,21.84
X$4248 336 17 337 644 645 cell_1rw
* cell instance $4249 r0 *1 95.88,21.84
X$4249 338 17 339 644 645 cell_1rw
* cell instance $4250 r0 *1 96.585,21.84
X$4250 340 17 341 644 645 cell_1rw
* cell instance $4251 r0 *1 97.29,21.84
X$4251 342 17 343 644 645 cell_1rw
* cell instance $4252 r0 *1 97.995,21.84
X$4252 344 17 345 644 645 cell_1rw
* cell instance $4253 r0 *1 98.7,21.84
X$4253 346 17 347 644 645 cell_1rw
* cell instance $4254 r0 *1 99.405,21.84
X$4254 348 17 349 644 645 cell_1rw
* cell instance $4255 r0 *1 100.11,21.84
X$4255 350 17 351 644 645 cell_1rw
* cell instance $4256 r0 *1 100.815,21.84
X$4256 352 17 353 644 645 cell_1rw
* cell instance $4257 r0 *1 101.52,21.84
X$4257 354 17 355 644 645 cell_1rw
* cell instance $4258 r0 *1 102.225,21.84
X$4258 356 17 357 644 645 cell_1rw
* cell instance $4259 r0 *1 102.93,21.84
X$4259 358 17 359 644 645 cell_1rw
* cell instance $4260 r0 *1 103.635,21.84
X$4260 360 17 361 644 645 cell_1rw
* cell instance $4261 r0 *1 104.34,21.84
X$4261 362 17 363 644 645 cell_1rw
* cell instance $4262 r0 *1 105.045,21.84
X$4262 364 17 365 644 645 cell_1rw
* cell instance $4263 r0 *1 105.75,21.84
X$4263 366 17 367 644 645 cell_1rw
* cell instance $4264 r0 *1 106.455,21.84
X$4264 368 17 369 644 645 cell_1rw
* cell instance $4265 r0 *1 107.16,21.84
X$4265 370 17 371 644 645 cell_1rw
* cell instance $4266 r0 *1 107.865,21.84
X$4266 372 17 373 644 645 cell_1rw
* cell instance $4267 r0 *1 108.57,21.84
X$4267 374 17 375 644 645 cell_1rw
* cell instance $4268 r0 *1 109.275,21.84
X$4268 376 17 377 644 645 cell_1rw
* cell instance $4269 r0 *1 109.98,21.84
X$4269 378 17 379 644 645 cell_1rw
* cell instance $4270 r0 *1 110.685,21.84
X$4270 380 17 381 644 645 cell_1rw
* cell instance $4271 r0 *1 111.39,21.84
X$4271 382 17 383 644 645 cell_1rw
* cell instance $4272 r0 *1 112.095,21.84
X$4272 384 17 385 644 645 cell_1rw
* cell instance $4273 r0 *1 112.8,21.84
X$4273 386 17 387 644 645 cell_1rw
* cell instance $4274 r0 *1 113.505,21.84
X$4274 388 17 389 644 645 cell_1rw
* cell instance $4275 r0 *1 114.21,21.84
X$4275 390 17 391 644 645 cell_1rw
* cell instance $4276 r0 *1 114.915,21.84
X$4276 392 17 393 644 645 cell_1rw
* cell instance $4277 r0 *1 115.62,21.84
X$4277 394 17 395 644 645 cell_1rw
* cell instance $4278 r0 *1 116.325,21.84
X$4278 396 17 397 644 645 cell_1rw
* cell instance $4279 r0 *1 117.03,21.84
X$4279 398 17 399 644 645 cell_1rw
* cell instance $4280 r0 *1 117.735,21.84
X$4280 400 17 401 644 645 cell_1rw
* cell instance $4281 r0 *1 118.44,21.84
X$4281 402 17 403 644 645 cell_1rw
* cell instance $4282 r0 *1 119.145,21.84
X$4282 404 17 405 644 645 cell_1rw
* cell instance $4283 r0 *1 119.85,21.84
X$4283 406 17 407 644 645 cell_1rw
* cell instance $4284 r0 *1 120.555,21.84
X$4284 408 17 409 644 645 cell_1rw
* cell instance $4285 r0 *1 121.26,21.84
X$4285 410 17 411 644 645 cell_1rw
* cell instance $4286 r0 *1 121.965,21.84
X$4286 412 17 413 644 645 cell_1rw
* cell instance $4287 r0 *1 122.67,21.84
X$4287 414 17 415 644 645 cell_1rw
* cell instance $4288 r0 *1 123.375,21.84
X$4288 416 17 417 644 645 cell_1rw
* cell instance $4289 r0 *1 124.08,21.84
X$4289 418 17 419 644 645 cell_1rw
* cell instance $4290 r0 *1 124.785,21.84
X$4290 420 17 421 644 645 cell_1rw
* cell instance $4291 r0 *1 125.49,21.84
X$4291 422 17 423 644 645 cell_1rw
* cell instance $4292 r0 *1 126.195,21.84
X$4292 424 17 425 644 645 cell_1rw
* cell instance $4293 r0 *1 126.9,21.84
X$4293 426 17 427 644 645 cell_1rw
* cell instance $4294 r0 *1 127.605,21.84
X$4294 428 17 429 644 645 cell_1rw
* cell instance $4295 r0 *1 128.31,21.84
X$4295 430 17 431 644 645 cell_1rw
* cell instance $4296 r0 *1 129.015,21.84
X$4296 432 17 433 644 645 cell_1rw
* cell instance $4297 r0 *1 129.72,21.84
X$4297 434 17 435 644 645 cell_1rw
* cell instance $4298 r0 *1 130.425,21.84
X$4298 436 17 437 644 645 cell_1rw
* cell instance $4299 r0 *1 131.13,21.84
X$4299 438 17 439 644 645 cell_1rw
* cell instance $4300 r0 *1 131.835,21.84
X$4300 440 17 441 644 645 cell_1rw
* cell instance $4301 r0 *1 132.54,21.84
X$4301 442 17 443 644 645 cell_1rw
* cell instance $4302 r0 *1 133.245,21.84
X$4302 444 17 445 644 645 cell_1rw
* cell instance $4303 r0 *1 133.95,21.84
X$4303 446 17 447 644 645 cell_1rw
* cell instance $4304 r0 *1 134.655,21.84
X$4304 448 17 449 644 645 cell_1rw
* cell instance $4305 r0 *1 135.36,21.84
X$4305 450 17 451 644 645 cell_1rw
* cell instance $4306 r0 *1 136.065,21.84
X$4306 452 17 453 644 645 cell_1rw
* cell instance $4307 r0 *1 136.77,21.84
X$4307 454 17 455 644 645 cell_1rw
* cell instance $4308 r0 *1 137.475,21.84
X$4308 456 17 457 644 645 cell_1rw
* cell instance $4309 r0 *1 138.18,21.84
X$4309 458 17 459 644 645 cell_1rw
* cell instance $4310 r0 *1 138.885,21.84
X$4310 460 17 461 644 645 cell_1rw
* cell instance $4311 r0 *1 139.59,21.84
X$4311 462 17 463 644 645 cell_1rw
* cell instance $4312 r0 *1 140.295,21.84
X$4312 464 17 465 644 645 cell_1rw
* cell instance $4313 r0 *1 141,21.84
X$4313 466 17 467 644 645 cell_1rw
* cell instance $4314 r0 *1 141.705,21.84
X$4314 468 17 469 644 645 cell_1rw
* cell instance $4315 r0 *1 142.41,21.84
X$4315 470 17 471 644 645 cell_1rw
* cell instance $4316 r0 *1 143.115,21.84
X$4316 472 17 473 644 645 cell_1rw
* cell instance $4317 r0 *1 143.82,21.84
X$4317 474 17 475 644 645 cell_1rw
* cell instance $4318 r0 *1 144.525,21.84
X$4318 476 17 477 644 645 cell_1rw
* cell instance $4319 r0 *1 145.23,21.84
X$4319 478 17 479 644 645 cell_1rw
* cell instance $4320 r0 *1 145.935,21.84
X$4320 480 17 481 644 645 cell_1rw
* cell instance $4321 r0 *1 146.64,21.84
X$4321 482 17 483 644 645 cell_1rw
* cell instance $4322 r0 *1 147.345,21.84
X$4322 484 17 485 644 645 cell_1rw
* cell instance $4323 r0 *1 148.05,21.84
X$4323 486 17 487 644 645 cell_1rw
* cell instance $4324 r0 *1 148.755,21.84
X$4324 488 17 489 644 645 cell_1rw
* cell instance $4325 r0 *1 149.46,21.84
X$4325 490 17 491 644 645 cell_1rw
* cell instance $4326 r0 *1 150.165,21.84
X$4326 492 17 493 644 645 cell_1rw
* cell instance $4327 r0 *1 150.87,21.84
X$4327 494 17 495 644 645 cell_1rw
* cell instance $4328 r0 *1 151.575,21.84
X$4328 496 17 497 644 645 cell_1rw
* cell instance $4329 r0 *1 152.28,21.84
X$4329 498 17 499 644 645 cell_1rw
* cell instance $4330 r0 *1 152.985,21.84
X$4330 500 17 501 644 645 cell_1rw
* cell instance $4331 r0 *1 153.69,21.84
X$4331 502 17 503 644 645 cell_1rw
* cell instance $4332 r0 *1 154.395,21.84
X$4332 504 17 505 644 645 cell_1rw
* cell instance $4333 r0 *1 155.1,21.84
X$4333 506 17 507 644 645 cell_1rw
* cell instance $4334 r0 *1 155.805,21.84
X$4334 508 17 509 644 645 cell_1rw
* cell instance $4335 r0 *1 156.51,21.84
X$4335 510 17 511 644 645 cell_1rw
* cell instance $4336 r0 *1 157.215,21.84
X$4336 512 17 513 644 645 cell_1rw
* cell instance $4337 r0 *1 157.92,21.84
X$4337 514 17 515 644 645 cell_1rw
* cell instance $4338 r0 *1 158.625,21.84
X$4338 516 17 517 644 645 cell_1rw
* cell instance $4339 r0 *1 159.33,21.84
X$4339 518 17 519 644 645 cell_1rw
* cell instance $4340 r0 *1 160.035,21.84
X$4340 520 17 521 644 645 cell_1rw
* cell instance $4341 r0 *1 160.74,21.84
X$4341 522 17 523 644 645 cell_1rw
* cell instance $4342 r0 *1 161.445,21.84
X$4342 524 17 525 644 645 cell_1rw
* cell instance $4343 r0 *1 162.15,21.84
X$4343 526 17 527 644 645 cell_1rw
* cell instance $4344 r0 *1 162.855,21.84
X$4344 528 17 529 644 645 cell_1rw
* cell instance $4345 r0 *1 163.56,21.84
X$4345 530 17 531 644 645 cell_1rw
* cell instance $4346 r0 *1 164.265,21.84
X$4346 532 17 533 644 645 cell_1rw
* cell instance $4347 r0 *1 164.97,21.84
X$4347 534 17 535 644 645 cell_1rw
* cell instance $4348 r0 *1 165.675,21.84
X$4348 536 17 537 644 645 cell_1rw
* cell instance $4349 r0 *1 166.38,21.84
X$4349 538 17 539 644 645 cell_1rw
* cell instance $4350 r0 *1 167.085,21.84
X$4350 540 17 541 644 645 cell_1rw
* cell instance $4351 r0 *1 167.79,21.84
X$4351 542 17 543 644 645 cell_1rw
* cell instance $4352 r0 *1 168.495,21.84
X$4352 544 17 545 644 645 cell_1rw
* cell instance $4353 r0 *1 169.2,21.84
X$4353 546 17 547 644 645 cell_1rw
* cell instance $4354 r0 *1 169.905,21.84
X$4354 548 17 549 644 645 cell_1rw
* cell instance $4355 r0 *1 170.61,21.84
X$4355 550 17 551 644 645 cell_1rw
* cell instance $4356 r0 *1 171.315,21.84
X$4356 552 17 553 644 645 cell_1rw
* cell instance $4357 r0 *1 172.02,21.84
X$4357 554 17 555 644 645 cell_1rw
* cell instance $4358 r0 *1 172.725,21.84
X$4358 556 17 557 644 645 cell_1rw
* cell instance $4359 r0 *1 173.43,21.84
X$4359 558 17 559 644 645 cell_1rw
* cell instance $4360 r0 *1 174.135,21.84
X$4360 560 17 561 644 645 cell_1rw
* cell instance $4361 r0 *1 174.84,21.84
X$4361 562 17 563 644 645 cell_1rw
* cell instance $4362 r0 *1 175.545,21.84
X$4362 564 17 565 644 645 cell_1rw
* cell instance $4363 r0 *1 176.25,21.84
X$4363 566 17 567 644 645 cell_1rw
* cell instance $4364 r0 *1 176.955,21.84
X$4364 568 17 569 644 645 cell_1rw
* cell instance $4365 r0 *1 177.66,21.84
X$4365 570 17 571 644 645 cell_1rw
* cell instance $4366 r0 *1 178.365,21.84
X$4366 572 17 573 644 645 cell_1rw
* cell instance $4367 r0 *1 179.07,21.84
X$4367 574 17 575 644 645 cell_1rw
* cell instance $4368 r0 *1 179.775,21.84
X$4368 576 17 577 644 645 cell_1rw
* cell instance $4369 r0 *1 180.48,21.84
X$4369 578 17 579 644 645 cell_1rw
* cell instance $4370 m0 *1 0.705,24.57
X$4370 67 18 68 644 645 cell_1rw
* cell instance $4371 m0 *1 0,24.57
X$4371 65 18 66 644 645 cell_1rw
* cell instance $4372 m0 *1 1.41,24.57
X$4372 69 18 70 644 645 cell_1rw
* cell instance $4373 m0 *1 2.115,24.57
X$4373 71 18 72 644 645 cell_1rw
* cell instance $4374 m0 *1 2.82,24.57
X$4374 73 18 74 644 645 cell_1rw
* cell instance $4375 m0 *1 3.525,24.57
X$4375 75 18 76 644 645 cell_1rw
* cell instance $4376 m0 *1 4.23,24.57
X$4376 77 18 78 644 645 cell_1rw
* cell instance $4377 m0 *1 4.935,24.57
X$4377 79 18 80 644 645 cell_1rw
* cell instance $4378 m0 *1 5.64,24.57
X$4378 81 18 82 644 645 cell_1rw
* cell instance $4379 m0 *1 6.345,24.57
X$4379 83 18 84 644 645 cell_1rw
* cell instance $4380 m0 *1 7.05,24.57
X$4380 85 18 86 644 645 cell_1rw
* cell instance $4381 m0 *1 7.755,24.57
X$4381 87 18 88 644 645 cell_1rw
* cell instance $4382 m0 *1 8.46,24.57
X$4382 89 18 90 644 645 cell_1rw
* cell instance $4383 m0 *1 9.165,24.57
X$4383 91 18 92 644 645 cell_1rw
* cell instance $4384 m0 *1 9.87,24.57
X$4384 93 18 94 644 645 cell_1rw
* cell instance $4385 m0 *1 10.575,24.57
X$4385 95 18 96 644 645 cell_1rw
* cell instance $4386 m0 *1 11.28,24.57
X$4386 97 18 98 644 645 cell_1rw
* cell instance $4387 m0 *1 11.985,24.57
X$4387 99 18 100 644 645 cell_1rw
* cell instance $4388 m0 *1 12.69,24.57
X$4388 101 18 102 644 645 cell_1rw
* cell instance $4389 m0 *1 13.395,24.57
X$4389 103 18 104 644 645 cell_1rw
* cell instance $4390 m0 *1 14.1,24.57
X$4390 105 18 106 644 645 cell_1rw
* cell instance $4391 m0 *1 14.805,24.57
X$4391 107 18 108 644 645 cell_1rw
* cell instance $4392 m0 *1 15.51,24.57
X$4392 109 18 110 644 645 cell_1rw
* cell instance $4393 m0 *1 16.215,24.57
X$4393 111 18 112 644 645 cell_1rw
* cell instance $4394 m0 *1 16.92,24.57
X$4394 113 18 114 644 645 cell_1rw
* cell instance $4395 m0 *1 17.625,24.57
X$4395 115 18 116 644 645 cell_1rw
* cell instance $4396 m0 *1 18.33,24.57
X$4396 117 18 118 644 645 cell_1rw
* cell instance $4397 m0 *1 19.035,24.57
X$4397 119 18 120 644 645 cell_1rw
* cell instance $4398 m0 *1 19.74,24.57
X$4398 121 18 122 644 645 cell_1rw
* cell instance $4399 m0 *1 20.445,24.57
X$4399 123 18 124 644 645 cell_1rw
* cell instance $4400 m0 *1 21.15,24.57
X$4400 125 18 126 644 645 cell_1rw
* cell instance $4401 m0 *1 21.855,24.57
X$4401 127 18 128 644 645 cell_1rw
* cell instance $4402 m0 *1 22.56,24.57
X$4402 129 18 130 644 645 cell_1rw
* cell instance $4403 m0 *1 23.265,24.57
X$4403 131 18 132 644 645 cell_1rw
* cell instance $4404 m0 *1 23.97,24.57
X$4404 133 18 134 644 645 cell_1rw
* cell instance $4405 m0 *1 24.675,24.57
X$4405 135 18 136 644 645 cell_1rw
* cell instance $4406 m0 *1 25.38,24.57
X$4406 137 18 138 644 645 cell_1rw
* cell instance $4407 m0 *1 26.085,24.57
X$4407 139 18 140 644 645 cell_1rw
* cell instance $4408 m0 *1 26.79,24.57
X$4408 141 18 142 644 645 cell_1rw
* cell instance $4409 m0 *1 27.495,24.57
X$4409 143 18 144 644 645 cell_1rw
* cell instance $4410 m0 *1 28.2,24.57
X$4410 145 18 146 644 645 cell_1rw
* cell instance $4411 m0 *1 28.905,24.57
X$4411 147 18 148 644 645 cell_1rw
* cell instance $4412 m0 *1 29.61,24.57
X$4412 149 18 150 644 645 cell_1rw
* cell instance $4413 m0 *1 30.315,24.57
X$4413 151 18 152 644 645 cell_1rw
* cell instance $4414 m0 *1 31.02,24.57
X$4414 153 18 154 644 645 cell_1rw
* cell instance $4415 m0 *1 31.725,24.57
X$4415 155 18 156 644 645 cell_1rw
* cell instance $4416 m0 *1 32.43,24.57
X$4416 157 18 158 644 645 cell_1rw
* cell instance $4417 m0 *1 33.135,24.57
X$4417 159 18 160 644 645 cell_1rw
* cell instance $4418 m0 *1 33.84,24.57
X$4418 161 18 162 644 645 cell_1rw
* cell instance $4419 m0 *1 34.545,24.57
X$4419 163 18 164 644 645 cell_1rw
* cell instance $4420 m0 *1 35.25,24.57
X$4420 165 18 166 644 645 cell_1rw
* cell instance $4421 m0 *1 35.955,24.57
X$4421 167 18 168 644 645 cell_1rw
* cell instance $4422 m0 *1 36.66,24.57
X$4422 169 18 170 644 645 cell_1rw
* cell instance $4423 m0 *1 37.365,24.57
X$4423 171 18 172 644 645 cell_1rw
* cell instance $4424 m0 *1 38.07,24.57
X$4424 173 18 174 644 645 cell_1rw
* cell instance $4425 m0 *1 38.775,24.57
X$4425 175 18 176 644 645 cell_1rw
* cell instance $4426 m0 *1 39.48,24.57
X$4426 177 18 178 644 645 cell_1rw
* cell instance $4427 m0 *1 40.185,24.57
X$4427 179 18 180 644 645 cell_1rw
* cell instance $4428 m0 *1 40.89,24.57
X$4428 181 18 182 644 645 cell_1rw
* cell instance $4429 m0 *1 41.595,24.57
X$4429 183 18 184 644 645 cell_1rw
* cell instance $4430 m0 *1 42.3,24.57
X$4430 185 18 186 644 645 cell_1rw
* cell instance $4431 m0 *1 43.005,24.57
X$4431 187 18 188 644 645 cell_1rw
* cell instance $4432 m0 *1 43.71,24.57
X$4432 189 18 190 644 645 cell_1rw
* cell instance $4433 m0 *1 44.415,24.57
X$4433 191 18 192 644 645 cell_1rw
* cell instance $4434 m0 *1 45.12,24.57
X$4434 193 18 194 644 645 cell_1rw
* cell instance $4435 m0 *1 45.825,24.57
X$4435 195 18 196 644 645 cell_1rw
* cell instance $4436 m0 *1 46.53,24.57
X$4436 197 18 198 644 645 cell_1rw
* cell instance $4437 m0 *1 47.235,24.57
X$4437 199 18 200 644 645 cell_1rw
* cell instance $4438 m0 *1 47.94,24.57
X$4438 201 18 202 644 645 cell_1rw
* cell instance $4439 m0 *1 48.645,24.57
X$4439 203 18 204 644 645 cell_1rw
* cell instance $4440 m0 *1 49.35,24.57
X$4440 205 18 206 644 645 cell_1rw
* cell instance $4441 m0 *1 50.055,24.57
X$4441 207 18 208 644 645 cell_1rw
* cell instance $4442 m0 *1 50.76,24.57
X$4442 209 18 210 644 645 cell_1rw
* cell instance $4443 m0 *1 51.465,24.57
X$4443 211 18 212 644 645 cell_1rw
* cell instance $4444 m0 *1 52.17,24.57
X$4444 213 18 214 644 645 cell_1rw
* cell instance $4445 m0 *1 52.875,24.57
X$4445 215 18 216 644 645 cell_1rw
* cell instance $4446 m0 *1 53.58,24.57
X$4446 217 18 218 644 645 cell_1rw
* cell instance $4447 m0 *1 54.285,24.57
X$4447 219 18 220 644 645 cell_1rw
* cell instance $4448 m0 *1 54.99,24.57
X$4448 221 18 222 644 645 cell_1rw
* cell instance $4449 m0 *1 55.695,24.57
X$4449 223 18 224 644 645 cell_1rw
* cell instance $4450 m0 *1 56.4,24.57
X$4450 225 18 226 644 645 cell_1rw
* cell instance $4451 m0 *1 57.105,24.57
X$4451 227 18 228 644 645 cell_1rw
* cell instance $4452 m0 *1 57.81,24.57
X$4452 229 18 230 644 645 cell_1rw
* cell instance $4453 m0 *1 58.515,24.57
X$4453 231 18 232 644 645 cell_1rw
* cell instance $4454 m0 *1 59.22,24.57
X$4454 233 18 234 644 645 cell_1rw
* cell instance $4455 m0 *1 59.925,24.57
X$4455 235 18 236 644 645 cell_1rw
* cell instance $4456 m0 *1 60.63,24.57
X$4456 237 18 238 644 645 cell_1rw
* cell instance $4457 m0 *1 61.335,24.57
X$4457 239 18 240 644 645 cell_1rw
* cell instance $4458 m0 *1 62.04,24.57
X$4458 241 18 242 644 645 cell_1rw
* cell instance $4459 m0 *1 62.745,24.57
X$4459 243 18 244 644 645 cell_1rw
* cell instance $4460 m0 *1 63.45,24.57
X$4460 245 18 246 644 645 cell_1rw
* cell instance $4461 m0 *1 64.155,24.57
X$4461 247 18 248 644 645 cell_1rw
* cell instance $4462 m0 *1 64.86,24.57
X$4462 249 18 250 644 645 cell_1rw
* cell instance $4463 m0 *1 65.565,24.57
X$4463 251 18 252 644 645 cell_1rw
* cell instance $4464 m0 *1 66.27,24.57
X$4464 253 18 254 644 645 cell_1rw
* cell instance $4465 m0 *1 66.975,24.57
X$4465 255 18 256 644 645 cell_1rw
* cell instance $4466 m0 *1 67.68,24.57
X$4466 257 18 258 644 645 cell_1rw
* cell instance $4467 m0 *1 68.385,24.57
X$4467 259 18 260 644 645 cell_1rw
* cell instance $4468 m0 *1 69.09,24.57
X$4468 261 18 262 644 645 cell_1rw
* cell instance $4469 m0 *1 69.795,24.57
X$4469 263 18 264 644 645 cell_1rw
* cell instance $4470 m0 *1 70.5,24.57
X$4470 265 18 266 644 645 cell_1rw
* cell instance $4471 m0 *1 71.205,24.57
X$4471 267 18 268 644 645 cell_1rw
* cell instance $4472 m0 *1 71.91,24.57
X$4472 269 18 270 644 645 cell_1rw
* cell instance $4473 m0 *1 72.615,24.57
X$4473 271 18 272 644 645 cell_1rw
* cell instance $4474 m0 *1 73.32,24.57
X$4474 273 18 274 644 645 cell_1rw
* cell instance $4475 m0 *1 74.025,24.57
X$4475 275 18 276 644 645 cell_1rw
* cell instance $4476 m0 *1 74.73,24.57
X$4476 277 18 278 644 645 cell_1rw
* cell instance $4477 m0 *1 75.435,24.57
X$4477 279 18 280 644 645 cell_1rw
* cell instance $4478 m0 *1 76.14,24.57
X$4478 281 18 282 644 645 cell_1rw
* cell instance $4479 m0 *1 76.845,24.57
X$4479 283 18 284 644 645 cell_1rw
* cell instance $4480 m0 *1 77.55,24.57
X$4480 285 18 286 644 645 cell_1rw
* cell instance $4481 m0 *1 78.255,24.57
X$4481 287 18 288 644 645 cell_1rw
* cell instance $4482 m0 *1 78.96,24.57
X$4482 289 18 290 644 645 cell_1rw
* cell instance $4483 m0 *1 79.665,24.57
X$4483 291 18 292 644 645 cell_1rw
* cell instance $4484 m0 *1 80.37,24.57
X$4484 293 18 294 644 645 cell_1rw
* cell instance $4485 m0 *1 81.075,24.57
X$4485 295 18 296 644 645 cell_1rw
* cell instance $4486 m0 *1 81.78,24.57
X$4486 297 18 298 644 645 cell_1rw
* cell instance $4487 m0 *1 82.485,24.57
X$4487 299 18 300 644 645 cell_1rw
* cell instance $4488 m0 *1 83.19,24.57
X$4488 301 18 302 644 645 cell_1rw
* cell instance $4489 m0 *1 83.895,24.57
X$4489 303 18 304 644 645 cell_1rw
* cell instance $4490 m0 *1 84.6,24.57
X$4490 305 18 306 644 645 cell_1rw
* cell instance $4491 m0 *1 85.305,24.57
X$4491 307 18 308 644 645 cell_1rw
* cell instance $4492 m0 *1 86.01,24.57
X$4492 309 18 310 644 645 cell_1rw
* cell instance $4493 m0 *1 86.715,24.57
X$4493 311 18 312 644 645 cell_1rw
* cell instance $4494 m0 *1 87.42,24.57
X$4494 313 18 314 644 645 cell_1rw
* cell instance $4495 m0 *1 88.125,24.57
X$4495 315 18 316 644 645 cell_1rw
* cell instance $4496 m0 *1 88.83,24.57
X$4496 317 18 318 644 645 cell_1rw
* cell instance $4497 m0 *1 89.535,24.57
X$4497 319 18 320 644 645 cell_1rw
* cell instance $4498 m0 *1 90.24,24.57
X$4498 321 18 323 644 645 cell_1rw
* cell instance $4499 m0 *1 90.945,24.57
X$4499 324 18 325 644 645 cell_1rw
* cell instance $4500 m0 *1 91.65,24.57
X$4500 326 18 327 644 645 cell_1rw
* cell instance $4501 m0 *1 92.355,24.57
X$4501 328 18 329 644 645 cell_1rw
* cell instance $4502 m0 *1 93.06,24.57
X$4502 330 18 331 644 645 cell_1rw
* cell instance $4503 m0 *1 93.765,24.57
X$4503 332 18 333 644 645 cell_1rw
* cell instance $4504 m0 *1 94.47,24.57
X$4504 334 18 335 644 645 cell_1rw
* cell instance $4505 m0 *1 95.175,24.57
X$4505 336 18 337 644 645 cell_1rw
* cell instance $4506 m0 *1 95.88,24.57
X$4506 338 18 339 644 645 cell_1rw
* cell instance $4507 m0 *1 96.585,24.57
X$4507 340 18 341 644 645 cell_1rw
* cell instance $4508 m0 *1 97.29,24.57
X$4508 342 18 343 644 645 cell_1rw
* cell instance $4509 m0 *1 97.995,24.57
X$4509 344 18 345 644 645 cell_1rw
* cell instance $4510 m0 *1 98.7,24.57
X$4510 346 18 347 644 645 cell_1rw
* cell instance $4511 m0 *1 99.405,24.57
X$4511 348 18 349 644 645 cell_1rw
* cell instance $4512 m0 *1 100.11,24.57
X$4512 350 18 351 644 645 cell_1rw
* cell instance $4513 m0 *1 100.815,24.57
X$4513 352 18 353 644 645 cell_1rw
* cell instance $4514 m0 *1 101.52,24.57
X$4514 354 18 355 644 645 cell_1rw
* cell instance $4515 m0 *1 102.225,24.57
X$4515 356 18 357 644 645 cell_1rw
* cell instance $4516 m0 *1 102.93,24.57
X$4516 358 18 359 644 645 cell_1rw
* cell instance $4517 m0 *1 103.635,24.57
X$4517 360 18 361 644 645 cell_1rw
* cell instance $4518 m0 *1 104.34,24.57
X$4518 362 18 363 644 645 cell_1rw
* cell instance $4519 m0 *1 105.045,24.57
X$4519 364 18 365 644 645 cell_1rw
* cell instance $4520 m0 *1 105.75,24.57
X$4520 366 18 367 644 645 cell_1rw
* cell instance $4521 m0 *1 106.455,24.57
X$4521 368 18 369 644 645 cell_1rw
* cell instance $4522 m0 *1 107.16,24.57
X$4522 370 18 371 644 645 cell_1rw
* cell instance $4523 m0 *1 107.865,24.57
X$4523 372 18 373 644 645 cell_1rw
* cell instance $4524 m0 *1 108.57,24.57
X$4524 374 18 375 644 645 cell_1rw
* cell instance $4525 m0 *1 109.275,24.57
X$4525 376 18 377 644 645 cell_1rw
* cell instance $4526 m0 *1 109.98,24.57
X$4526 378 18 379 644 645 cell_1rw
* cell instance $4527 m0 *1 110.685,24.57
X$4527 380 18 381 644 645 cell_1rw
* cell instance $4528 m0 *1 111.39,24.57
X$4528 382 18 383 644 645 cell_1rw
* cell instance $4529 m0 *1 112.095,24.57
X$4529 384 18 385 644 645 cell_1rw
* cell instance $4530 m0 *1 112.8,24.57
X$4530 386 18 387 644 645 cell_1rw
* cell instance $4531 m0 *1 113.505,24.57
X$4531 388 18 389 644 645 cell_1rw
* cell instance $4532 m0 *1 114.21,24.57
X$4532 390 18 391 644 645 cell_1rw
* cell instance $4533 m0 *1 114.915,24.57
X$4533 392 18 393 644 645 cell_1rw
* cell instance $4534 m0 *1 115.62,24.57
X$4534 394 18 395 644 645 cell_1rw
* cell instance $4535 m0 *1 116.325,24.57
X$4535 396 18 397 644 645 cell_1rw
* cell instance $4536 m0 *1 117.03,24.57
X$4536 398 18 399 644 645 cell_1rw
* cell instance $4537 m0 *1 117.735,24.57
X$4537 400 18 401 644 645 cell_1rw
* cell instance $4538 m0 *1 118.44,24.57
X$4538 402 18 403 644 645 cell_1rw
* cell instance $4539 m0 *1 119.145,24.57
X$4539 404 18 405 644 645 cell_1rw
* cell instance $4540 m0 *1 119.85,24.57
X$4540 406 18 407 644 645 cell_1rw
* cell instance $4541 m0 *1 120.555,24.57
X$4541 408 18 409 644 645 cell_1rw
* cell instance $4542 m0 *1 121.26,24.57
X$4542 410 18 411 644 645 cell_1rw
* cell instance $4543 m0 *1 121.965,24.57
X$4543 412 18 413 644 645 cell_1rw
* cell instance $4544 m0 *1 122.67,24.57
X$4544 414 18 415 644 645 cell_1rw
* cell instance $4545 m0 *1 123.375,24.57
X$4545 416 18 417 644 645 cell_1rw
* cell instance $4546 m0 *1 124.08,24.57
X$4546 418 18 419 644 645 cell_1rw
* cell instance $4547 m0 *1 124.785,24.57
X$4547 420 18 421 644 645 cell_1rw
* cell instance $4548 m0 *1 125.49,24.57
X$4548 422 18 423 644 645 cell_1rw
* cell instance $4549 m0 *1 126.195,24.57
X$4549 424 18 425 644 645 cell_1rw
* cell instance $4550 m0 *1 126.9,24.57
X$4550 426 18 427 644 645 cell_1rw
* cell instance $4551 m0 *1 127.605,24.57
X$4551 428 18 429 644 645 cell_1rw
* cell instance $4552 m0 *1 128.31,24.57
X$4552 430 18 431 644 645 cell_1rw
* cell instance $4553 m0 *1 129.015,24.57
X$4553 432 18 433 644 645 cell_1rw
* cell instance $4554 m0 *1 129.72,24.57
X$4554 434 18 435 644 645 cell_1rw
* cell instance $4555 m0 *1 130.425,24.57
X$4555 436 18 437 644 645 cell_1rw
* cell instance $4556 m0 *1 131.13,24.57
X$4556 438 18 439 644 645 cell_1rw
* cell instance $4557 m0 *1 131.835,24.57
X$4557 440 18 441 644 645 cell_1rw
* cell instance $4558 m0 *1 132.54,24.57
X$4558 442 18 443 644 645 cell_1rw
* cell instance $4559 m0 *1 133.245,24.57
X$4559 444 18 445 644 645 cell_1rw
* cell instance $4560 m0 *1 133.95,24.57
X$4560 446 18 447 644 645 cell_1rw
* cell instance $4561 m0 *1 134.655,24.57
X$4561 448 18 449 644 645 cell_1rw
* cell instance $4562 m0 *1 135.36,24.57
X$4562 450 18 451 644 645 cell_1rw
* cell instance $4563 m0 *1 136.065,24.57
X$4563 452 18 453 644 645 cell_1rw
* cell instance $4564 m0 *1 136.77,24.57
X$4564 454 18 455 644 645 cell_1rw
* cell instance $4565 m0 *1 137.475,24.57
X$4565 456 18 457 644 645 cell_1rw
* cell instance $4566 m0 *1 138.18,24.57
X$4566 458 18 459 644 645 cell_1rw
* cell instance $4567 m0 *1 138.885,24.57
X$4567 460 18 461 644 645 cell_1rw
* cell instance $4568 m0 *1 139.59,24.57
X$4568 462 18 463 644 645 cell_1rw
* cell instance $4569 m0 *1 140.295,24.57
X$4569 464 18 465 644 645 cell_1rw
* cell instance $4570 m0 *1 141,24.57
X$4570 466 18 467 644 645 cell_1rw
* cell instance $4571 m0 *1 141.705,24.57
X$4571 468 18 469 644 645 cell_1rw
* cell instance $4572 m0 *1 142.41,24.57
X$4572 470 18 471 644 645 cell_1rw
* cell instance $4573 m0 *1 143.115,24.57
X$4573 472 18 473 644 645 cell_1rw
* cell instance $4574 m0 *1 143.82,24.57
X$4574 474 18 475 644 645 cell_1rw
* cell instance $4575 m0 *1 144.525,24.57
X$4575 476 18 477 644 645 cell_1rw
* cell instance $4576 m0 *1 145.23,24.57
X$4576 478 18 479 644 645 cell_1rw
* cell instance $4577 m0 *1 145.935,24.57
X$4577 480 18 481 644 645 cell_1rw
* cell instance $4578 m0 *1 146.64,24.57
X$4578 482 18 483 644 645 cell_1rw
* cell instance $4579 m0 *1 147.345,24.57
X$4579 484 18 485 644 645 cell_1rw
* cell instance $4580 m0 *1 148.05,24.57
X$4580 486 18 487 644 645 cell_1rw
* cell instance $4581 m0 *1 148.755,24.57
X$4581 488 18 489 644 645 cell_1rw
* cell instance $4582 m0 *1 149.46,24.57
X$4582 490 18 491 644 645 cell_1rw
* cell instance $4583 m0 *1 150.165,24.57
X$4583 492 18 493 644 645 cell_1rw
* cell instance $4584 m0 *1 150.87,24.57
X$4584 494 18 495 644 645 cell_1rw
* cell instance $4585 m0 *1 151.575,24.57
X$4585 496 18 497 644 645 cell_1rw
* cell instance $4586 m0 *1 152.28,24.57
X$4586 498 18 499 644 645 cell_1rw
* cell instance $4587 m0 *1 152.985,24.57
X$4587 500 18 501 644 645 cell_1rw
* cell instance $4588 m0 *1 153.69,24.57
X$4588 502 18 503 644 645 cell_1rw
* cell instance $4589 m0 *1 154.395,24.57
X$4589 504 18 505 644 645 cell_1rw
* cell instance $4590 m0 *1 155.1,24.57
X$4590 506 18 507 644 645 cell_1rw
* cell instance $4591 m0 *1 155.805,24.57
X$4591 508 18 509 644 645 cell_1rw
* cell instance $4592 m0 *1 156.51,24.57
X$4592 510 18 511 644 645 cell_1rw
* cell instance $4593 m0 *1 157.215,24.57
X$4593 512 18 513 644 645 cell_1rw
* cell instance $4594 m0 *1 157.92,24.57
X$4594 514 18 515 644 645 cell_1rw
* cell instance $4595 m0 *1 158.625,24.57
X$4595 516 18 517 644 645 cell_1rw
* cell instance $4596 m0 *1 159.33,24.57
X$4596 518 18 519 644 645 cell_1rw
* cell instance $4597 m0 *1 160.035,24.57
X$4597 520 18 521 644 645 cell_1rw
* cell instance $4598 m0 *1 160.74,24.57
X$4598 522 18 523 644 645 cell_1rw
* cell instance $4599 m0 *1 161.445,24.57
X$4599 524 18 525 644 645 cell_1rw
* cell instance $4600 m0 *1 162.15,24.57
X$4600 526 18 527 644 645 cell_1rw
* cell instance $4601 m0 *1 162.855,24.57
X$4601 528 18 529 644 645 cell_1rw
* cell instance $4602 m0 *1 163.56,24.57
X$4602 530 18 531 644 645 cell_1rw
* cell instance $4603 m0 *1 164.265,24.57
X$4603 532 18 533 644 645 cell_1rw
* cell instance $4604 m0 *1 164.97,24.57
X$4604 534 18 535 644 645 cell_1rw
* cell instance $4605 m0 *1 165.675,24.57
X$4605 536 18 537 644 645 cell_1rw
* cell instance $4606 m0 *1 166.38,24.57
X$4606 538 18 539 644 645 cell_1rw
* cell instance $4607 m0 *1 167.085,24.57
X$4607 540 18 541 644 645 cell_1rw
* cell instance $4608 m0 *1 167.79,24.57
X$4608 542 18 543 644 645 cell_1rw
* cell instance $4609 m0 *1 168.495,24.57
X$4609 544 18 545 644 645 cell_1rw
* cell instance $4610 m0 *1 169.2,24.57
X$4610 546 18 547 644 645 cell_1rw
* cell instance $4611 m0 *1 169.905,24.57
X$4611 548 18 549 644 645 cell_1rw
* cell instance $4612 m0 *1 170.61,24.57
X$4612 550 18 551 644 645 cell_1rw
* cell instance $4613 m0 *1 171.315,24.57
X$4613 552 18 553 644 645 cell_1rw
* cell instance $4614 m0 *1 172.02,24.57
X$4614 554 18 555 644 645 cell_1rw
* cell instance $4615 m0 *1 172.725,24.57
X$4615 556 18 557 644 645 cell_1rw
* cell instance $4616 m0 *1 173.43,24.57
X$4616 558 18 559 644 645 cell_1rw
* cell instance $4617 m0 *1 174.135,24.57
X$4617 560 18 561 644 645 cell_1rw
* cell instance $4618 m0 *1 174.84,24.57
X$4618 562 18 563 644 645 cell_1rw
* cell instance $4619 m0 *1 175.545,24.57
X$4619 564 18 565 644 645 cell_1rw
* cell instance $4620 m0 *1 176.25,24.57
X$4620 566 18 567 644 645 cell_1rw
* cell instance $4621 m0 *1 176.955,24.57
X$4621 568 18 569 644 645 cell_1rw
* cell instance $4622 m0 *1 177.66,24.57
X$4622 570 18 571 644 645 cell_1rw
* cell instance $4623 m0 *1 178.365,24.57
X$4623 572 18 573 644 645 cell_1rw
* cell instance $4624 m0 *1 179.07,24.57
X$4624 574 18 575 644 645 cell_1rw
* cell instance $4625 m0 *1 179.775,24.57
X$4625 576 18 577 644 645 cell_1rw
* cell instance $4626 m0 *1 180.48,24.57
X$4626 578 18 579 644 645 cell_1rw
* cell instance $4627 r0 *1 0.705,24.57
X$4627 67 19 68 644 645 cell_1rw
* cell instance $4628 r0 *1 0,24.57
X$4628 65 19 66 644 645 cell_1rw
* cell instance $4629 r0 *1 1.41,24.57
X$4629 69 19 70 644 645 cell_1rw
* cell instance $4630 r0 *1 2.115,24.57
X$4630 71 19 72 644 645 cell_1rw
* cell instance $4631 r0 *1 2.82,24.57
X$4631 73 19 74 644 645 cell_1rw
* cell instance $4632 r0 *1 3.525,24.57
X$4632 75 19 76 644 645 cell_1rw
* cell instance $4633 r0 *1 4.23,24.57
X$4633 77 19 78 644 645 cell_1rw
* cell instance $4634 r0 *1 4.935,24.57
X$4634 79 19 80 644 645 cell_1rw
* cell instance $4635 r0 *1 5.64,24.57
X$4635 81 19 82 644 645 cell_1rw
* cell instance $4636 r0 *1 6.345,24.57
X$4636 83 19 84 644 645 cell_1rw
* cell instance $4637 r0 *1 7.05,24.57
X$4637 85 19 86 644 645 cell_1rw
* cell instance $4638 r0 *1 7.755,24.57
X$4638 87 19 88 644 645 cell_1rw
* cell instance $4639 r0 *1 8.46,24.57
X$4639 89 19 90 644 645 cell_1rw
* cell instance $4640 r0 *1 9.165,24.57
X$4640 91 19 92 644 645 cell_1rw
* cell instance $4641 r0 *1 9.87,24.57
X$4641 93 19 94 644 645 cell_1rw
* cell instance $4642 r0 *1 10.575,24.57
X$4642 95 19 96 644 645 cell_1rw
* cell instance $4643 r0 *1 11.28,24.57
X$4643 97 19 98 644 645 cell_1rw
* cell instance $4644 r0 *1 11.985,24.57
X$4644 99 19 100 644 645 cell_1rw
* cell instance $4645 r0 *1 12.69,24.57
X$4645 101 19 102 644 645 cell_1rw
* cell instance $4646 r0 *1 13.395,24.57
X$4646 103 19 104 644 645 cell_1rw
* cell instance $4647 r0 *1 14.1,24.57
X$4647 105 19 106 644 645 cell_1rw
* cell instance $4648 r0 *1 14.805,24.57
X$4648 107 19 108 644 645 cell_1rw
* cell instance $4649 r0 *1 15.51,24.57
X$4649 109 19 110 644 645 cell_1rw
* cell instance $4650 r0 *1 16.215,24.57
X$4650 111 19 112 644 645 cell_1rw
* cell instance $4651 r0 *1 16.92,24.57
X$4651 113 19 114 644 645 cell_1rw
* cell instance $4652 r0 *1 17.625,24.57
X$4652 115 19 116 644 645 cell_1rw
* cell instance $4653 r0 *1 18.33,24.57
X$4653 117 19 118 644 645 cell_1rw
* cell instance $4654 r0 *1 19.035,24.57
X$4654 119 19 120 644 645 cell_1rw
* cell instance $4655 r0 *1 19.74,24.57
X$4655 121 19 122 644 645 cell_1rw
* cell instance $4656 r0 *1 20.445,24.57
X$4656 123 19 124 644 645 cell_1rw
* cell instance $4657 r0 *1 21.15,24.57
X$4657 125 19 126 644 645 cell_1rw
* cell instance $4658 r0 *1 21.855,24.57
X$4658 127 19 128 644 645 cell_1rw
* cell instance $4659 r0 *1 22.56,24.57
X$4659 129 19 130 644 645 cell_1rw
* cell instance $4660 r0 *1 23.265,24.57
X$4660 131 19 132 644 645 cell_1rw
* cell instance $4661 r0 *1 23.97,24.57
X$4661 133 19 134 644 645 cell_1rw
* cell instance $4662 r0 *1 24.675,24.57
X$4662 135 19 136 644 645 cell_1rw
* cell instance $4663 r0 *1 25.38,24.57
X$4663 137 19 138 644 645 cell_1rw
* cell instance $4664 r0 *1 26.085,24.57
X$4664 139 19 140 644 645 cell_1rw
* cell instance $4665 r0 *1 26.79,24.57
X$4665 141 19 142 644 645 cell_1rw
* cell instance $4666 r0 *1 27.495,24.57
X$4666 143 19 144 644 645 cell_1rw
* cell instance $4667 r0 *1 28.2,24.57
X$4667 145 19 146 644 645 cell_1rw
* cell instance $4668 r0 *1 28.905,24.57
X$4668 147 19 148 644 645 cell_1rw
* cell instance $4669 r0 *1 29.61,24.57
X$4669 149 19 150 644 645 cell_1rw
* cell instance $4670 r0 *1 30.315,24.57
X$4670 151 19 152 644 645 cell_1rw
* cell instance $4671 r0 *1 31.02,24.57
X$4671 153 19 154 644 645 cell_1rw
* cell instance $4672 r0 *1 31.725,24.57
X$4672 155 19 156 644 645 cell_1rw
* cell instance $4673 r0 *1 32.43,24.57
X$4673 157 19 158 644 645 cell_1rw
* cell instance $4674 r0 *1 33.135,24.57
X$4674 159 19 160 644 645 cell_1rw
* cell instance $4675 r0 *1 33.84,24.57
X$4675 161 19 162 644 645 cell_1rw
* cell instance $4676 r0 *1 34.545,24.57
X$4676 163 19 164 644 645 cell_1rw
* cell instance $4677 r0 *1 35.25,24.57
X$4677 165 19 166 644 645 cell_1rw
* cell instance $4678 r0 *1 35.955,24.57
X$4678 167 19 168 644 645 cell_1rw
* cell instance $4679 r0 *1 36.66,24.57
X$4679 169 19 170 644 645 cell_1rw
* cell instance $4680 r0 *1 37.365,24.57
X$4680 171 19 172 644 645 cell_1rw
* cell instance $4681 r0 *1 38.07,24.57
X$4681 173 19 174 644 645 cell_1rw
* cell instance $4682 r0 *1 38.775,24.57
X$4682 175 19 176 644 645 cell_1rw
* cell instance $4683 r0 *1 39.48,24.57
X$4683 177 19 178 644 645 cell_1rw
* cell instance $4684 r0 *1 40.185,24.57
X$4684 179 19 180 644 645 cell_1rw
* cell instance $4685 r0 *1 40.89,24.57
X$4685 181 19 182 644 645 cell_1rw
* cell instance $4686 r0 *1 41.595,24.57
X$4686 183 19 184 644 645 cell_1rw
* cell instance $4687 r0 *1 42.3,24.57
X$4687 185 19 186 644 645 cell_1rw
* cell instance $4688 r0 *1 43.005,24.57
X$4688 187 19 188 644 645 cell_1rw
* cell instance $4689 r0 *1 43.71,24.57
X$4689 189 19 190 644 645 cell_1rw
* cell instance $4690 r0 *1 44.415,24.57
X$4690 191 19 192 644 645 cell_1rw
* cell instance $4691 r0 *1 45.12,24.57
X$4691 193 19 194 644 645 cell_1rw
* cell instance $4692 r0 *1 45.825,24.57
X$4692 195 19 196 644 645 cell_1rw
* cell instance $4693 r0 *1 46.53,24.57
X$4693 197 19 198 644 645 cell_1rw
* cell instance $4694 r0 *1 47.235,24.57
X$4694 199 19 200 644 645 cell_1rw
* cell instance $4695 r0 *1 47.94,24.57
X$4695 201 19 202 644 645 cell_1rw
* cell instance $4696 r0 *1 48.645,24.57
X$4696 203 19 204 644 645 cell_1rw
* cell instance $4697 r0 *1 49.35,24.57
X$4697 205 19 206 644 645 cell_1rw
* cell instance $4698 r0 *1 50.055,24.57
X$4698 207 19 208 644 645 cell_1rw
* cell instance $4699 r0 *1 50.76,24.57
X$4699 209 19 210 644 645 cell_1rw
* cell instance $4700 r0 *1 51.465,24.57
X$4700 211 19 212 644 645 cell_1rw
* cell instance $4701 r0 *1 52.17,24.57
X$4701 213 19 214 644 645 cell_1rw
* cell instance $4702 r0 *1 52.875,24.57
X$4702 215 19 216 644 645 cell_1rw
* cell instance $4703 r0 *1 53.58,24.57
X$4703 217 19 218 644 645 cell_1rw
* cell instance $4704 r0 *1 54.285,24.57
X$4704 219 19 220 644 645 cell_1rw
* cell instance $4705 r0 *1 54.99,24.57
X$4705 221 19 222 644 645 cell_1rw
* cell instance $4706 r0 *1 55.695,24.57
X$4706 223 19 224 644 645 cell_1rw
* cell instance $4707 r0 *1 56.4,24.57
X$4707 225 19 226 644 645 cell_1rw
* cell instance $4708 r0 *1 57.105,24.57
X$4708 227 19 228 644 645 cell_1rw
* cell instance $4709 r0 *1 57.81,24.57
X$4709 229 19 230 644 645 cell_1rw
* cell instance $4710 r0 *1 58.515,24.57
X$4710 231 19 232 644 645 cell_1rw
* cell instance $4711 r0 *1 59.22,24.57
X$4711 233 19 234 644 645 cell_1rw
* cell instance $4712 r0 *1 59.925,24.57
X$4712 235 19 236 644 645 cell_1rw
* cell instance $4713 r0 *1 60.63,24.57
X$4713 237 19 238 644 645 cell_1rw
* cell instance $4714 r0 *1 61.335,24.57
X$4714 239 19 240 644 645 cell_1rw
* cell instance $4715 r0 *1 62.04,24.57
X$4715 241 19 242 644 645 cell_1rw
* cell instance $4716 r0 *1 62.745,24.57
X$4716 243 19 244 644 645 cell_1rw
* cell instance $4717 r0 *1 63.45,24.57
X$4717 245 19 246 644 645 cell_1rw
* cell instance $4718 r0 *1 64.155,24.57
X$4718 247 19 248 644 645 cell_1rw
* cell instance $4719 r0 *1 64.86,24.57
X$4719 249 19 250 644 645 cell_1rw
* cell instance $4720 r0 *1 65.565,24.57
X$4720 251 19 252 644 645 cell_1rw
* cell instance $4721 r0 *1 66.27,24.57
X$4721 253 19 254 644 645 cell_1rw
* cell instance $4722 r0 *1 66.975,24.57
X$4722 255 19 256 644 645 cell_1rw
* cell instance $4723 r0 *1 67.68,24.57
X$4723 257 19 258 644 645 cell_1rw
* cell instance $4724 r0 *1 68.385,24.57
X$4724 259 19 260 644 645 cell_1rw
* cell instance $4725 r0 *1 69.09,24.57
X$4725 261 19 262 644 645 cell_1rw
* cell instance $4726 r0 *1 69.795,24.57
X$4726 263 19 264 644 645 cell_1rw
* cell instance $4727 r0 *1 70.5,24.57
X$4727 265 19 266 644 645 cell_1rw
* cell instance $4728 r0 *1 71.205,24.57
X$4728 267 19 268 644 645 cell_1rw
* cell instance $4729 r0 *1 71.91,24.57
X$4729 269 19 270 644 645 cell_1rw
* cell instance $4730 r0 *1 72.615,24.57
X$4730 271 19 272 644 645 cell_1rw
* cell instance $4731 r0 *1 73.32,24.57
X$4731 273 19 274 644 645 cell_1rw
* cell instance $4732 r0 *1 74.025,24.57
X$4732 275 19 276 644 645 cell_1rw
* cell instance $4733 r0 *1 74.73,24.57
X$4733 277 19 278 644 645 cell_1rw
* cell instance $4734 r0 *1 75.435,24.57
X$4734 279 19 280 644 645 cell_1rw
* cell instance $4735 r0 *1 76.14,24.57
X$4735 281 19 282 644 645 cell_1rw
* cell instance $4736 r0 *1 76.845,24.57
X$4736 283 19 284 644 645 cell_1rw
* cell instance $4737 r0 *1 77.55,24.57
X$4737 285 19 286 644 645 cell_1rw
* cell instance $4738 r0 *1 78.255,24.57
X$4738 287 19 288 644 645 cell_1rw
* cell instance $4739 r0 *1 78.96,24.57
X$4739 289 19 290 644 645 cell_1rw
* cell instance $4740 r0 *1 79.665,24.57
X$4740 291 19 292 644 645 cell_1rw
* cell instance $4741 r0 *1 80.37,24.57
X$4741 293 19 294 644 645 cell_1rw
* cell instance $4742 r0 *1 81.075,24.57
X$4742 295 19 296 644 645 cell_1rw
* cell instance $4743 r0 *1 81.78,24.57
X$4743 297 19 298 644 645 cell_1rw
* cell instance $4744 r0 *1 82.485,24.57
X$4744 299 19 300 644 645 cell_1rw
* cell instance $4745 r0 *1 83.19,24.57
X$4745 301 19 302 644 645 cell_1rw
* cell instance $4746 r0 *1 83.895,24.57
X$4746 303 19 304 644 645 cell_1rw
* cell instance $4747 r0 *1 84.6,24.57
X$4747 305 19 306 644 645 cell_1rw
* cell instance $4748 r0 *1 85.305,24.57
X$4748 307 19 308 644 645 cell_1rw
* cell instance $4749 r0 *1 86.01,24.57
X$4749 309 19 310 644 645 cell_1rw
* cell instance $4750 r0 *1 86.715,24.57
X$4750 311 19 312 644 645 cell_1rw
* cell instance $4751 r0 *1 87.42,24.57
X$4751 313 19 314 644 645 cell_1rw
* cell instance $4752 r0 *1 88.125,24.57
X$4752 315 19 316 644 645 cell_1rw
* cell instance $4753 r0 *1 88.83,24.57
X$4753 317 19 318 644 645 cell_1rw
* cell instance $4754 r0 *1 89.535,24.57
X$4754 319 19 320 644 645 cell_1rw
* cell instance $4755 r0 *1 90.24,24.57
X$4755 321 19 323 644 645 cell_1rw
* cell instance $4756 r0 *1 90.945,24.57
X$4756 324 19 325 644 645 cell_1rw
* cell instance $4757 r0 *1 91.65,24.57
X$4757 326 19 327 644 645 cell_1rw
* cell instance $4758 r0 *1 92.355,24.57
X$4758 328 19 329 644 645 cell_1rw
* cell instance $4759 r0 *1 93.06,24.57
X$4759 330 19 331 644 645 cell_1rw
* cell instance $4760 r0 *1 93.765,24.57
X$4760 332 19 333 644 645 cell_1rw
* cell instance $4761 r0 *1 94.47,24.57
X$4761 334 19 335 644 645 cell_1rw
* cell instance $4762 r0 *1 95.175,24.57
X$4762 336 19 337 644 645 cell_1rw
* cell instance $4763 r0 *1 95.88,24.57
X$4763 338 19 339 644 645 cell_1rw
* cell instance $4764 r0 *1 96.585,24.57
X$4764 340 19 341 644 645 cell_1rw
* cell instance $4765 r0 *1 97.29,24.57
X$4765 342 19 343 644 645 cell_1rw
* cell instance $4766 r0 *1 97.995,24.57
X$4766 344 19 345 644 645 cell_1rw
* cell instance $4767 r0 *1 98.7,24.57
X$4767 346 19 347 644 645 cell_1rw
* cell instance $4768 r0 *1 99.405,24.57
X$4768 348 19 349 644 645 cell_1rw
* cell instance $4769 r0 *1 100.11,24.57
X$4769 350 19 351 644 645 cell_1rw
* cell instance $4770 r0 *1 100.815,24.57
X$4770 352 19 353 644 645 cell_1rw
* cell instance $4771 r0 *1 101.52,24.57
X$4771 354 19 355 644 645 cell_1rw
* cell instance $4772 r0 *1 102.225,24.57
X$4772 356 19 357 644 645 cell_1rw
* cell instance $4773 r0 *1 102.93,24.57
X$4773 358 19 359 644 645 cell_1rw
* cell instance $4774 r0 *1 103.635,24.57
X$4774 360 19 361 644 645 cell_1rw
* cell instance $4775 r0 *1 104.34,24.57
X$4775 362 19 363 644 645 cell_1rw
* cell instance $4776 r0 *1 105.045,24.57
X$4776 364 19 365 644 645 cell_1rw
* cell instance $4777 r0 *1 105.75,24.57
X$4777 366 19 367 644 645 cell_1rw
* cell instance $4778 r0 *1 106.455,24.57
X$4778 368 19 369 644 645 cell_1rw
* cell instance $4779 r0 *1 107.16,24.57
X$4779 370 19 371 644 645 cell_1rw
* cell instance $4780 r0 *1 107.865,24.57
X$4780 372 19 373 644 645 cell_1rw
* cell instance $4781 r0 *1 108.57,24.57
X$4781 374 19 375 644 645 cell_1rw
* cell instance $4782 r0 *1 109.275,24.57
X$4782 376 19 377 644 645 cell_1rw
* cell instance $4783 r0 *1 109.98,24.57
X$4783 378 19 379 644 645 cell_1rw
* cell instance $4784 r0 *1 110.685,24.57
X$4784 380 19 381 644 645 cell_1rw
* cell instance $4785 r0 *1 111.39,24.57
X$4785 382 19 383 644 645 cell_1rw
* cell instance $4786 r0 *1 112.095,24.57
X$4786 384 19 385 644 645 cell_1rw
* cell instance $4787 r0 *1 112.8,24.57
X$4787 386 19 387 644 645 cell_1rw
* cell instance $4788 r0 *1 113.505,24.57
X$4788 388 19 389 644 645 cell_1rw
* cell instance $4789 r0 *1 114.21,24.57
X$4789 390 19 391 644 645 cell_1rw
* cell instance $4790 r0 *1 114.915,24.57
X$4790 392 19 393 644 645 cell_1rw
* cell instance $4791 r0 *1 115.62,24.57
X$4791 394 19 395 644 645 cell_1rw
* cell instance $4792 r0 *1 116.325,24.57
X$4792 396 19 397 644 645 cell_1rw
* cell instance $4793 r0 *1 117.03,24.57
X$4793 398 19 399 644 645 cell_1rw
* cell instance $4794 r0 *1 117.735,24.57
X$4794 400 19 401 644 645 cell_1rw
* cell instance $4795 r0 *1 118.44,24.57
X$4795 402 19 403 644 645 cell_1rw
* cell instance $4796 r0 *1 119.145,24.57
X$4796 404 19 405 644 645 cell_1rw
* cell instance $4797 r0 *1 119.85,24.57
X$4797 406 19 407 644 645 cell_1rw
* cell instance $4798 r0 *1 120.555,24.57
X$4798 408 19 409 644 645 cell_1rw
* cell instance $4799 r0 *1 121.26,24.57
X$4799 410 19 411 644 645 cell_1rw
* cell instance $4800 r0 *1 121.965,24.57
X$4800 412 19 413 644 645 cell_1rw
* cell instance $4801 r0 *1 122.67,24.57
X$4801 414 19 415 644 645 cell_1rw
* cell instance $4802 r0 *1 123.375,24.57
X$4802 416 19 417 644 645 cell_1rw
* cell instance $4803 r0 *1 124.08,24.57
X$4803 418 19 419 644 645 cell_1rw
* cell instance $4804 r0 *1 124.785,24.57
X$4804 420 19 421 644 645 cell_1rw
* cell instance $4805 r0 *1 125.49,24.57
X$4805 422 19 423 644 645 cell_1rw
* cell instance $4806 r0 *1 126.195,24.57
X$4806 424 19 425 644 645 cell_1rw
* cell instance $4807 r0 *1 126.9,24.57
X$4807 426 19 427 644 645 cell_1rw
* cell instance $4808 r0 *1 127.605,24.57
X$4808 428 19 429 644 645 cell_1rw
* cell instance $4809 r0 *1 128.31,24.57
X$4809 430 19 431 644 645 cell_1rw
* cell instance $4810 r0 *1 129.015,24.57
X$4810 432 19 433 644 645 cell_1rw
* cell instance $4811 r0 *1 129.72,24.57
X$4811 434 19 435 644 645 cell_1rw
* cell instance $4812 r0 *1 130.425,24.57
X$4812 436 19 437 644 645 cell_1rw
* cell instance $4813 r0 *1 131.13,24.57
X$4813 438 19 439 644 645 cell_1rw
* cell instance $4814 r0 *1 131.835,24.57
X$4814 440 19 441 644 645 cell_1rw
* cell instance $4815 r0 *1 132.54,24.57
X$4815 442 19 443 644 645 cell_1rw
* cell instance $4816 r0 *1 133.245,24.57
X$4816 444 19 445 644 645 cell_1rw
* cell instance $4817 r0 *1 133.95,24.57
X$4817 446 19 447 644 645 cell_1rw
* cell instance $4818 r0 *1 134.655,24.57
X$4818 448 19 449 644 645 cell_1rw
* cell instance $4819 r0 *1 135.36,24.57
X$4819 450 19 451 644 645 cell_1rw
* cell instance $4820 r0 *1 136.065,24.57
X$4820 452 19 453 644 645 cell_1rw
* cell instance $4821 r0 *1 136.77,24.57
X$4821 454 19 455 644 645 cell_1rw
* cell instance $4822 r0 *1 137.475,24.57
X$4822 456 19 457 644 645 cell_1rw
* cell instance $4823 r0 *1 138.18,24.57
X$4823 458 19 459 644 645 cell_1rw
* cell instance $4824 r0 *1 138.885,24.57
X$4824 460 19 461 644 645 cell_1rw
* cell instance $4825 r0 *1 139.59,24.57
X$4825 462 19 463 644 645 cell_1rw
* cell instance $4826 r0 *1 140.295,24.57
X$4826 464 19 465 644 645 cell_1rw
* cell instance $4827 r0 *1 141,24.57
X$4827 466 19 467 644 645 cell_1rw
* cell instance $4828 r0 *1 141.705,24.57
X$4828 468 19 469 644 645 cell_1rw
* cell instance $4829 r0 *1 142.41,24.57
X$4829 470 19 471 644 645 cell_1rw
* cell instance $4830 r0 *1 143.115,24.57
X$4830 472 19 473 644 645 cell_1rw
* cell instance $4831 r0 *1 143.82,24.57
X$4831 474 19 475 644 645 cell_1rw
* cell instance $4832 r0 *1 144.525,24.57
X$4832 476 19 477 644 645 cell_1rw
* cell instance $4833 r0 *1 145.23,24.57
X$4833 478 19 479 644 645 cell_1rw
* cell instance $4834 r0 *1 145.935,24.57
X$4834 480 19 481 644 645 cell_1rw
* cell instance $4835 r0 *1 146.64,24.57
X$4835 482 19 483 644 645 cell_1rw
* cell instance $4836 r0 *1 147.345,24.57
X$4836 484 19 485 644 645 cell_1rw
* cell instance $4837 r0 *1 148.05,24.57
X$4837 486 19 487 644 645 cell_1rw
* cell instance $4838 r0 *1 148.755,24.57
X$4838 488 19 489 644 645 cell_1rw
* cell instance $4839 r0 *1 149.46,24.57
X$4839 490 19 491 644 645 cell_1rw
* cell instance $4840 r0 *1 150.165,24.57
X$4840 492 19 493 644 645 cell_1rw
* cell instance $4841 r0 *1 150.87,24.57
X$4841 494 19 495 644 645 cell_1rw
* cell instance $4842 r0 *1 151.575,24.57
X$4842 496 19 497 644 645 cell_1rw
* cell instance $4843 r0 *1 152.28,24.57
X$4843 498 19 499 644 645 cell_1rw
* cell instance $4844 r0 *1 152.985,24.57
X$4844 500 19 501 644 645 cell_1rw
* cell instance $4845 r0 *1 153.69,24.57
X$4845 502 19 503 644 645 cell_1rw
* cell instance $4846 r0 *1 154.395,24.57
X$4846 504 19 505 644 645 cell_1rw
* cell instance $4847 r0 *1 155.1,24.57
X$4847 506 19 507 644 645 cell_1rw
* cell instance $4848 r0 *1 155.805,24.57
X$4848 508 19 509 644 645 cell_1rw
* cell instance $4849 r0 *1 156.51,24.57
X$4849 510 19 511 644 645 cell_1rw
* cell instance $4850 r0 *1 157.215,24.57
X$4850 512 19 513 644 645 cell_1rw
* cell instance $4851 r0 *1 157.92,24.57
X$4851 514 19 515 644 645 cell_1rw
* cell instance $4852 r0 *1 158.625,24.57
X$4852 516 19 517 644 645 cell_1rw
* cell instance $4853 r0 *1 159.33,24.57
X$4853 518 19 519 644 645 cell_1rw
* cell instance $4854 r0 *1 160.035,24.57
X$4854 520 19 521 644 645 cell_1rw
* cell instance $4855 r0 *1 160.74,24.57
X$4855 522 19 523 644 645 cell_1rw
* cell instance $4856 r0 *1 161.445,24.57
X$4856 524 19 525 644 645 cell_1rw
* cell instance $4857 r0 *1 162.15,24.57
X$4857 526 19 527 644 645 cell_1rw
* cell instance $4858 r0 *1 162.855,24.57
X$4858 528 19 529 644 645 cell_1rw
* cell instance $4859 r0 *1 163.56,24.57
X$4859 530 19 531 644 645 cell_1rw
* cell instance $4860 r0 *1 164.265,24.57
X$4860 532 19 533 644 645 cell_1rw
* cell instance $4861 r0 *1 164.97,24.57
X$4861 534 19 535 644 645 cell_1rw
* cell instance $4862 r0 *1 165.675,24.57
X$4862 536 19 537 644 645 cell_1rw
* cell instance $4863 r0 *1 166.38,24.57
X$4863 538 19 539 644 645 cell_1rw
* cell instance $4864 r0 *1 167.085,24.57
X$4864 540 19 541 644 645 cell_1rw
* cell instance $4865 r0 *1 167.79,24.57
X$4865 542 19 543 644 645 cell_1rw
* cell instance $4866 r0 *1 168.495,24.57
X$4866 544 19 545 644 645 cell_1rw
* cell instance $4867 r0 *1 169.2,24.57
X$4867 546 19 547 644 645 cell_1rw
* cell instance $4868 r0 *1 169.905,24.57
X$4868 548 19 549 644 645 cell_1rw
* cell instance $4869 r0 *1 170.61,24.57
X$4869 550 19 551 644 645 cell_1rw
* cell instance $4870 r0 *1 171.315,24.57
X$4870 552 19 553 644 645 cell_1rw
* cell instance $4871 r0 *1 172.02,24.57
X$4871 554 19 555 644 645 cell_1rw
* cell instance $4872 r0 *1 172.725,24.57
X$4872 556 19 557 644 645 cell_1rw
* cell instance $4873 r0 *1 173.43,24.57
X$4873 558 19 559 644 645 cell_1rw
* cell instance $4874 r0 *1 174.135,24.57
X$4874 560 19 561 644 645 cell_1rw
* cell instance $4875 r0 *1 174.84,24.57
X$4875 562 19 563 644 645 cell_1rw
* cell instance $4876 r0 *1 175.545,24.57
X$4876 564 19 565 644 645 cell_1rw
* cell instance $4877 r0 *1 176.25,24.57
X$4877 566 19 567 644 645 cell_1rw
* cell instance $4878 r0 *1 176.955,24.57
X$4878 568 19 569 644 645 cell_1rw
* cell instance $4879 r0 *1 177.66,24.57
X$4879 570 19 571 644 645 cell_1rw
* cell instance $4880 r0 *1 178.365,24.57
X$4880 572 19 573 644 645 cell_1rw
* cell instance $4881 r0 *1 179.07,24.57
X$4881 574 19 575 644 645 cell_1rw
* cell instance $4882 r0 *1 179.775,24.57
X$4882 576 19 577 644 645 cell_1rw
* cell instance $4883 r0 *1 180.48,24.57
X$4883 578 19 579 644 645 cell_1rw
* cell instance $4884 m0 *1 0.705,27.3
X$4884 67 20 68 644 645 cell_1rw
* cell instance $4885 m0 *1 0,27.3
X$4885 65 20 66 644 645 cell_1rw
* cell instance $4886 m0 *1 1.41,27.3
X$4886 69 20 70 644 645 cell_1rw
* cell instance $4887 m0 *1 2.115,27.3
X$4887 71 20 72 644 645 cell_1rw
* cell instance $4888 m0 *1 2.82,27.3
X$4888 73 20 74 644 645 cell_1rw
* cell instance $4889 m0 *1 3.525,27.3
X$4889 75 20 76 644 645 cell_1rw
* cell instance $4890 m0 *1 4.23,27.3
X$4890 77 20 78 644 645 cell_1rw
* cell instance $4891 m0 *1 4.935,27.3
X$4891 79 20 80 644 645 cell_1rw
* cell instance $4892 m0 *1 5.64,27.3
X$4892 81 20 82 644 645 cell_1rw
* cell instance $4893 m0 *1 6.345,27.3
X$4893 83 20 84 644 645 cell_1rw
* cell instance $4894 m0 *1 7.05,27.3
X$4894 85 20 86 644 645 cell_1rw
* cell instance $4895 m0 *1 7.755,27.3
X$4895 87 20 88 644 645 cell_1rw
* cell instance $4896 m0 *1 8.46,27.3
X$4896 89 20 90 644 645 cell_1rw
* cell instance $4897 m0 *1 9.165,27.3
X$4897 91 20 92 644 645 cell_1rw
* cell instance $4898 m0 *1 9.87,27.3
X$4898 93 20 94 644 645 cell_1rw
* cell instance $4899 m0 *1 10.575,27.3
X$4899 95 20 96 644 645 cell_1rw
* cell instance $4900 m0 *1 11.28,27.3
X$4900 97 20 98 644 645 cell_1rw
* cell instance $4901 m0 *1 11.985,27.3
X$4901 99 20 100 644 645 cell_1rw
* cell instance $4902 m0 *1 12.69,27.3
X$4902 101 20 102 644 645 cell_1rw
* cell instance $4903 m0 *1 13.395,27.3
X$4903 103 20 104 644 645 cell_1rw
* cell instance $4904 m0 *1 14.1,27.3
X$4904 105 20 106 644 645 cell_1rw
* cell instance $4905 m0 *1 14.805,27.3
X$4905 107 20 108 644 645 cell_1rw
* cell instance $4906 m0 *1 15.51,27.3
X$4906 109 20 110 644 645 cell_1rw
* cell instance $4907 m0 *1 16.215,27.3
X$4907 111 20 112 644 645 cell_1rw
* cell instance $4908 m0 *1 16.92,27.3
X$4908 113 20 114 644 645 cell_1rw
* cell instance $4909 m0 *1 17.625,27.3
X$4909 115 20 116 644 645 cell_1rw
* cell instance $4910 m0 *1 18.33,27.3
X$4910 117 20 118 644 645 cell_1rw
* cell instance $4911 m0 *1 19.035,27.3
X$4911 119 20 120 644 645 cell_1rw
* cell instance $4912 m0 *1 19.74,27.3
X$4912 121 20 122 644 645 cell_1rw
* cell instance $4913 m0 *1 20.445,27.3
X$4913 123 20 124 644 645 cell_1rw
* cell instance $4914 m0 *1 21.15,27.3
X$4914 125 20 126 644 645 cell_1rw
* cell instance $4915 m0 *1 21.855,27.3
X$4915 127 20 128 644 645 cell_1rw
* cell instance $4916 m0 *1 22.56,27.3
X$4916 129 20 130 644 645 cell_1rw
* cell instance $4917 m0 *1 23.265,27.3
X$4917 131 20 132 644 645 cell_1rw
* cell instance $4918 m0 *1 23.97,27.3
X$4918 133 20 134 644 645 cell_1rw
* cell instance $4919 m0 *1 24.675,27.3
X$4919 135 20 136 644 645 cell_1rw
* cell instance $4920 m0 *1 25.38,27.3
X$4920 137 20 138 644 645 cell_1rw
* cell instance $4921 m0 *1 26.085,27.3
X$4921 139 20 140 644 645 cell_1rw
* cell instance $4922 m0 *1 26.79,27.3
X$4922 141 20 142 644 645 cell_1rw
* cell instance $4923 m0 *1 27.495,27.3
X$4923 143 20 144 644 645 cell_1rw
* cell instance $4924 m0 *1 28.2,27.3
X$4924 145 20 146 644 645 cell_1rw
* cell instance $4925 m0 *1 28.905,27.3
X$4925 147 20 148 644 645 cell_1rw
* cell instance $4926 m0 *1 29.61,27.3
X$4926 149 20 150 644 645 cell_1rw
* cell instance $4927 m0 *1 30.315,27.3
X$4927 151 20 152 644 645 cell_1rw
* cell instance $4928 m0 *1 31.02,27.3
X$4928 153 20 154 644 645 cell_1rw
* cell instance $4929 m0 *1 31.725,27.3
X$4929 155 20 156 644 645 cell_1rw
* cell instance $4930 m0 *1 32.43,27.3
X$4930 157 20 158 644 645 cell_1rw
* cell instance $4931 m0 *1 33.135,27.3
X$4931 159 20 160 644 645 cell_1rw
* cell instance $4932 m0 *1 33.84,27.3
X$4932 161 20 162 644 645 cell_1rw
* cell instance $4933 m0 *1 34.545,27.3
X$4933 163 20 164 644 645 cell_1rw
* cell instance $4934 m0 *1 35.25,27.3
X$4934 165 20 166 644 645 cell_1rw
* cell instance $4935 m0 *1 35.955,27.3
X$4935 167 20 168 644 645 cell_1rw
* cell instance $4936 m0 *1 36.66,27.3
X$4936 169 20 170 644 645 cell_1rw
* cell instance $4937 m0 *1 37.365,27.3
X$4937 171 20 172 644 645 cell_1rw
* cell instance $4938 m0 *1 38.07,27.3
X$4938 173 20 174 644 645 cell_1rw
* cell instance $4939 m0 *1 38.775,27.3
X$4939 175 20 176 644 645 cell_1rw
* cell instance $4940 m0 *1 39.48,27.3
X$4940 177 20 178 644 645 cell_1rw
* cell instance $4941 m0 *1 40.185,27.3
X$4941 179 20 180 644 645 cell_1rw
* cell instance $4942 m0 *1 40.89,27.3
X$4942 181 20 182 644 645 cell_1rw
* cell instance $4943 m0 *1 41.595,27.3
X$4943 183 20 184 644 645 cell_1rw
* cell instance $4944 m0 *1 42.3,27.3
X$4944 185 20 186 644 645 cell_1rw
* cell instance $4945 m0 *1 43.005,27.3
X$4945 187 20 188 644 645 cell_1rw
* cell instance $4946 m0 *1 43.71,27.3
X$4946 189 20 190 644 645 cell_1rw
* cell instance $4947 m0 *1 44.415,27.3
X$4947 191 20 192 644 645 cell_1rw
* cell instance $4948 m0 *1 45.12,27.3
X$4948 193 20 194 644 645 cell_1rw
* cell instance $4949 m0 *1 45.825,27.3
X$4949 195 20 196 644 645 cell_1rw
* cell instance $4950 m0 *1 46.53,27.3
X$4950 197 20 198 644 645 cell_1rw
* cell instance $4951 m0 *1 47.235,27.3
X$4951 199 20 200 644 645 cell_1rw
* cell instance $4952 m0 *1 47.94,27.3
X$4952 201 20 202 644 645 cell_1rw
* cell instance $4953 m0 *1 48.645,27.3
X$4953 203 20 204 644 645 cell_1rw
* cell instance $4954 m0 *1 49.35,27.3
X$4954 205 20 206 644 645 cell_1rw
* cell instance $4955 m0 *1 50.055,27.3
X$4955 207 20 208 644 645 cell_1rw
* cell instance $4956 m0 *1 50.76,27.3
X$4956 209 20 210 644 645 cell_1rw
* cell instance $4957 m0 *1 51.465,27.3
X$4957 211 20 212 644 645 cell_1rw
* cell instance $4958 m0 *1 52.17,27.3
X$4958 213 20 214 644 645 cell_1rw
* cell instance $4959 m0 *1 52.875,27.3
X$4959 215 20 216 644 645 cell_1rw
* cell instance $4960 m0 *1 53.58,27.3
X$4960 217 20 218 644 645 cell_1rw
* cell instance $4961 m0 *1 54.285,27.3
X$4961 219 20 220 644 645 cell_1rw
* cell instance $4962 m0 *1 54.99,27.3
X$4962 221 20 222 644 645 cell_1rw
* cell instance $4963 m0 *1 55.695,27.3
X$4963 223 20 224 644 645 cell_1rw
* cell instance $4964 m0 *1 56.4,27.3
X$4964 225 20 226 644 645 cell_1rw
* cell instance $4965 m0 *1 57.105,27.3
X$4965 227 20 228 644 645 cell_1rw
* cell instance $4966 m0 *1 57.81,27.3
X$4966 229 20 230 644 645 cell_1rw
* cell instance $4967 m0 *1 58.515,27.3
X$4967 231 20 232 644 645 cell_1rw
* cell instance $4968 m0 *1 59.22,27.3
X$4968 233 20 234 644 645 cell_1rw
* cell instance $4969 m0 *1 59.925,27.3
X$4969 235 20 236 644 645 cell_1rw
* cell instance $4970 m0 *1 60.63,27.3
X$4970 237 20 238 644 645 cell_1rw
* cell instance $4971 m0 *1 61.335,27.3
X$4971 239 20 240 644 645 cell_1rw
* cell instance $4972 m0 *1 62.04,27.3
X$4972 241 20 242 644 645 cell_1rw
* cell instance $4973 m0 *1 62.745,27.3
X$4973 243 20 244 644 645 cell_1rw
* cell instance $4974 m0 *1 63.45,27.3
X$4974 245 20 246 644 645 cell_1rw
* cell instance $4975 m0 *1 64.155,27.3
X$4975 247 20 248 644 645 cell_1rw
* cell instance $4976 m0 *1 64.86,27.3
X$4976 249 20 250 644 645 cell_1rw
* cell instance $4977 m0 *1 65.565,27.3
X$4977 251 20 252 644 645 cell_1rw
* cell instance $4978 m0 *1 66.27,27.3
X$4978 253 20 254 644 645 cell_1rw
* cell instance $4979 m0 *1 66.975,27.3
X$4979 255 20 256 644 645 cell_1rw
* cell instance $4980 m0 *1 67.68,27.3
X$4980 257 20 258 644 645 cell_1rw
* cell instance $4981 m0 *1 68.385,27.3
X$4981 259 20 260 644 645 cell_1rw
* cell instance $4982 m0 *1 69.09,27.3
X$4982 261 20 262 644 645 cell_1rw
* cell instance $4983 m0 *1 69.795,27.3
X$4983 263 20 264 644 645 cell_1rw
* cell instance $4984 m0 *1 70.5,27.3
X$4984 265 20 266 644 645 cell_1rw
* cell instance $4985 m0 *1 71.205,27.3
X$4985 267 20 268 644 645 cell_1rw
* cell instance $4986 m0 *1 71.91,27.3
X$4986 269 20 270 644 645 cell_1rw
* cell instance $4987 m0 *1 72.615,27.3
X$4987 271 20 272 644 645 cell_1rw
* cell instance $4988 m0 *1 73.32,27.3
X$4988 273 20 274 644 645 cell_1rw
* cell instance $4989 m0 *1 74.025,27.3
X$4989 275 20 276 644 645 cell_1rw
* cell instance $4990 m0 *1 74.73,27.3
X$4990 277 20 278 644 645 cell_1rw
* cell instance $4991 m0 *1 75.435,27.3
X$4991 279 20 280 644 645 cell_1rw
* cell instance $4992 m0 *1 76.14,27.3
X$4992 281 20 282 644 645 cell_1rw
* cell instance $4993 m0 *1 76.845,27.3
X$4993 283 20 284 644 645 cell_1rw
* cell instance $4994 m0 *1 77.55,27.3
X$4994 285 20 286 644 645 cell_1rw
* cell instance $4995 m0 *1 78.255,27.3
X$4995 287 20 288 644 645 cell_1rw
* cell instance $4996 m0 *1 78.96,27.3
X$4996 289 20 290 644 645 cell_1rw
* cell instance $4997 m0 *1 79.665,27.3
X$4997 291 20 292 644 645 cell_1rw
* cell instance $4998 m0 *1 80.37,27.3
X$4998 293 20 294 644 645 cell_1rw
* cell instance $4999 m0 *1 81.075,27.3
X$4999 295 20 296 644 645 cell_1rw
* cell instance $5000 m0 *1 81.78,27.3
X$5000 297 20 298 644 645 cell_1rw
* cell instance $5001 m0 *1 82.485,27.3
X$5001 299 20 300 644 645 cell_1rw
* cell instance $5002 m0 *1 83.19,27.3
X$5002 301 20 302 644 645 cell_1rw
* cell instance $5003 m0 *1 83.895,27.3
X$5003 303 20 304 644 645 cell_1rw
* cell instance $5004 m0 *1 84.6,27.3
X$5004 305 20 306 644 645 cell_1rw
* cell instance $5005 m0 *1 85.305,27.3
X$5005 307 20 308 644 645 cell_1rw
* cell instance $5006 m0 *1 86.01,27.3
X$5006 309 20 310 644 645 cell_1rw
* cell instance $5007 m0 *1 86.715,27.3
X$5007 311 20 312 644 645 cell_1rw
* cell instance $5008 m0 *1 87.42,27.3
X$5008 313 20 314 644 645 cell_1rw
* cell instance $5009 m0 *1 88.125,27.3
X$5009 315 20 316 644 645 cell_1rw
* cell instance $5010 m0 *1 88.83,27.3
X$5010 317 20 318 644 645 cell_1rw
* cell instance $5011 m0 *1 89.535,27.3
X$5011 319 20 320 644 645 cell_1rw
* cell instance $5012 m0 *1 90.24,27.3
X$5012 321 20 323 644 645 cell_1rw
* cell instance $5013 m0 *1 90.945,27.3
X$5013 324 20 325 644 645 cell_1rw
* cell instance $5014 m0 *1 91.65,27.3
X$5014 326 20 327 644 645 cell_1rw
* cell instance $5015 m0 *1 92.355,27.3
X$5015 328 20 329 644 645 cell_1rw
* cell instance $5016 m0 *1 93.06,27.3
X$5016 330 20 331 644 645 cell_1rw
* cell instance $5017 m0 *1 93.765,27.3
X$5017 332 20 333 644 645 cell_1rw
* cell instance $5018 m0 *1 94.47,27.3
X$5018 334 20 335 644 645 cell_1rw
* cell instance $5019 m0 *1 95.175,27.3
X$5019 336 20 337 644 645 cell_1rw
* cell instance $5020 m0 *1 95.88,27.3
X$5020 338 20 339 644 645 cell_1rw
* cell instance $5021 m0 *1 96.585,27.3
X$5021 340 20 341 644 645 cell_1rw
* cell instance $5022 m0 *1 97.29,27.3
X$5022 342 20 343 644 645 cell_1rw
* cell instance $5023 m0 *1 97.995,27.3
X$5023 344 20 345 644 645 cell_1rw
* cell instance $5024 m0 *1 98.7,27.3
X$5024 346 20 347 644 645 cell_1rw
* cell instance $5025 m0 *1 99.405,27.3
X$5025 348 20 349 644 645 cell_1rw
* cell instance $5026 m0 *1 100.11,27.3
X$5026 350 20 351 644 645 cell_1rw
* cell instance $5027 m0 *1 100.815,27.3
X$5027 352 20 353 644 645 cell_1rw
* cell instance $5028 m0 *1 101.52,27.3
X$5028 354 20 355 644 645 cell_1rw
* cell instance $5029 m0 *1 102.225,27.3
X$5029 356 20 357 644 645 cell_1rw
* cell instance $5030 m0 *1 102.93,27.3
X$5030 358 20 359 644 645 cell_1rw
* cell instance $5031 m0 *1 103.635,27.3
X$5031 360 20 361 644 645 cell_1rw
* cell instance $5032 m0 *1 104.34,27.3
X$5032 362 20 363 644 645 cell_1rw
* cell instance $5033 m0 *1 105.045,27.3
X$5033 364 20 365 644 645 cell_1rw
* cell instance $5034 m0 *1 105.75,27.3
X$5034 366 20 367 644 645 cell_1rw
* cell instance $5035 m0 *1 106.455,27.3
X$5035 368 20 369 644 645 cell_1rw
* cell instance $5036 m0 *1 107.16,27.3
X$5036 370 20 371 644 645 cell_1rw
* cell instance $5037 m0 *1 107.865,27.3
X$5037 372 20 373 644 645 cell_1rw
* cell instance $5038 m0 *1 108.57,27.3
X$5038 374 20 375 644 645 cell_1rw
* cell instance $5039 m0 *1 109.275,27.3
X$5039 376 20 377 644 645 cell_1rw
* cell instance $5040 m0 *1 109.98,27.3
X$5040 378 20 379 644 645 cell_1rw
* cell instance $5041 m0 *1 110.685,27.3
X$5041 380 20 381 644 645 cell_1rw
* cell instance $5042 m0 *1 111.39,27.3
X$5042 382 20 383 644 645 cell_1rw
* cell instance $5043 m0 *1 112.095,27.3
X$5043 384 20 385 644 645 cell_1rw
* cell instance $5044 m0 *1 112.8,27.3
X$5044 386 20 387 644 645 cell_1rw
* cell instance $5045 m0 *1 113.505,27.3
X$5045 388 20 389 644 645 cell_1rw
* cell instance $5046 m0 *1 114.21,27.3
X$5046 390 20 391 644 645 cell_1rw
* cell instance $5047 m0 *1 114.915,27.3
X$5047 392 20 393 644 645 cell_1rw
* cell instance $5048 m0 *1 115.62,27.3
X$5048 394 20 395 644 645 cell_1rw
* cell instance $5049 m0 *1 116.325,27.3
X$5049 396 20 397 644 645 cell_1rw
* cell instance $5050 m0 *1 117.03,27.3
X$5050 398 20 399 644 645 cell_1rw
* cell instance $5051 m0 *1 117.735,27.3
X$5051 400 20 401 644 645 cell_1rw
* cell instance $5052 m0 *1 118.44,27.3
X$5052 402 20 403 644 645 cell_1rw
* cell instance $5053 m0 *1 119.145,27.3
X$5053 404 20 405 644 645 cell_1rw
* cell instance $5054 m0 *1 119.85,27.3
X$5054 406 20 407 644 645 cell_1rw
* cell instance $5055 m0 *1 120.555,27.3
X$5055 408 20 409 644 645 cell_1rw
* cell instance $5056 m0 *1 121.26,27.3
X$5056 410 20 411 644 645 cell_1rw
* cell instance $5057 m0 *1 121.965,27.3
X$5057 412 20 413 644 645 cell_1rw
* cell instance $5058 m0 *1 122.67,27.3
X$5058 414 20 415 644 645 cell_1rw
* cell instance $5059 m0 *1 123.375,27.3
X$5059 416 20 417 644 645 cell_1rw
* cell instance $5060 m0 *1 124.08,27.3
X$5060 418 20 419 644 645 cell_1rw
* cell instance $5061 m0 *1 124.785,27.3
X$5061 420 20 421 644 645 cell_1rw
* cell instance $5062 m0 *1 125.49,27.3
X$5062 422 20 423 644 645 cell_1rw
* cell instance $5063 m0 *1 126.195,27.3
X$5063 424 20 425 644 645 cell_1rw
* cell instance $5064 m0 *1 126.9,27.3
X$5064 426 20 427 644 645 cell_1rw
* cell instance $5065 m0 *1 127.605,27.3
X$5065 428 20 429 644 645 cell_1rw
* cell instance $5066 m0 *1 128.31,27.3
X$5066 430 20 431 644 645 cell_1rw
* cell instance $5067 m0 *1 129.015,27.3
X$5067 432 20 433 644 645 cell_1rw
* cell instance $5068 m0 *1 129.72,27.3
X$5068 434 20 435 644 645 cell_1rw
* cell instance $5069 m0 *1 130.425,27.3
X$5069 436 20 437 644 645 cell_1rw
* cell instance $5070 m0 *1 131.13,27.3
X$5070 438 20 439 644 645 cell_1rw
* cell instance $5071 m0 *1 131.835,27.3
X$5071 440 20 441 644 645 cell_1rw
* cell instance $5072 m0 *1 132.54,27.3
X$5072 442 20 443 644 645 cell_1rw
* cell instance $5073 m0 *1 133.245,27.3
X$5073 444 20 445 644 645 cell_1rw
* cell instance $5074 m0 *1 133.95,27.3
X$5074 446 20 447 644 645 cell_1rw
* cell instance $5075 m0 *1 134.655,27.3
X$5075 448 20 449 644 645 cell_1rw
* cell instance $5076 m0 *1 135.36,27.3
X$5076 450 20 451 644 645 cell_1rw
* cell instance $5077 m0 *1 136.065,27.3
X$5077 452 20 453 644 645 cell_1rw
* cell instance $5078 m0 *1 136.77,27.3
X$5078 454 20 455 644 645 cell_1rw
* cell instance $5079 m0 *1 137.475,27.3
X$5079 456 20 457 644 645 cell_1rw
* cell instance $5080 m0 *1 138.18,27.3
X$5080 458 20 459 644 645 cell_1rw
* cell instance $5081 m0 *1 138.885,27.3
X$5081 460 20 461 644 645 cell_1rw
* cell instance $5082 m0 *1 139.59,27.3
X$5082 462 20 463 644 645 cell_1rw
* cell instance $5083 m0 *1 140.295,27.3
X$5083 464 20 465 644 645 cell_1rw
* cell instance $5084 m0 *1 141,27.3
X$5084 466 20 467 644 645 cell_1rw
* cell instance $5085 m0 *1 141.705,27.3
X$5085 468 20 469 644 645 cell_1rw
* cell instance $5086 m0 *1 142.41,27.3
X$5086 470 20 471 644 645 cell_1rw
* cell instance $5087 m0 *1 143.115,27.3
X$5087 472 20 473 644 645 cell_1rw
* cell instance $5088 m0 *1 143.82,27.3
X$5088 474 20 475 644 645 cell_1rw
* cell instance $5089 m0 *1 144.525,27.3
X$5089 476 20 477 644 645 cell_1rw
* cell instance $5090 m0 *1 145.23,27.3
X$5090 478 20 479 644 645 cell_1rw
* cell instance $5091 m0 *1 145.935,27.3
X$5091 480 20 481 644 645 cell_1rw
* cell instance $5092 m0 *1 146.64,27.3
X$5092 482 20 483 644 645 cell_1rw
* cell instance $5093 m0 *1 147.345,27.3
X$5093 484 20 485 644 645 cell_1rw
* cell instance $5094 m0 *1 148.05,27.3
X$5094 486 20 487 644 645 cell_1rw
* cell instance $5095 m0 *1 148.755,27.3
X$5095 488 20 489 644 645 cell_1rw
* cell instance $5096 m0 *1 149.46,27.3
X$5096 490 20 491 644 645 cell_1rw
* cell instance $5097 m0 *1 150.165,27.3
X$5097 492 20 493 644 645 cell_1rw
* cell instance $5098 m0 *1 150.87,27.3
X$5098 494 20 495 644 645 cell_1rw
* cell instance $5099 m0 *1 151.575,27.3
X$5099 496 20 497 644 645 cell_1rw
* cell instance $5100 m0 *1 152.28,27.3
X$5100 498 20 499 644 645 cell_1rw
* cell instance $5101 m0 *1 152.985,27.3
X$5101 500 20 501 644 645 cell_1rw
* cell instance $5102 m0 *1 153.69,27.3
X$5102 502 20 503 644 645 cell_1rw
* cell instance $5103 m0 *1 154.395,27.3
X$5103 504 20 505 644 645 cell_1rw
* cell instance $5104 m0 *1 155.1,27.3
X$5104 506 20 507 644 645 cell_1rw
* cell instance $5105 m0 *1 155.805,27.3
X$5105 508 20 509 644 645 cell_1rw
* cell instance $5106 m0 *1 156.51,27.3
X$5106 510 20 511 644 645 cell_1rw
* cell instance $5107 m0 *1 157.215,27.3
X$5107 512 20 513 644 645 cell_1rw
* cell instance $5108 m0 *1 157.92,27.3
X$5108 514 20 515 644 645 cell_1rw
* cell instance $5109 m0 *1 158.625,27.3
X$5109 516 20 517 644 645 cell_1rw
* cell instance $5110 m0 *1 159.33,27.3
X$5110 518 20 519 644 645 cell_1rw
* cell instance $5111 m0 *1 160.035,27.3
X$5111 520 20 521 644 645 cell_1rw
* cell instance $5112 m0 *1 160.74,27.3
X$5112 522 20 523 644 645 cell_1rw
* cell instance $5113 m0 *1 161.445,27.3
X$5113 524 20 525 644 645 cell_1rw
* cell instance $5114 m0 *1 162.15,27.3
X$5114 526 20 527 644 645 cell_1rw
* cell instance $5115 m0 *1 162.855,27.3
X$5115 528 20 529 644 645 cell_1rw
* cell instance $5116 m0 *1 163.56,27.3
X$5116 530 20 531 644 645 cell_1rw
* cell instance $5117 m0 *1 164.265,27.3
X$5117 532 20 533 644 645 cell_1rw
* cell instance $5118 m0 *1 164.97,27.3
X$5118 534 20 535 644 645 cell_1rw
* cell instance $5119 m0 *1 165.675,27.3
X$5119 536 20 537 644 645 cell_1rw
* cell instance $5120 m0 *1 166.38,27.3
X$5120 538 20 539 644 645 cell_1rw
* cell instance $5121 m0 *1 167.085,27.3
X$5121 540 20 541 644 645 cell_1rw
* cell instance $5122 m0 *1 167.79,27.3
X$5122 542 20 543 644 645 cell_1rw
* cell instance $5123 m0 *1 168.495,27.3
X$5123 544 20 545 644 645 cell_1rw
* cell instance $5124 m0 *1 169.2,27.3
X$5124 546 20 547 644 645 cell_1rw
* cell instance $5125 m0 *1 169.905,27.3
X$5125 548 20 549 644 645 cell_1rw
* cell instance $5126 m0 *1 170.61,27.3
X$5126 550 20 551 644 645 cell_1rw
* cell instance $5127 m0 *1 171.315,27.3
X$5127 552 20 553 644 645 cell_1rw
* cell instance $5128 m0 *1 172.02,27.3
X$5128 554 20 555 644 645 cell_1rw
* cell instance $5129 m0 *1 172.725,27.3
X$5129 556 20 557 644 645 cell_1rw
* cell instance $5130 m0 *1 173.43,27.3
X$5130 558 20 559 644 645 cell_1rw
* cell instance $5131 m0 *1 174.135,27.3
X$5131 560 20 561 644 645 cell_1rw
* cell instance $5132 m0 *1 174.84,27.3
X$5132 562 20 563 644 645 cell_1rw
* cell instance $5133 m0 *1 175.545,27.3
X$5133 564 20 565 644 645 cell_1rw
* cell instance $5134 m0 *1 176.25,27.3
X$5134 566 20 567 644 645 cell_1rw
* cell instance $5135 m0 *1 176.955,27.3
X$5135 568 20 569 644 645 cell_1rw
* cell instance $5136 m0 *1 177.66,27.3
X$5136 570 20 571 644 645 cell_1rw
* cell instance $5137 m0 *1 178.365,27.3
X$5137 572 20 573 644 645 cell_1rw
* cell instance $5138 m0 *1 179.07,27.3
X$5138 574 20 575 644 645 cell_1rw
* cell instance $5139 m0 *1 179.775,27.3
X$5139 576 20 577 644 645 cell_1rw
* cell instance $5140 m0 *1 180.48,27.3
X$5140 578 20 579 644 645 cell_1rw
* cell instance $5141 r0 *1 0.705,27.3
X$5141 67 21 68 644 645 cell_1rw
* cell instance $5142 r0 *1 0,27.3
X$5142 65 21 66 644 645 cell_1rw
* cell instance $5143 r0 *1 1.41,27.3
X$5143 69 21 70 644 645 cell_1rw
* cell instance $5144 r0 *1 2.115,27.3
X$5144 71 21 72 644 645 cell_1rw
* cell instance $5145 r0 *1 2.82,27.3
X$5145 73 21 74 644 645 cell_1rw
* cell instance $5146 r0 *1 3.525,27.3
X$5146 75 21 76 644 645 cell_1rw
* cell instance $5147 r0 *1 4.23,27.3
X$5147 77 21 78 644 645 cell_1rw
* cell instance $5148 r0 *1 4.935,27.3
X$5148 79 21 80 644 645 cell_1rw
* cell instance $5149 r0 *1 5.64,27.3
X$5149 81 21 82 644 645 cell_1rw
* cell instance $5150 r0 *1 6.345,27.3
X$5150 83 21 84 644 645 cell_1rw
* cell instance $5151 r0 *1 7.05,27.3
X$5151 85 21 86 644 645 cell_1rw
* cell instance $5152 r0 *1 7.755,27.3
X$5152 87 21 88 644 645 cell_1rw
* cell instance $5153 r0 *1 8.46,27.3
X$5153 89 21 90 644 645 cell_1rw
* cell instance $5154 r0 *1 9.165,27.3
X$5154 91 21 92 644 645 cell_1rw
* cell instance $5155 r0 *1 9.87,27.3
X$5155 93 21 94 644 645 cell_1rw
* cell instance $5156 r0 *1 10.575,27.3
X$5156 95 21 96 644 645 cell_1rw
* cell instance $5157 r0 *1 11.28,27.3
X$5157 97 21 98 644 645 cell_1rw
* cell instance $5158 r0 *1 11.985,27.3
X$5158 99 21 100 644 645 cell_1rw
* cell instance $5159 r0 *1 12.69,27.3
X$5159 101 21 102 644 645 cell_1rw
* cell instance $5160 r0 *1 13.395,27.3
X$5160 103 21 104 644 645 cell_1rw
* cell instance $5161 r0 *1 14.1,27.3
X$5161 105 21 106 644 645 cell_1rw
* cell instance $5162 r0 *1 14.805,27.3
X$5162 107 21 108 644 645 cell_1rw
* cell instance $5163 r0 *1 15.51,27.3
X$5163 109 21 110 644 645 cell_1rw
* cell instance $5164 r0 *1 16.215,27.3
X$5164 111 21 112 644 645 cell_1rw
* cell instance $5165 r0 *1 16.92,27.3
X$5165 113 21 114 644 645 cell_1rw
* cell instance $5166 r0 *1 17.625,27.3
X$5166 115 21 116 644 645 cell_1rw
* cell instance $5167 r0 *1 18.33,27.3
X$5167 117 21 118 644 645 cell_1rw
* cell instance $5168 r0 *1 19.035,27.3
X$5168 119 21 120 644 645 cell_1rw
* cell instance $5169 r0 *1 19.74,27.3
X$5169 121 21 122 644 645 cell_1rw
* cell instance $5170 r0 *1 20.445,27.3
X$5170 123 21 124 644 645 cell_1rw
* cell instance $5171 r0 *1 21.15,27.3
X$5171 125 21 126 644 645 cell_1rw
* cell instance $5172 r0 *1 21.855,27.3
X$5172 127 21 128 644 645 cell_1rw
* cell instance $5173 r0 *1 22.56,27.3
X$5173 129 21 130 644 645 cell_1rw
* cell instance $5174 r0 *1 23.265,27.3
X$5174 131 21 132 644 645 cell_1rw
* cell instance $5175 r0 *1 23.97,27.3
X$5175 133 21 134 644 645 cell_1rw
* cell instance $5176 r0 *1 24.675,27.3
X$5176 135 21 136 644 645 cell_1rw
* cell instance $5177 r0 *1 25.38,27.3
X$5177 137 21 138 644 645 cell_1rw
* cell instance $5178 r0 *1 26.085,27.3
X$5178 139 21 140 644 645 cell_1rw
* cell instance $5179 r0 *1 26.79,27.3
X$5179 141 21 142 644 645 cell_1rw
* cell instance $5180 r0 *1 27.495,27.3
X$5180 143 21 144 644 645 cell_1rw
* cell instance $5181 r0 *1 28.2,27.3
X$5181 145 21 146 644 645 cell_1rw
* cell instance $5182 r0 *1 28.905,27.3
X$5182 147 21 148 644 645 cell_1rw
* cell instance $5183 r0 *1 29.61,27.3
X$5183 149 21 150 644 645 cell_1rw
* cell instance $5184 r0 *1 30.315,27.3
X$5184 151 21 152 644 645 cell_1rw
* cell instance $5185 r0 *1 31.02,27.3
X$5185 153 21 154 644 645 cell_1rw
* cell instance $5186 r0 *1 31.725,27.3
X$5186 155 21 156 644 645 cell_1rw
* cell instance $5187 r0 *1 32.43,27.3
X$5187 157 21 158 644 645 cell_1rw
* cell instance $5188 r0 *1 33.135,27.3
X$5188 159 21 160 644 645 cell_1rw
* cell instance $5189 r0 *1 33.84,27.3
X$5189 161 21 162 644 645 cell_1rw
* cell instance $5190 r0 *1 34.545,27.3
X$5190 163 21 164 644 645 cell_1rw
* cell instance $5191 r0 *1 35.25,27.3
X$5191 165 21 166 644 645 cell_1rw
* cell instance $5192 r0 *1 35.955,27.3
X$5192 167 21 168 644 645 cell_1rw
* cell instance $5193 r0 *1 36.66,27.3
X$5193 169 21 170 644 645 cell_1rw
* cell instance $5194 r0 *1 37.365,27.3
X$5194 171 21 172 644 645 cell_1rw
* cell instance $5195 r0 *1 38.07,27.3
X$5195 173 21 174 644 645 cell_1rw
* cell instance $5196 r0 *1 38.775,27.3
X$5196 175 21 176 644 645 cell_1rw
* cell instance $5197 r0 *1 39.48,27.3
X$5197 177 21 178 644 645 cell_1rw
* cell instance $5198 r0 *1 40.185,27.3
X$5198 179 21 180 644 645 cell_1rw
* cell instance $5199 r0 *1 40.89,27.3
X$5199 181 21 182 644 645 cell_1rw
* cell instance $5200 r0 *1 41.595,27.3
X$5200 183 21 184 644 645 cell_1rw
* cell instance $5201 r0 *1 42.3,27.3
X$5201 185 21 186 644 645 cell_1rw
* cell instance $5202 r0 *1 43.005,27.3
X$5202 187 21 188 644 645 cell_1rw
* cell instance $5203 r0 *1 43.71,27.3
X$5203 189 21 190 644 645 cell_1rw
* cell instance $5204 r0 *1 44.415,27.3
X$5204 191 21 192 644 645 cell_1rw
* cell instance $5205 r0 *1 45.12,27.3
X$5205 193 21 194 644 645 cell_1rw
* cell instance $5206 r0 *1 45.825,27.3
X$5206 195 21 196 644 645 cell_1rw
* cell instance $5207 r0 *1 46.53,27.3
X$5207 197 21 198 644 645 cell_1rw
* cell instance $5208 r0 *1 47.235,27.3
X$5208 199 21 200 644 645 cell_1rw
* cell instance $5209 r0 *1 47.94,27.3
X$5209 201 21 202 644 645 cell_1rw
* cell instance $5210 r0 *1 48.645,27.3
X$5210 203 21 204 644 645 cell_1rw
* cell instance $5211 r0 *1 49.35,27.3
X$5211 205 21 206 644 645 cell_1rw
* cell instance $5212 r0 *1 50.055,27.3
X$5212 207 21 208 644 645 cell_1rw
* cell instance $5213 r0 *1 50.76,27.3
X$5213 209 21 210 644 645 cell_1rw
* cell instance $5214 r0 *1 51.465,27.3
X$5214 211 21 212 644 645 cell_1rw
* cell instance $5215 r0 *1 52.17,27.3
X$5215 213 21 214 644 645 cell_1rw
* cell instance $5216 r0 *1 52.875,27.3
X$5216 215 21 216 644 645 cell_1rw
* cell instance $5217 r0 *1 53.58,27.3
X$5217 217 21 218 644 645 cell_1rw
* cell instance $5218 r0 *1 54.285,27.3
X$5218 219 21 220 644 645 cell_1rw
* cell instance $5219 r0 *1 54.99,27.3
X$5219 221 21 222 644 645 cell_1rw
* cell instance $5220 r0 *1 55.695,27.3
X$5220 223 21 224 644 645 cell_1rw
* cell instance $5221 r0 *1 56.4,27.3
X$5221 225 21 226 644 645 cell_1rw
* cell instance $5222 r0 *1 57.105,27.3
X$5222 227 21 228 644 645 cell_1rw
* cell instance $5223 r0 *1 57.81,27.3
X$5223 229 21 230 644 645 cell_1rw
* cell instance $5224 r0 *1 58.515,27.3
X$5224 231 21 232 644 645 cell_1rw
* cell instance $5225 r0 *1 59.22,27.3
X$5225 233 21 234 644 645 cell_1rw
* cell instance $5226 r0 *1 59.925,27.3
X$5226 235 21 236 644 645 cell_1rw
* cell instance $5227 r0 *1 60.63,27.3
X$5227 237 21 238 644 645 cell_1rw
* cell instance $5228 r0 *1 61.335,27.3
X$5228 239 21 240 644 645 cell_1rw
* cell instance $5229 r0 *1 62.04,27.3
X$5229 241 21 242 644 645 cell_1rw
* cell instance $5230 r0 *1 62.745,27.3
X$5230 243 21 244 644 645 cell_1rw
* cell instance $5231 r0 *1 63.45,27.3
X$5231 245 21 246 644 645 cell_1rw
* cell instance $5232 r0 *1 64.155,27.3
X$5232 247 21 248 644 645 cell_1rw
* cell instance $5233 r0 *1 64.86,27.3
X$5233 249 21 250 644 645 cell_1rw
* cell instance $5234 r0 *1 65.565,27.3
X$5234 251 21 252 644 645 cell_1rw
* cell instance $5235 r0 *1 66.27,27.3
X$5235 253 21 254 644 645 cell_1rw
* cell instance $5236 r0 *1 66.975,27.3
X$5236 255 21 256 644 645 cell_1rw
* cell instance $5237 r0 *1 67.68,27.3
X$5237 257 21 258 644 645 cell_1rw
* cell instance $5238 r0 *1 68.385,27.3
X$5238 259 21 260 644 645 cell_1rw
* cell instance $5239 r0 *1 69.09,27.3
X$5239 261 21 262 644 645 cell_1rw
* cell instance $5240 r0 *1 69.795,27.3
X$5240 263 21 264 644 645 cell_1rw
* cell instance $5241 r0 *1 70.5,27.3
X$5241 265 21 266 644 645 cell_1rw
* cell instance $5242 r0 *1 71.205,27.3
X$5242 267 21 268 644 645 cell_1rw
* cell instance $5243 r0 *1 71.91,27.3
X$5243 269 21 270 644 645 cell_1rw
* cell instance $5244 r0 *1 72.615,27.3
X$5244 271 21 272 644 645 cell_1rw
* cell instance $5245 r0 *1 73.32,27.3
X$5245 273 21 274 644 645 cell_1rw
* cell instance $5246 r0 *1 74.025,27.3
X$5246 275 21 276 644 645 cell_1rw
* cell instance $5247 r0 *1 74.73,27.3
X$5247 277 21 278 644 645 cell_1rw
* cell instance $5248 r0 *1 75.435,27.3
X$5248 279 21 280 644 645 cell_1rw
* cell instance $5249 r0 *1 76.14,27.3
X$5249 281 21 282 644 645 cell_1rw
* cell instance $5250 r0 *1 76.845,27.3
X$5250 283 21 284 644 645 cell_1rw
* cell instance $5251 r0 *1 77.55,27.3
X$5251 285 21 286 644 645 cell_1rw
* cell instance $5252 r0 *1 78.255,27.3
X$5252 287 21 288 644 645 cell_1rw
* cell instance $5253 r0 *1 78.96,27.3
X$5253 289 21 290 644 645 cell_1rw
* cell instance $5254 r0 *1 79.665,27.3
X$5254 291 21 292 644 645 cell_1rw
* cell instance $5255 r0 *1 80.37,27.3
X$5255 293 21 294 644 645 cell_1rw
* cell instance $5256 r0 *1 81.075,27.3
X$5256 295 21 296 644 645 cell_1rw
* cell instance $5257 r0 *1 81.78,27.3
X$5257 297 21 298 644 645 cell_1rw
* cell instance $5258 r0 *1 82.485,27.3
X$5258 299 21 300 644 645 cell_1rw
* cell instance $5259 r0 *1 83.19,27.3
X$5259 301 21 302 644 645 cell_1rw
* cell instance $5260 r0 *1 83.895,27.3
X$5260 303 21 304 644 645 cell_1rw
* cell instance $5261 r0 *1 84.6,27.3
X$5261 305 21 306 644 645 cell_1rw
* cell instance $5262 r0 *1 85.305,27.3
X$5262 307 21 308 644 645 cell_1rw
* cell instance $5263 r0 *1 86.01,27.3
X$5263 309 21 310 644 645 cell_1rw
* cell instance $5264 r0 *1 86.715,27.3
X$5264 311 21 312 644 645 cell_1rw
* cell instance $5265 r0 *1 87.42,27.3
X$5265 313 21 314 644 645 cell_1rw
* cell instance $5266 r0 *1 88.125,27.3
X$5266 315 21 316 644 645 cell_1rw
* cell instance $5267 r0 *1 88.83,27.3
X$5267 317 21 318 644 645 cell_1rw
* cell instance $5268 r0 *1 89.535,27.3
X$5268 319 21 320 644 645 cell_1rw
* cell instance $5269 r0 *1 90.24,27.3
X$5269 321 21 323 644 645 cell_1rw
* cell instance $5270 r0 *1 90.945,27.3
X$5270 324 21 325 644 645 cell_1rw
* cell instance $5271 r0 *1 91.65,27.3
X$5271 326 21 327 644 645 cell_1rw
* cell instance $5272 r0 *1 92.355,27.3
X$5272 328 21 329 644 645 cell_1rw
* cell instance $5273 r0 *1 93.06,27.3
X$5273 330 21 331 644 645 cell_1rw
* cell instance $5274 r0 *1 93.765,27.3
X$5274 332 21 333 644 645 cell_1rw
* cell instance $5275 r0 *1 94.47,27.3
X$5275 334 21 335 644 645 cell_1rw
* cell instance $5276 r0 *1 95.175,27.3
X$5276 336 21 337 644 645 cell_1rw
* cell instance $5277 r0 *1 95.88,27.3
X$5277 338 21 339 644 645 cell_1rw
* cell instance $5278 r0 *1 96.585,27.3
X$5278 340 21 341 644 645 cell_1rw
* cell instance $5279 r0 *1 97.29,27.3
X$5279 342 21 343 644 645 cell_1rw
* cell instance $5280 r0 *1 97.995,27.3
X$5280 344 21 345 644 645 cell_1rw
* cell instance $5281 r0 *1 98.7,27.3
X$5281 346 21 347 644 645 cell_1rw
* cell instance $5282 r0 *1 99.405,27.3
X$5282 348 21 349 644 645 cell_1rw
* cell instance $5283 r0 *1 100.11,27.3
X$5283 350 21 351 644 645 cell_1rw
* cell instance $5284 r0 *1 100.815,27.3
X$5284 352 21 353 644 645 cell_1rw
* cell instance $5285 r0 *1 101.52,27.3
X$5285 354 21 355 644 645 cell_1rw
* cell instance $5286 r0 *1 102.225,27.3
X$5286 356 21 357 644 645 cell_1rw
* cell instance $5287 r0 *1 102.93,27.3
X$5287 358 21 359 644 645 cell_1rw
* cell instance $5288 r0 *1 103.635,27.3
X$5288 360 21 361 644 645 cell_1rw
* cell instance $5289 r0 *1 104.34,27.3
X$5289 362 21 363 644 645 cell_1rw
* cell instance $5290 r0 *1 105.045,27.3
X$5290 364 21 365 644 645 cell_1rw
* cell instance $5291 r0 *1 105.75,27.3
X$5291 366 21 367 644 645 cell_1rw
* cell instance $5292 r0 *1 106.455,27.3
X$5292 368 21 369 644 645 cell_1rw
* cell instance $5293 r0 *1 107.16,27.3
X$5293 370 21 371 644 645 cell_1rw
* cell instance $5294 r0 *1 107.865,27.3
X$5294 372 21 373 644 645 cell_1rw
* cell instance $5295 r0 *1 108.57,27.3
X$5295 374 21 375 644 645 cell_1rw
* cell instance $5296 r0 *1 109.275,27.3
X$5296 376 21 377 644 645 cell_1rw
* cell instance $5297 r0 *1 109.98,27.3
X$5297 378 21 379 644 645 cell_1rw
* cell instance $5298 r0 *1 110.685,27.3
X$5298 380 21 381 644 645 cell_1rw
* cell instance $5299 r0 *1 111.39,27.3
X$5299 382 21 383 644 645 cell_1rw
* cell instance $5300 r0 *1 112.095,27.3
X$5300 384 21 385 644 645 cell_1rw
* cell instance $5301 r0 *1 112.8,27.3
X$5301 386 21 387 644 645 cell_1rw
* cell instance $5302 r0 *1 113.505,27.3
X$5302 388 21 389 644 645 cell_1rw
* cell instance $5303 r0 *1 114.21,27.3
X$5303 390 21 391 644 645 cell_1rw
* cell instance $5304 r0 *1 114.915,27.3
X$5304 392 21 393 644 645 cell_1rw
* cell instance $5305 r0 *1 115.62,27.3
X$5305 394 21 395 644 645 cell_1rw
* cell instance $5306 r0 *1 116.325,27.3
X$5306 396 21 397 644 645 cell_1rw
* cell instance $5307 r0 *1 117.03,27.3
X$5307 398 21 399 644 645 cell_1rw
* cell instance $5308 r0 *1 117.735,27.3
X$5308 400 21 401 644 645 cell_1rw
* cell instance $5309 r0 *1 118.44,27.3
X$5309 402 21 403 644 645 cell_1rw
* cell instance $5310 r0 *1 119.145,27.3
X$5310 404 21 405 644 645 cell_1rw
* cell instance $5311 r0 *1 119.85,27.3
X$5311 406 21 407 644 645 cell_1rw
* cell instance $5312 r0 *1 120.555,27.3
X$5312 408 21 409 644 645 cell_1rw
* cell instance $5313 r0 *1 121.26,27.3
X$5313 410 21 411 644 645 cell_1rw
* cell instance $5314 r0 *1 121.965,27.3
X$5314 412 21 413 644 645 cell_1rw
* cell instance $5315 r0 *1 122.67,27.3
X$5315 414 21 415 644 645 cell_1rw
* cell instance $5316 r0 *1 123.375,27.3
X$5316 416 21 417 644 645 cell_1rw
* cell instance $5317 r0 *1 124.08,27.3
X$5317 418 21 419 644 645 cell_1rw
* cell instance $5318 r0 *1 124.785,27.3
X$5318 420 21 421 644 645 cell_1rw
* cell instance $5319 r0 *1 125.49,27.3
X$5319 422 21 423 644 645 cell_1rw
* cell instance $5320 r0 *1 126.195,27.3
X$5320 424 21 425 644 645 cell_1rw
* cell instance $5321 r0 *1 126.9,27.3
X$5321 426 21 427 644 645 cell_1rw
* cell instance $5322 r0 *1 127.605,27.3
X$5322 428 21 429 644 645 cell_1rw
* cell instance $5323 r0 *1 128.31,27.3
X$5323 430 21 431 644 645 cell_1rw
* cell instance $5324 r0 *1 129.015,27.3
X$5324 432 21 433 644 645 cell_1rw
* cell instance $5325 r0 *1 129.72,27.3
X$5325 434 21 435 644 645 cell_1rw
* cell instance $5326 r0 *1 130.425,27.3
X$5326 436 21 437 644 645 cell_1rw
* cell instance $5327 r0 *1 131.13,27.3
X$5327 438 21 439 644 645 cell_1rw
* cell instance $5328 r0 *1 131.835,27.3
X$5328 440 21 441 644 645 cell_1rw
* cell instance $5329 r0 *1 132.54,27.3
X$5329 442 21 443 644 645 cell_1rw
* cell instance $5330 r0 *1 133.245,27.3
X$5330 444 21 445 644 645 cell_1rw
* cell instance $5331 r0 *1 133.95,27.3
X$5331 446 21 447 644 645 cell_1rw
* cell instance $5332 r0 *1 134.655,27.3
X$5332 448 21 449 644 645 cell_1rw
* cell instance $5333 r0 *1 135.36,27.3
X$5333 450 21 451 644 645 cell_1rw
* cell instance $5334 r0 *1 136.065,27.3
X$5334 452 21 453 644 645 cell_1rw
* cell instance $5335 r0 *1 136.77,27.3
X$5335 454 21 455 644 645 cell_1rw
* cell instance $5336 r0 *1 137.475,27.3
X$5336 456 21 457 644 645 cell_1rw
* cell instance $5337 r0 *1 138.18,27.3
X$5337 458 21 459 644 645 cell_1rw
* cell instance $5338 r0 *1 138.885,27.3
X$5338 460 21 461 644 645 cell_1rw
* cell instance $5339 r0 *1 139.59,27.3
X$5339 462 21 463 644 645 cell_1rw
* cell instance $5340 r0 *1 140.295,27.3
X$5340 464 21 465 644 645 cell_1rw
* cell instance $5341 r0 *1 141,27.3
X$5341 466 21 467 644 645 cell_1rw
* cell instance $5342 r0 *1 141.705,27.3
X$5342 468 21 469 644 645 cell_1rw
* cell instance $5343 r0 *1 142.41,27.3
X$5343 470 21 471 644 645 cell_1rw
* cell instance $5344 r0 *1 143.115,27.3
X$5344 472 21 473 644 645 cell_1rw
* cell instance $5345 r0 *1 143.82,27.3
X$5345 474 21 475 644 645 cell_1rw
* cell instance $5346 r0 *1 144.525,27.3
X$5346 476 21 477 644 645 cell_1rw
* cell instance $5347 r0 *1 145.23,27.3
X$5347 478 21 479 644 645 cell_1rw
* cell instance $5348 r0 *1 145.935,27.3
X$5348 480 21 481 644 645 cell_1rw
* cell instance $5349 r0 *1 146.64,27.3
X$5349 482 21 483 644 645 cell_1rw
* cell instance $5350 r0 *1 147.345,27.3
X$5350 484 21 485 644 645 cell_1rw
* cell instance $5351 r0 *1 148.05,27.3
X$5351 486 21 487 644 645 cell_1rw
* cell instance $5352 r0 *1 148.755,27.3
X$5352 488 21 489 644 645 cell_1rw
* cell instance $5353 r0 *1 149.46,27.3
X$5353 490 21 491 644 645 cell_1rw
* cell instance $5354 r0 *1 150.165,27.3
X$5354 492 21 493 644 645 cell_1rw
* cell instance $5355 r0 *1 150.87,27.3
X$5355 494 21 495 644 645 cell_1rw
* cell instance $5356 r0 *1 151.575,27.3
X$5356 496 21 497 644 645 cell_1rw
* cell instance $5357 r0 *1 152.28,27.3
X$5357 498 21 499 644 645 cell_1rw
* cell instance $5358 r0 *1 152.985,27.3
X$5358 500 21 501 644 645 cell_1rw
* cell instance $5359 r0 *1 153.69,27.3
X$5359 502 21 503 644 645 cell_1rw
* cell instance $5360 r0 *1 154.395,27.3
X$5360 504 21 505 644 645 cell_1rw
* cell instance $5361 r0 *1 155.1,27.3
X$5361 506 21 507 644 645 cell_1rw
* cell instance $5362 r0 *1 155.805,27.3
X$5362 508 21 509 644 645 cell_1rw
* cell instance $5363 r0 *1 156.51,27.3
X$5363 510 21 511 644 645 cell_1rw
* cell instance $5364 r0 *1 157.215,27.3
X$5364 512 21 513 644 645 cell_1rw
* cell instance $5365 r0 *1 157.92,27.3
X$5365 514 21 515 644 645 cell_1rw
* cell instance $5366 r0 *1 158.625,27.3
X$5366 516 21 517 644 645 cell_1rw
* cell instance $5367 r0 *1 159.33,27.3
X$5367 518 21 519 644 645 cell_1rw
* cell instance $5368 r0 *1 160.035,27.3
X$5368 520 21 521 644 645 cell_1rw
* cell instance $5369 r0 *1 160.74,27.3
X$5369 522 21 523 644 645 cell_1rw
* cell instance $5370 r0 *1 161.445,27.3
X$5370 524 21 525 644 645 cell_1rw
* cell instance $5371 r0 *1 162.15,27.3
X$5371 526 21 527 644 645 cell_1rw
* cell instance $5372 r0 *1 162.855,27.3
X$5372 528 21 529 644 645 cell_1rw
* cell instance $5373 r0 *1 163.56,27.3
X$5373 530 21 531 644 645 cell_1rw
* cell instance $5374 r0 *1 164.265,27.3
X$5374 532 21 533 644 645 cell_1rw
* cell instance $5375 r0 *1 164.97,27.3
X$5375 534 21 535 644 645 cell_1rw
* cell instance $5376 r0 *1 165.675,27.3
X$5376 536 21 537 644 645 cell_1rw
* cell instance $5377 r0 *1 166.38,27.3
X$5377 538 21 539 644 645 cell_1rw
* cell instance $5378 r0 *1 167.085,27.3
X$5378 540 21 541 644 645 cell_1rw
* cell instance $5379 r0 *1 167.79,27.3
X$5379 542 21 543 644 645 cell_1rw
* cell instance $5380 r0 *1 168.495,27.3
X$5380 544 21 545 644 645 cell_1rw
* cell instance $5381 r0 *1 169.2,27.3
X$5381 546 21 547 644 645 cell_1rw
* cell instance $5382 r0 *1 169.905,27.3
X$5382 548 21 549 644 645 cell_1rw
* cell instance $5383 r0 *1 170.61,27.3
X$5383 550 21 551 644 645 cell_1rw
* cell instance $5384 r0 *1 171.315,27.3
X$5384 552 21 553 644 645 cell_1rw
* cell instance $5385 r0 *1 172.02,27.3
X$5385 554 21 555 644 645 cell_1rw
* cell instance $5386 r0 *1 172.725,27.3
X$5386 556 21 557 644 645 cell_1rw
* cell instance $5387 r0 *1 173.43,27.3
X$5387 558 21 559 644 645 cell_1rw
* cell instance $5388 r0 *1 174.135,27.3
X$5388 560 21 561 644 645 cell_1rw
* cell instance $5389 r0 *1 174.84,27.3
X$5389 562 21 563 644 645 cell_1rw
* cell instance $5390 r0 *1 175.545,27.3
X$5390 564 21 565 644 645 cell_1rw
* cell instance $5391 r0 *1 176.25,27.3
X$5391 566 21 567 644 645 cell_1rw
* cell instance $5392 r0 *1 176.955,27.3
X$5392 568 21 569 644 645 cell_1rw
* cell instance $5393 r0 *1 177.66,27.3
X$5393 570 21 571 644 645 cell_1rw
* cell instance $5394 r0 *1 178.365,27.3
X$5394 572 21 573 644 645 cell_1rw
* cell instance $5395 r0 *1 179.07,27.3
X$5395 574 21 575 644 645 cell_1rw
* cell instance $5396 r0 *1 179.775,27.3
X$5396 576 21 577 644 645 cell_1rw
* cell instance $5397 r0 *1 180.48,27.3
X$5397 578 21 579 644 645 cell_1rw
* cell instance $5398 m0 *1 0.705,30.03
X$5398 67 22 68 644 645 cell_1rw
* cell instance $5399 m0 *1 0,30.03
X$5399 65 22 66 644 645 cell_1rw
* cell instance $5400 m0 *1 1.41,30.03
X$5400 69 22 70 644 645 cell_1rw
* cell instance $5401 m0 *1 2.115,30.03
X$5401 71 22 72 644 645 cell_1rw
* cell instance $5402 m0 *1 2.82,30.03
X$5402 73 22 74 644 645 cell_1rw
* cell instance $5403 m0 *1 3.525,30.03
X$5403 75 22 76 644 645 cell_1rw
* cell instance $5404 m0 *1 4.23,30.03
X$5404 77 22 78 644 645 cell_1rw
* cell instance $5405 m0 *1 4.935,30.03
X$5405 79 22 80 644 645 cell_1rw
* cell instance $5406 m0 *1 5.64,30.03
X$5406 81 22 82 644 645 cell_1rw
* cell instance $5407 m0 *1 6.345,30.03
X$5407 83 22 84 644 645 cell_1rw
* cell instance $5408 m0 *1 7.05,30.03
X$5408 85 22 86 644 645 cell_1rw
* cell instance $5409 m0 *1 7.755,30.03
X$5409 87 22 88 644 645 cell_1rw
* cell instance $5410 m0 *1 8.46,30.03
X$5410 89 22 90 644 645 cell_1rw
* cell instance $5411 m0 *1 9.165,30.03
X$5411 91 22 92 644 645 cell_1rw
* cell instance $5412 m0 *1 9.87,30.03
X$5412 93 22 94 644 645 cell_1rw
* cell instance $5413 m0 *1 10.575,30.03
X$5413 95 22 96 644 645 cell_1rw
* cell instance $5414 m0 *1 11.28,30.03
X$5414 97 22 98 644 645 cell_1rw
* cell instance $5415 m0 *1 11.985,30.03
X$5415 99 22 100 644 645 cell_1rw
* cell instance $5416 m0 *1 12.69,30.03
X$5416 101 22 102 644 645 cell_1rw
* cell instance $5417 m0 *1 13.395,30.03
X$5417 103 22 104 644 645 cell_1rw
* cell instance $5418 m0 *1 14.1,30.03
X$5418 105 22 106 644 645 cell_1rw
* cell instance $5419 m0 *1 14.805,30.03
X$5419 107 22 108 644 645 cell_1rw
* cell instance $5420 m0 *1 15.51,30.03
X$5420 109 22 110 644 645 cell_1rw
* cell instance $5421 m0 *1 16.215,30.03
X$5421 111 22 112 644 645 cell_1rw
* cell instance $5422 m0 *1 16.92,30.03
X$5422 113 22 114 644 645 cell_1rw
* cell instance $5423 m0 *1 17.625,30.03
X$5423 115 22 116 644 645 cell_1rw
* cell instance $5424 m0 *1 18.33,30.03
X$5424 117 22 118 644 645 cell_1rw
* cell instance $5425 m0 *1 19.035,30.03
X$5425 119 22 120 644 645 cell_1rw
* cell instance $5426 m0 *1 19.74,30.03
X$5426 121 22 122 644 645 cell_1rw
* cell instance $5427 m0 *1 20.445,30.03
X$5427 123 22 124 644 645 cell_1rw
* cell instance $5428 m0 *1 21.15,30.03
X$5428 125 22 126 644 645 cell_1rw
* cell instance $5429 m0 *1 21.855,30.03
X$5429 127 22 128 644 645 cell_1rw
* cell instance $5430 m0 *1 22.56,30.03
X$5430 129 22 130 644 645 cell_1rw
* cell instance $5431 m0 *1 23.265,30.03
X$5431 131 22 132 644 645 cell_1rw
* cell instance $5432 m0 *1 23.97,30.03
X$5432 133 22 134 644 645 cell_1rw
* cell instance $5433 m0 *1 24.675,30.03
X$5433 135 22 136 644 645 cell_1rw
* cell instance $5434 m0 *1 25.38,30.03
X$5434 137 22 138 644 645 cell_1rw
* cell instance $5435 m0 *1 26.085,30.03
X$5435 139 22 140 644 645 cell_1rw
* cell instance $5436 m0 *1 26.79,30.03
X$5436 141 22 142 644 645 cell_1rw
* cell instance $5437 m0 *1 27.495,30.03
X$5437 143 22 144 644 645 cell_1rw
* cell instance $5438 m0 *1 28.2,30.03
X$5438 145 22 146 644 645 cell_1rw
* cell instance $5439 m0 *1 28.905,30.03
X$5439 147 22 148 644 645 cell_1rw
* cell instance $5440 m0 *1 29.61,30.03
X$5440 149 22 150 644 645 cell_1rw
* cell instance $5441 m0 *1 30.315,30.03
X$5441 151 22 152 644 645 cell_1rw
* cell instance $5442 m0 *1 31.02,30.03
X$5442 153 22 154 644 645 cell_1rw
* cell instance $5443 m0 *1 31.725,30.03
X$5443 155 22 156 644 645 cell_1rw
* cell instance $5444 m0 *1 32.43,30.03
X$5444 157 22 158 644 645 cell_1rw
* cell instance $5445 m0 *1 33.135,30.03
X$5445 159 22 160 644 645 cell_1rw
* cell instance $5446 m0 *1 33.84,30.03
X$5446 161 22 162 644 645 cell_1rw
* cell instance $5447 m0 *1 34.545,30.03
X$5447 163 22 164 644 645 cell_1rw
* cell instance $5448 m0 *1 35.25,30.03
X$5448 165 22 166 644 645 cell_1rw
* cell instance $5449 m0 *1 35.955,30.03
X$5449 167 22 168 644 645 cell_1rw
* cell instance $5450 m0 *1 36.66,30.03
X$5450 169 22 170 644 645 cell_1rw
* cell instance $5451 m0 *1 37.365,30.03
X$5451 171 22 172 644 645 cell_1rw
* cell instance $5452 m0 *1 38.07,30.03
X$5452 173 22 174 644 645 cell_1rw
* cell instance $5453 m0 *1 38.775,30.03
X$5453 175 22 176 644 645 cell_1rw
* cell instance $5454 m0 *1 39.48,30.03
X$5454 177 22 178 644 645 cell_1rw
* cell instance $5455 m0 *1 40.185,30.03
X$5455 179 22 180 644 645 cell_1rw
* cell instance $5456 m0 *1 40.89,30.03
X$5456 181 22 182 644 645 cell_1rw
* cell instance $5457 m0 *1 41.595,30.03
X$5457 183 22 184 644 645 cell_1rw
* cell instance $5458 m0 *1 42.3,30.03
X$5458 185 22 186 644 645 cell_1rw
* cell instance $5459 m0 *1 43.005,30.03
X$5459 187 22 188 644 645 cell_1rw
* cell instance $5460 m0 *1 43.71,30.03
X$5460 189 22 190 644 645 cell_1rw
* cell instance $5461 m0 *1 44.415,30.03
X$5461 191 22 192 644 645 cell_1rw
* cell instance $5462 m0 *1 45.12,30.03
X$5462 193 22 194 644 645 cell_1rw
* cell instance $5463 m0 *1 45.825,30.03
X$5463 195 22 196 644 645 cell_1rw
* cell instance $5464 m0 *1 46.53,30.03
X$5464 197 22 198 644 645 cell_1rw
* cell instance $5465 m0 *1 47.235,30.03
X$5465 199 22 200 644 645 cell_1rw
* cell instance $5466 m0 *1 47.94,30.03
X$5466 201 22 202 644 645 cell_1rw
* cell instance $5467 m0 *1 48.645,30.03
X$5467 203 22 204 644 645 cell_1rw
* cell instance $5468 m0 *1 49.35,30.03
X$5468 205 22 206 644 645 cell_1rw
* cell instance $5469 m0 *1 50.055,30.03
X$5469 207 22 208 644 645 cell_1rw
* cell instance $5470 m0 *1 50.76,30.03
X$5470 209 22 210 644 645 cell_1rw
* cell instance $5471 m0 *1 51.465,30.03
X$5471 211 22 212 644 645 cell_1rw
* cell instance $5472 m0 *1 52.17,30.03
X$5472 213 22 214 644 645 cell_1rw
* cell instance $5473 m0 *1 52.875,30.03
X$5473 215 22 216 644 645 cell_1rw
* cell instance $5474 m0 *1 53.58,30.03
X$5474 217 22 218 644 645 cell_1rw
* cell instance $5475 m0 *1 54.285,30.03
X$5475 219 22 220 644 645 cell_1rw
* cell instance $5476 m0 *1 54.99,30.03
X$5476 221 22 222 644 645 cell_1rw
* cell instance $5477 m0 *1 55.695,30.03
X$5477 223 22 224 644 645 cell_1rw
* cell instance $5478 m0 *1 56.4,30.03
X$5478 225 22 226 644 645 cell_1rw
* cell instance $5479 m0 *1 57.105,30.03
X$5479 227 22 228 644 645 cell_1rw
* cell instance $5480 m0 *1 57.81,30.03
X$5480 229 22 230 644 645 cell_1rw
* cell instance $5481 m0 *1 58.515,30.03
X$5481 231 22 232 644 645 cell_1rw
* cell instance $5482 m0 *1 59.22,30.03
X$5482 233 22 234 644 645 cell_1rw
* cell instance $5483 m0 *1 59.925,30.03
X$5483 235 22 236 644 645 cell_1rw
* cell instance $5484 m0 *1 60.63,30.03
X$5484 237 22 238 644 645 cell_1rw
* cell instance $5485 m0 *1 61.335,30.03
X$5485 239 22 240 644 645 cell_1rw
* cell instance $5486 m0 *1 62.04,30.03
X$5486 241 22 242 644 645 cell_1rw
* cell instance $5487 m0 *1 62.745,30.03
X$5487 243 22 244 644 645 cell_1rw
* cell instance $5488 m0 *1 63.45,30.03
X$5488 245 22 246 644 645 cell_1rw
* cell instance $5489 m0 *1 64.155,30.03
X$5489 247 22 248 644 645 cell_1rw
* cell instance $5490 m0 *1 64.86,30.03
X$5490 249 22 250 644 645 cell_1rw
* cell instance $5491 m0 *1 65.565,30.03
X$5491 251 22 252 644 645 cell_1rw
* cell instance $5492 m0 *1 66.27,30.03
X$5492 253 22 254 644 645 cell_1rw
* cell instance $5493 m0 *1 66.975,30.03
X$5493 255 22 256 644 645 cell_1rw
* cell instance $5494 m0 *1 67.68,30.03
X$5494 257 22 258 644 645 cell_1rw
* cell instance $5495 m0 *1 68.385,30.03
X$5495 259 22 260 644 645 cell_1rw
* cell instance $5496 m0 *1 69.09,30.03
X$5496 261 22 262 644 645 cell_1rw
* cell instance $5497 m0 *1 69.795,30.03
X$5497 263 22 264 644 645 cell_1rw
* cell instance $5498 m0 *1 70.5,30.03
X$5498 265 22 266 644 645 cell_1rw
* cell instance $5499 m0 *1 71.205,30.03
X$5499 267 22 268 644 645 cell_1rw
* cell instance $5500 m0 *1 71.91,30.03
X$5500 269 22 270 644 645 cell_1rw
* cell instance $5501 m0 *1 72.615,30.03
X$5501 271 22 272 644 645 cell_1rw
* cell instance $5502 m0 *1 73.32,30.03
X$5502 273 22 274 644 645 cell_1rw
* cell instance $5503 m0 *1 74.025,30.03
X$5503 275 22 276 644 645 cell_1rw
* cell instance $5504 m0 *1 74.73,30.03
X$5504 277 22 278 644 645 cell_1rw
* cell instance $5505 m0 *1 75.435,30.03
X$5505 279 22 280 644 645 cell_1rw
* cell instance $5506 m0 *1 76.14,30.03
X$5506 281 22 282 644 645 cell_1rw
* cell instance $5507 m0 *1 76.845,30.03
X$5507 283 22 284 644 645 cell_1rw
* cell instance $5508 m0 *1 77.55,30.03
X$5508 285 22 286 644 645 cell_1rw
* cell instance $5509 m0 *1 78.255,30.03
X$5509 287 22 288 644 645 cell_1rw
* cell instance $5510 m0 *1 78.96,30.03
X$5510 289 22 290 644 645 cell_1rw
* cell instance $5511 m0 *1 79.665,30.03
X$5511 291 22 292 644 645 cell_1rw
* cell instance $5512 m0 *1 80.37,30.03
X$5512 293 22 294 644 645 cell_1rw
* cell instance $5513 m0 *1 81.075,30.03
X$5513 295 22 296 644 645 cell_1rw
* cell instance $5514 m0 *1 81.78,30.03
X$5514 297 22 298 644 645 cell_1rw
* cell instance $5515 m0 *1 82.485,30.03
X$5515 299 22 300 644 645 cell_1rw
* cell instance $5516 m0 *1 83.19,30.03
X$5516 301 22 302 644 645 cell_1rw
* cell instance $5517 m0 *1 83.895,30.03
X$5517 303 22 304 644 645 cell_1rw
* cell instance $5518 m0 *1 84.6,30.03
X$5518 305 22 306 644 645 cell_1rw
* cell instance $5519 m0 *1 85.305,30.03
X$5519 307 22 308 644 645 cell_1rw
* cell instance $5520 m0 *1 86.01,30.03
X$5520 309 22 310 644 645 cell_1rw
* cell instance $5521 m0 *1 86.715,30.03
X$5521 311 22 312 644 645 cell_1rw
* cell instance $5522 m0 *1 87.42,30.03
X$5522 313 22 314 644 645 cell_1rw
* cell instance $5523 m0 *1 88.125,30.03
X$5523 315 22 316 644 645 cell_1rw
* cell instance $5524 m0 *1 88.83,30.03
X$5524 317 22 318 644 645 cell_1rw
* cell instance $5525 m0 *1 89.535,30.03
X$5525 319 22 320 644 645 cell_1rw
* cell instance $5526 m0 *1 90.24,30.03
X$5526 321 22 323 644 645 cell_1rw
* cell instance $5527 m0 *1 90.945,30.03
X$5527 324 22 325 644 645 cell_1rw
* cell instance $5528 m0 *1 91.65,30.03
X$5528 326 22 327 644 645 cell_1rw
* cell instance $5529 m0 *1 92.355,30.03
X$5529 328 22 329 644 645 cell_1rw
* cell instance $5530 m0 *1 93.06,30.03
X$5530 330 22 331 644 645 cell_1rw
* cell instance $5531 m0 *1 93.765,30.03
X$5531 332 22 333 644 645 cell_1rw
* cell instance $5532 m0 *1 94.47,30.03
X$5532 334 22 335 644 645 cell_1rw
* cell instance $5533 m0 *1 95.175,30.03
X$5533 336 22 337 644 645 cell_1rw
* cell instance $5534 m0 *1 95.88,30.03
X$5534 338 22 339 644 645 cell_1rw
* cell instance $5535 m0 *1 96.585,30.03
X$5535 340 22 341 644 645 cell_1rw
* cell instance $5536 m0 *1 97.29,30.03
X$5536 342 22 343 644 645 cell_1rw
* cell instance $5537 m0 *1 97.995,30.03
X$5537 344 22 345 644 645 cell_1rw
* cell instance $5538 m0 *1 98.7,30.03
X$5538 346 22 347 644 645 cell_1rw
* cell instance $5539 m0 *1 99.405,30.03
X$5539 348 22 349 644 645 cell_1rw
* cell instance $5540 m0 *1 100.11,30.03
X$5540 350 22 351 644 645 cell_1rw
* cell instance $5541 m0 *1 100.815,30.03
X$5541 352 22 353 644 645 cell_1rw
* cell instance $5542 m0 *1 101.52,30.03
X$5542 354 22 355 644 645 cell_1rw
* cell instance $5543 m0 *1 102.225,30.03
X$5543 356 22 357 644 645 cell_1rw
* cell instance $5544 m0 *1 102.93,30.03
X$5544 358 22 359 644 645 cell_1rw
* cell instance $5545 m0 *1 103.635,30.03
X$5545 360 22 361 644 645 cell_1rw
* cell instance $5546 m0 *1 104.34,30.03
X$5546 362 22 363 644 645 cell_1rw
* cell instance $5547 m0 *1 105.045,30.03
X$5547 364 22 365 644 645 cell_1rw
* cell instance $5548 m0 *1 105.75,30.03
X$5548 366 22 367 644 645 cell_1rw
* cell instance $5549 m0 *1 106.455,30.03
X$5549 368 22 369 644 645 cell_1rw
* cell instance $5550 m0 *1 107.16,30.03
X$5550 370 22 371 644 645 cell_1rw
* cell instance $5551 m0 *1 107.865,30.03
X$5551 372 22 373 644 645 cell_1rw
* cell instance $5552 m0 *1 108.57,30.03
X$5552 374 22 375 644 645 cell_1rw
* cell instance $5553 m0 *1 109.275,30.03
X$5553 376 22 377 644 645 cell_1rw
* cell instance $5554 m0 *1 109.98,30.03
X$5554 378 22 379 644 645 cell_1rw
* cell instance $5555 m0 *1 110.685,30.03
X$5555 380 22 381 644 645 cell_1rw
* cell instance $5556 m0 *1 111.39,30.03
X$5556 382 22 383 644 645 cell_1rw
* cell instance $5557 m0 *1 112.095,30.03
X$5557 384 22 385 644 645 cell_1rw
* cell instance $5558 m0 *1 112.8,30.03
X$5558 386 22 387 644 645 cell_1rw
* cell instance $5559 m0 *1 113.505,30.03
X$5559 388 22 389 644 645 cell_1rw
* cell instance $5560 m0 *1 114.21,30.03
X$5560 390 22 391 644 645 cell_1rw
* cell instance $5561 m0 *1 114.915,30.03
X$5561 392 22 393 644 645 cell_1rw
* cell instance $5562 m0 *1 115.62,30.03
X$5562 394 22 395 644 645 cell_1rw
* cell instance $5563 m0 *1 116.325,30.03
X$5563 396 22 397 644 645 cell_1rw
* cell instance $5564 m0 *1 117.03,30.03
X$5564 398 22 399 644 645 cell_1rw
* cell instance $5565 m0 *1 117.735,30.03
X$5565 400 22 401 644 645 cell_1rw
* cell instance $5566 m0 *1 118.44,30.03
X$5566 402 22 403 644 645 cell_1rw
* cell instance $5567 m0 *1 119.145,30.03
X$5567 404 22 405 644 645 cell_1rw
* cell instance $5568 m0 *1 119.85,30.03
X$5568 406 22 407 644 645 cell_1rw
* cell instance $5569 m0 *1 120.555,30.03
X$5569 408 22 409 644 645 cell_1rw
* cell instance $5570 m0 *1 121.26,30.03
X$5570 410 22 411 644 645 cell_1rw
* cell instance $5571 m0 *1 121.965,30.03
X$5571 412 22 413 644 645 cell_1rw
* cell instance $5572 m0 *1 122.67,30.03
X$5572 414 22 415 644 645 cell_1rw
* cell instance $5573 m0 *1 123.375,30.03
X$5573 416 22 417 644 645 cell_1rw
* cell instance $5574 m0 *1 124.08,30.03
X$5574 418 22 419 644 645 cell_1rw
* cell instance $5575 m0 *1 124.785,30.03
X$5575 420 22 421 644 645 cell_1rw
* cell instance $5576 m0 *1 125.49,30.03
X$5576 422 22 423 644 645 cell_1rw
* cell instance $5577 m0 *1 126.195,30.03
X$5577 424 22 425 644 645 cell_1rw
* cell instance $5578 m0 *1 126.9,30.03
X$5578 426 22 427 644 645 cell_1rw
* cell instance $5579 m0 *1 127.605,30.03
X$5579 428 22 429 644 645 cell_1rw
* cell instance $5580 m0 *1 128.31,30.03
X$5580 430 22 431 644 645 cell_1rw
* cell instance $5581 m0 *1 129.015,30.03
X$5581 432 22 433 644 645 cell_1rw
* cell instance $5582 m0 *1 129.72,30.03
X$5582 434 22 435 644 645 cell_1rw
* cell instance $5583 m0 *1 130.425,30.03
X$5583 436 22 437 644 645 cell_1rw
* cell instance $5584 m0 *1 131.13,30.03
X$5584 438 22 439 644 645 cell_1rw
* cell instance $5585 m0 *1 131.835,30.03
X$5585 440 22 441 644 645 cell_1rw
* cell instance $5586 m0 *1 132.54,30.03
X$5586 442 22 443 644 645 cell_1rw
* cell instance $5587 m0 *1 133.245,30.03
X$5587 444 22 445 644 645 cell_1rw
* cell instance $5588 m0 *1 133.95,30.03
X$5588 446 22 447 644 645 cell_1rw
* cell instance $5589 m0 *1 134.655,30.03
X$5589 448 22 449 644 645 cell_1rw
* cell instance $5590 m0 *1 135.36,30.03
X$5590 450 22 451 644 645 cell_1rw
* cell instance $5591 m0 *1 136.065,30.03
X$5591 452 22 453 644 645 cell_1rw
* cell instance $5592 m0 *1 136.77,30.03
X$5592 454 22 455 644 645 cell_1rw
* cell instance $5593 m0 *1 137.475,30.03
X$5593 456 22 457 644 645 cell_1rw
* cell instance $5594 m0 *1 138.18,30.03
X$5594 458 22 459 644 645 cell_1rw
* cell instance $5595 m0 *1 138.885,30.03
X$5595 460 22 461 644 645 cell_1rw
* cell instance $5596 m0 *1 139.59,30.03
X$5596 462 22 463 644 645 cell_1rw
* cell instance $5597 m0 *1 140.295,30.03
X$5597 464 22 465 644 645 cell_1rw
* cell instance $5598 m0 *1 141,30.03
X$5598 466 22 467 644 645 cell_1rw
* cell instance $5599 m0 *1 141.705,30.03
X$5599 468 22 469 644 645 cell_1rw
* cell instance $5600 m0 *1 142.41,30.03
X$5600 470 22 471 644 645 cell_1rw
* cell instance $5601 m0 *1 143.115,30.03
X$5601 472 22 473 644 645 cell_1rw
* cell instance $5602 m0 *1 143.82,30.03
X$5602 474 22 475 644 645 cell_1rw
* cell instance $5603 m0 *1 144.525,30.03
X$5603 476 22 477 644 645 cell_1rw
* cell instance $5604 m0 *1 145.23,30.03
X$5604 478 22 479 644 645 cell_1rw
* cell instance $5605 m0 *1 145.935,30.03
X$5605 480 22 481 644 645 cell_1rw
* cell instance $5606 m0 *1 146.64,30.03
X$5606 482 22 483 644 645 cell_1rw
* cell instance $5607 m0 *1 147.345,30.03
X$5607 484 22 485 644 645 cell_1rw
* cell instance $5608 m0 *1 148.05,30.03
X$5608 486 22 487 644 645 cell_1rw
* cell instance $5609 m0 *1 148.755,30.03
X$5609 488 22 489 644 645 cell_1rw
* cell instance $5610 m0 *1 149.46,30.03
X$5610 490 22 491 644 645 cell_1rw
* cell instance $5611 m0 *1 150.165,30.03
X$5611 492 22 493 644 645 cell_1rw
* cell instance $5612 m0 *1 150.87,30.03
X$5612 494 22 495 644 645 cell_1rw
* cell instance $5613 m0 *1 151.575,30.03
X$5613 496 22 497 644 645 cell_1rw
* cell instance $5614 m0 *1 152.28,30.03
X$5614 498 22 499 644 645 cell_1rw
* cell instance $5615 m0 *1 152.985,30.03
X$5615 500 22 501 644 645 cell_1rw
* cell instance $5616 m0 *1 153.69,30.03
X$5616 502 22 503 644 645 cell_1rw
* cell instance $5617 m0 *1 154.395,30.03
X$5617 504 22 505 644 645 cell_1rw
* cell instance $5618 m0 *1 155.1,30.03
X$5618 506 22 507 644 645 cell_1rw
* cell instance $5619 m0 *1 155.805,30.03
X$5619 508 22 509 644 645 cell_1rw
* cell instance $5620 m0 *1 156.51,30.03
X$5620 510 22 511 644 645 cell_1rw
* cell instance $5621 m0 *1 157.215,30.03
X$5621 512 22 513 644 645 cell_1rw
* cell instance $5622 m0 *1 157.92,30.03
X$5622 514 22 515 644 645 cell_1rw
* cell instance $5623 m0 *1 158.625,30.03
X$5623 516 22 517 644 645 cell_1rw
* cell instance $5624 m0 *1 159.33,30.03
X$5624 518 22 519 644 645 cell_1rw
* cell instance $5625 m0 *1 160.035,30.03
X$5625 520 22 521 644 645 cell_1rw
* cell instance $5626 m0 *1 160.74,30.03
X$5626 522 22 523 644 645 cell_1rw
* cell instance $5627 m0 *1 161.445,30.03
X$5627 524 22 525 644 645 cell_1rw
* cell instance $5628 m0 *1 162.15,30.03
X$5628 526 22 527 644 645 cell_1rw
* cell instance $5629 m0 *1 162.855,30.03
X$5629 528 22 529 644 645 cell_1rw
* cell instance $5630 m0 *1 163.56,30.03
X$5630 530 22 531 644 645 cell_1rw
* cell instance $5631 m0 *1 164.265,30.03
X$5631 532 22 533 644 645 cell_1rw
* cell instance $5632 m0 *1 164.97,30.03
X$5632 534 22 535 644 645 cell_1rw
* cell instance $5633 m0 *1 165.675,30.03
X$5633 536 22 537 644 645 cell_1rw
* cell instance $5634 m0 *1 166.38,30.03
X$5634 538 22 539 644 645 cell_1rw
* cell instance $5635 m0 *1 167.085,30.03
X$5635 540 22 541 644 645 cell_1rw
* cell instance $5636 m0 *1 167.79,30.03
X$5636 542 22 543 644 645 cell_1rw
* cell instance $5637 m0 *1 168.495,30.03
X$5637 544 22 545 644 645 cell_1rw
* cell instance $5638 m0 *1 169.2,30.03
X$5638 546 22 547 644 645 cell_1rw
* cell instance $5639 m0 *1 169.905,30.03
X$5639 548 22 549 644 645 cell_1rw
* cell instance $5640 m0 *1 170.61,30.03
X$5640 550 22 551 644 645 cell_1rw
* cell instance $5641 m0 *1 171.315,30.03
X$5641 552 22 553 644 645 cell_1rw
* cell instance $5642 m0 *1 172.02,30.03
X$5642 554 22 555 644 645 cell_1rw
* cell instance $5643 m0 *1 172.725,30.03
X$5643 556 22 557 644 645 cell_1rw
* cell instance $5644 m0 *1 173.43,30.03
X$5644 558 22 559 644 645 cell_1rw
* cell instance $5645 m0 *1 174.135,30.03
X$5645 560 22 561 644 645 cell_1rw
* cell instance $5646 m0 *1 174.84,30.03
X$5646 562 22 563 644 645 cell_1rw
* cell instance $5647 m0 *1 175.545,30.03
X$5647 564 22 565 644 645 cell_1rw
* cell instance $5648 m0 *1 176.25,30.03
X$5648 566 22 567 644 645 cell_1rw
* cell instance $5649 m0 *1 176.955,30.03
X$5649 568 22 569 644 645 cell_1rw
* cell instance $5650 m0 *1 177.66,30.03
X$5650 570 22 571 644 645 cell_1rw
* cell instance $5651 m0 *1 178.365,30.03
X$5651 572 22 573 644 645 cell_1rw
* cell instance $5652 m0 *1 179.07,30.03
X$5652 574 22 575 644 645 cell_1rw
* cell instance $5653 m0 *1 179.775,30.03
X$5653 576 22 577 644 645 cell_1rw
* cell instance $5654 m0 *1 180.48,30.03
X$5654 578 22 579 644 645 cell_1rw
* cell instance $5655 r0 *1 0.705,30.03
X$5655 67 23 68 644 645 cell_1rw
* cell instance $5656 r0 *1 0,30.03
X$5656 65 23 66 644 645 cell_1rw
* cell instance $5657 r0 *1 1.41,30.03
X$5657 69 23 70 644 645 cell_1rw
* cell instance $5658 r0 *1 2.115,30.03
X$5658 71 23 72 644 645 cell_1rw
* cell instance $5659 r0 *1 2.82,30.03
X$5659 73 23 74 644 645 cell_1rw
* cell instance $5660 r0 *1 3.525,30.03
X$5660 75 23 76 644 645 cell_1rw
* cell instance $5661 r0 *1 4.23,30.03
X$5661 77 23 78 644 645 cell_1rw
* cell instance $5662 r0 *1 4.935,30.03
X$5662 79 23 80 644 645 cell_1rw
* cell instance $5663 r0 *1 5.64,30.03
X$5663 81 23 82 644 645 cell_1rw
* cell instance $5664 r0 *1 6.345,30.03
X$5664 83 23 84 644 645 cell_1rw
* cell instance $5665 r0 *1 7.05,30.03
X$5665 85 23 86 644 645 cell_1rw
* cell instance $5666 r0 *1 7.755,30.03
X$5666 87 23 88 644 645 cell_1rw
* cell instance $5667 r0 *1 8.46,30.03
X$5667 89 23 90 644 645 cell_1rw
* cell instance $5668 r0 *1 9.165,30.03
X$5668 91 23 92 644 645 cell_1rw
* cell instance $5669 r0 *1 9.87,30.03
X$5669 93 23 94 644 645 cell_1rw
* cell instance $5670 r0 *1 10.575,30.03
X$5670 95 23 96 644 645 cell_1rw
* cell instance $5671 r0 *1 11.28,30.03
X$5671 97 23 98 644 645 cell_1rw
* cell instance $5672 r0 *1 11.985,30.03
X$5672 99 23 100 644 645 cell_1rw
* cell instance $5673 r0 *1 12.69,30.03
X$5673 101 23 102 644 645 cell_1rw
* cell instance $5674 r0 *1 13.395,30.03
X$5674 103 23 104 644 645 cell_1rw
* cell instance $5675 r0 *1 14.1,30.03
X$5675 105 23 106 644 645 cell_1rw
* cell instance $5676 r0 *1 14.805,30.03
X$5676 107 23 108 644 645 cell_1rw
* cell instance $5677 r0 *1 15.51,30.03
X$5677 109 23 110 644 645 cell_1rw
* cell instance $5678 r0 *1 16.215,30.03
X$5678 111 23 112 644 645 cell_1rw
* cell instance $5679 r0 *1 16.92,30.03
X$5679 113 23 114 644 645 cell_1rw
* cell instance $5680 r0 *1 17.625,30.03
X$5680 115 23 116 644 645 cell_1rw
* cell instance $5681 r0 *1 18.33,30.03
X$5681 117 23 118 644 645 cell_1rw
* cell instance $5682 r0 *1 19.035,30.03
X$5682 119 23 120 644 645 cell_1rw
* cell instance $5683 r0 *1 19.74,30.03
X$5683 121 23 122 644 645 cell_1rw
* cell instance $5684 r0 *1 20.445,30.03
X$5684 123 23 124 644 645 cell_1rw
* cell instance $5685 r0 *1 21.15,30.03
X$5685 125 23 126 644 645 cell_1rw
* cell instance $5686 r0 *1 21.855,30.03
X$5686 127 23 128 644 645 cell_1rw
* cell instance $5687 r0 *1 22.56,30.03
X$5687 129 23 130 644 645 cell_1rw
* cell instance $5688 r0 *1 23.265,30.03
X$5688 131 23 132 644 645 cell_1rw
* cell instance $5689 r0 *1 23.97,30.03
X$5689 133 23 134 644 645 cell_1rw
* cell instance $5690 r0 *1 24.675,30.03
X$5690 135 23 136 644 645 cell_1rw
* cell instance $5691 r0 *1 25.38,30.03
X$5691 137 23 138 644 645 cell_1rw
* cell instance $5692 r0 *1 26.085,30.03
X$5692 139 23 140 644 645 cell_1rw
* cell instance $5693 r0 *1 26.79,30.03
X$5693 141 23 142 644 645 cell_1rw
* cell instance $5694 r0 *1 27.495,30.03
X$5694 143 23 144 644 645 cell_1rw
* cell instance $5695 r0 *1 28.2,30.03
X$5695 145 23 146 644 645 cell_1rw
* cell instance $5696 r0 *1 28.905,30.03
X$5696 147 23 148 644 645 cell_1rw
* cell instance $5697 r0 *1 29.61,30.03
X$5697 149 23 150 644 645 cell_1rw
* cell instance $5698 r0 *1 30.315,30.03
X$5698 151 23 152 644 645 cell_1rw
* cell instance $5699 r0 *1 31.02,30.03
X$5699 153 23 154 644 645 cell_1rw
* cell instance $5700 r0 *1 31.725,30.03
X$5700 155 23 156 644 645 cell_1rw
* cell instance $5701 r0 *1 32.43,30.03
X$5701 157 23 158 644 645 cell_1rw
* cell instance $5702 r0 *1 33.135,30.03
X$5702 159 23 160 644 645 cell_1rw
* cell instance $5703 r0 *1 33.84,30.03
X$5703 161 23 162 644 645 cell_1rw
* cell instance $5704 r0 *1 34.545,30.03
X$5704 163 23 164 644 645 cell_1rw
* cell instance $5705 r0 *1 35.25,30.03
X$5705 165 23 166 644 645 cell_1rw
* cell instance $5706 r0 *1 35.955,30.03
X$5706 167 23 168 644 645 cell_1rw
* cell instance $5707 r0 *1 36.66,30.03
X$5707 169 23 170 644 645 cell_1rw
* cell instance $5708 r0 *1 37.365,30.03
X$5708 171 23 172 644 645 cell_1rw
* cell instance $5709 r0 *1 38.07,30.03
X$5709 173 23 174 644 645 cell_1rw
* cell instance $5710 r0 *1 38.775,30.03
X$5710 175 23 176 644 645 cell_1rw
* cell instance $5711 r0 *1 39.48,30.03
X$5711 177 23 178 644 645 cell_1rw
* cell instance $5712 r0 *1 40.185,30.03
X$5712 179 23 180 644 645 cell_1rw
* cell instance $5713 r0 *1 40.89,30.03
X$5713 181 23 182 644 645 cell_1rw
* cell instance $5714 r0 *1 41.595,30.03
X$5714 183 23 184 644 645 cell_1rw
* cell instance $5715 r0 *1 42.3,30.03
X$5715 185 23 186 644 645 cell_1rw
* cell instance $5716 r0 *1 43.005,30.03
X$5716 187 23 188 644 645 cell_1rw
* cell instance $5717 r0 *1 43.71,30.03
X$5717 189 23 190 644 645 cell_1rw
* cell instance $5718 r0 *1 44.415,30.03
X$5718 191 23 192 644 645 cell_1rw
* cell instance $5719 r0 *1 45.12,30.03
X$5719 193 23 194 644 645 cell_1rw
* cell instance $5720 r0 *1 45.825,30.03
X$5720 195 23 196 644 645 cell_1rw
* cell instance $5721 r0 *1 46.53,30.03
X$5721 197 23 198 644 645 cell_1rw
* cell instance $5722 r0 *1 47.235,30.03
X$5722 199 23 200 644 645 cell_1rw
* cell instance $5723 r0 *1 47.94,30.03
X$5723 201 23 202 644 645 cell_1rw
* cell instance $5724 r0 *1 48.645,30.03
X$5724 203 23 204 644 645 cell_1rw
* cell instance $5725 r0 *1 49.35,30.03
X$5725 205 23 206 644 645 cell_1rw
* cell instance $5726 r0 *1 50.055,30.03
X$5726 207 23 208 644 645 cell_1rw
* cell instance $5727 r0 *1 50.76,30.03
X$5727 209 23 210 644 645 cell_1rw
* cell instance $5728 r0 *1 51.465,30.03
X$5728 211 23 212 644 645 cell_1rw
* cell instance $5729 r0 *1 52.17,30.03
X$5729 213 23 214 644 645 cell_1rw
* cell instance $5730 r0 *1 52.875,30.03
X$5730 215 23 216 644 645 cell_1rw
* cell instance $5731 r0 *1 53.58,30.03
X$5731 217 23 218 644 645 cell_1rw
* cell instance $5732 r0 *1 54.285,30.03
X$5732 219 23 220 644 645 cell_1rw
* cell instance $5733 r0 *1 54.99,30.03
X$5733 221 23 222 644 645 cell_1rw
* cell instance $5734 r0 *1 55.695,30.03
X$5734 223 23 224 644 645 cell_1rw
* cell instance $5735 r0 *1 56.4,30.03
X$5735 225 23 226 644 645 cell_1rw
* cell instance $5736 r0 *1 57.105,30.03
X$5736 227 23 228 644 645 cell_1rw
* cell instance $5737 r0 *1 57.81,30.03
X$5737 229 23 230 644 645 cell_1rw
* cell instance $5738 r0 *1 58.515,30.03
X$5738 231 23 232 644 645 cell_1rw
* cell instance $5739 r0 *1 59.22,30.03
X$5739 233 23 234 644 645 cell_1rw
* cell instance $5740 r0 *1 59.925,30.03
X$5740 235 23 236 644 645 cell_1rw
* cell instance $5741 r0 *1 60.63,30.03
X$5741 237 23 238 644 645 cell_1rw
* cell instance $5742 r0 *1 61.335,30.03
X$5742 239 23 240 644 645 cell_1rw
* cell instance $5743 r0 *1 62.04,30.03
X$5743 241 23 242 644 645 cell_1rw
* cell instance $5744 r0 *1 62.745,30.03
X$5744 243 23 244 644 645 cell_1rw
* cell instance $5745 r0 *1 63.45,30.03
X$5745 245 23 246 644 645 cell_1rw
* cell instance $5746 r0 *1 64.155,30.03
X$5746 247 23 248 644 645 cell_1rw
* cell instance $5747 r0 *1 64.86,30.03
X$5747 249 23 250 644 645 cell_1rw
* cell instance $5748 r0 *1 65.565,30.03
X$5748 251 23 252 644 645 cell_1rw
* cell instance $5749 r0 *1 66.27,30.03
X$5749 253 23 254 644 645 cell_1rw
* cell instance $5750 r0 *1 66.975,30.03
X$5750 255 23 256 644 645 cell_1rw
* cell instance $5751 r0 *1 67.68,30.03
X$5751 257 23 258 644 645 cell_1rw
* cell instance $5752 r0 *1 68.385,30.03
X$5752 259 23 260 644 645 cell_1rw
* cell instance $5753 r0 *1 69.09,30.03
X$5753 261 23 262 644 645 cell_1rw
* cell instance $5754 r0 *1 69.795,30.03
X$5754 263 23 264 644 645 cell_1rw
* cell instance $5755 r0 *1 70.5,30.03
X$5755 265 23 266 644 645 cell_1rw
* cell instance $5756 r0 *1 71.205,30.03
X$5756 267 23 268 644 645 cell_1rw
* cell instance $5757 r0 *1 71.91,30.03
X$5757 269 23 270 644 645 cell_1rw
* cell instance $5758 r0 *1 72.615,30.03
X$5758 271 23 272 644 645 cell_1rw
* cell instance $5759 r0 *1 73.32,30.03
X$5759 273 23 274 644 645 cell_1rw
* cell instance $5760 r0 *1 74.025,30.03
X$5760 275 23 276 644 645 cell_1rw
* cell instance $5761 r0 *1 74.73,30.03
X$5761 277 23 278 644 645 cell_1rw
* cell instance $5762 r0 *1 75.435,30.03
X$5762 279 23 280 644 645 cell_1rw
* cell instance $5763 r0 *1 76.14,30.03
X$5763 281 23 282 644 645 cell_1rw
* cell instance $5764 r0 *1 76.845,30.03
X$5764 283 23 284 644 645 cell_1rw
* cell instance $5765 r0 *1 77.55,30.03
X$5765 285 23 286 644 645 cell_1rw
* cell instance $5766 r0 *1 78.255,30.03
X$5766 287 23 288 644 645 cell_1rw
* cell instance $5767 r0 *1 78.96,30.03
X$5767 289 23 290 644 645 cell_1rw
* cell instance $5768 r0 *1 79.665,30.03
X$5768 291 23 292 644 645 cell_1rw
* cell instance $5769 r0 *1 80.37,30.03
X$5769 293 23 294 644 645 cell_1rw
* cell instance $5770 r0 *1 81.075,30.03
X$5770 295 23 296 644 645 cell_1rw
* cell instance $5771 r0 *1 81.78,30.03
X$5771 297 23 298 644 645 cell_1rw
* cell instance $5772 r0 *1 82.485,30.03
X$5772 299 23 300 644 645 cell_1rw
* cell instance $5773 r0 *1 83.19,30.03
X$5773 301 23 302 644 645 cell_1rw
* cell instance $5774 r0 *1 83.895,30.03
X$5774 303 23 304 644 645 cell_1rw
* cell instance $5775 r0 *1 84.6,30.03
X$5775 305 23 306 644 645 cell_1rw
* cell instance $5776 r0 *1 85.305,30.03
X$5776 307 23 308 644 645 cell_1rw
* cell instance $5777 r0 *1 86.01,30.03
X$5777 309 23 310 644 645 cell_1rw
* cell instance $5778 r0 *1 86.715,30.03
X$5778 311 23 312 644 645 cell_1rw
* cell instance $5779 r0 *1 87.42,30.03
X$5779 313 23 314 644 645 cell_1rw
* cell instance $5780 r0 *1 88.125,30.03
X$5780 315 23 316 644 645 cell_1rw
* cell instance $5781 r0 *1 88.83,30.03
X$5781 317 23 318 644 645 cell_1rw
* cell instance $5782 r0 *1 89.535,30.03
X$5782 319 23 320 644 645 cell_1rw
* cell instance $5783 r0 *1 90.24,30.03
X$5783 321 23 323 644 645 cell_1rw
* cell instance $5784 r0 *1 90.945,30.03
X$5784 324 23 325 644 645 cell_1rw
* cell instance $5785 r0 *1 91.65,30.03
X$5785 326 23 327 644 645 cell_1rw
* cell instance $5786 r0 *1 92.355,30.03
X$5786 328 23 329 644 645 cell_1rw
* cell instance $5787 r0 *1 93.06,30.03
X$5787 330 23 331 644 645 cell_1rw
* cell instance $5788 r0 *1 93.765,30.03
X$5788 332 23 333 644 645 cell_1rw
* cell instance $5789 r0 *1 94.47,30.03
X$5789 334 23 335 644 645 cell_1rw
* cell instance $5790 r0 *1 95.175,30.03
X$5790 336 23 337 644 645 cell_1rw
* cell instance $5791 r0 *1 95.88,30.03
X$5791 338 23 339 644 645 cell_1rw
* cell instance $5792 r0 *1 96.585,30.03
X$5792 340 23 341 644 645 cell_1rw
* cell instance $5793 r0 *1 97.29,30.03
X$5793 342 23 343 644 645 cell_1rw
* cell instance $5794 r0 *1 97.995,30.03
X$5794 344 23 345 644 645 cell_1rw
* cell instance $5795 r0 *1 98.7,30.03
X$5795 346 23 347 644 645 cell_1rw
* cell instance $5796 r0 *1 99.405,30.03
X$5796 348 23 349 644 645 cell_1rw
* cell instance $5797 r0 *1 100.11,30.03
X$5797 350 23 351 644 645 cell_1rw
* cell instance $5798 r0 *1 100.815,30.03
X$5798 352 23 353 644 645 cell_1rw
* cell instance $5799 r0 *1 101.52,30.03
X$5799 354 23 355 644 645 cell_1rw
* cell instance $5800 r0 *1 102.225,30.03
X$5800 356 23 357 644 645 cell_1rw
* cell instance $5801 r0 *1 102.93,30.03
X$5801 358 23 359 644 645 cell_1rw
* cell instance $5802 r0 *1 103.635,30.03
X$5802 360 23 361 644 645 cell_1rw
* cell instance $5803 r0 *1 104.34,30.03
X$5803 362 23 363 644 645 cell_1rw
* cell instance $5804 r0 *1 105.045,30.03
X$5804 364 23 365 644 645 cell_1rw
* cell instance $5805 r0 *1 105.75,30.03
X$5805 366 23 367 644 645 cell_1rw
* cell instance $5806 r0 *1 106.455,30.03
X$5806 368 23 369 644 645 cell_1rw
* cell instance $5807 r0 *1 107.16,30.03
X$5807 370 23 371 644 645 cell_1rw
* cell instance $5808 r0 *1 107.865,30.03
X$5808 372 23 373 644 645 cell_1rw
* cell instance $5809 r0 *1 108.57,30.03
X$5809 374 23 375 644 645 cell_1rw
* cell instance $5810 r0 *1 109.275,30.03
X$5810 376 23 377 644 645 cell_1rw
* cell instance $5811 r0 *1 109.98,30.03
X$5811 378 23 379 644 645 cell_1rw
* cell instance $5812 r0 *1 110.685,30.03
X$5812 380 23 381 644 645 cell_1rw
* cell instance $5813 r0 *1 111.39,30.03
X$5813 382 23 383 644 645 cell_1rw
* cell instance $5814 r0 *1 112.095,30.03
X$5814 384 23 385 644 645 cell_1rw
* cell instance $5815 r0 *1 112.8,30.03
X$5815 386 23 387 644 645 cell_1rw
* cell instance $5816 r0 *1 113.505,30.03
X$5816 388 23 389 644 645 cell_1rw
* cell instance $5817 r0 *1 114.21,30.03
X$5817 390 23 391 644 645 cell_1rw
* cell instance $5818 r0 *1 114.915,30.03
X$5818 392 23 393 644 645 cell_1rw
* cell instance $5819 r0 *1 115.62,30.03
X$5819 394 23 395 644 645 cell_1rw
* cell instance $5820 r0 *1 116.325,30.03
X$5820 396 23 397 644 645 cell_1rw
* cell instance $5821 r0 *1 117.03,30.03
X$5821 398 23 399 644 645 cell_1rw
* cell instance $5822 r0 *1 117.735,30.03
X$5822 400 23 401 644 645 cell_1rw
* cell instance $5823 r0 *1 118.44,30.03
X$5823 402 23 403 644 645 cell_1rw
* cell instance $5824 r0 *1 119.145,30.03
X$5824 404 23 405 644 645 cell_1rw
* cell instance $5825 r0 *1 119.85,30.03
X$5825 406 23 407 644 645 cell_1rw
* cell instance $5826 r0 *1 120.555,30.03
X$5826 408 23 409 644 645 cell_1rw
* cell instance $5827 r0 *1 121.26,30.03
X$5827 410 23 411 644 645 cell_1rw
* cell instance $5828 r0 *1 121.965,30.03
X$5828 412 23 413 644 645 cell_1rw
* cell instance $5829 r0 *1 122.67,30.03
X$5829 414 23 415 644 645 cell_1rw
* cell instance $5830 r0 *1 123.375,30.03
X$5830 416 23 417 644 645 cell_1rw
* cell instance $5831 r0 *1 124.08,30.03
X$5831 418 23 419 644 645 cell_1rw
* cell instance $5832 r0 *1 124.785,30.03
X$5832 420 23 421 644 645 cell_1rw
* cell instance $5833 r0 *1 125.49,30.03
X$5833 422 23 423 644 645 cell_1rw
* cell instance $5834 r0 *1 126.195,30.03
X$5834 424 23 425 644 645 cell_1rw
* cell instance $5835 r0 *1 126.9,30.03
X$5835 426 23 427 644 645 cell_1rw
* cell instance $5836 r0 *1 127.605,30.03
X$5836 428 23 429 644 645 cell_1rw
* cell instance $5837 r0 *1 128.31,30.03
X$5837 430 23 431 644 645 cell_1rw
* cell instance $5838 r0 *1 129.015,30.03
X$5838 432 23 433 644 645 cell_1rw
* cell instance $5839 r0 *1 129.72,30.03
X$5839 434 23 435 644 645 cell_1rw
* cell instance $5840 r0 *1 130.425,30.03
X$5840 436 23 437 644 645 cell_1rw
* cell instance $5841 r0 *1 131.13,30.03
X$5841 438 23 439 644 645 cell_1rw
* cell instance $5842 r0 *1 131.835,30.03
X$5842 440 23 441 644 645 cell_1rw
* cell instance $5843 r0 *1 132.54,30.03
X$5843 442 23 443 644 645 cell_1rw
* cell instance $5844 r0 *1 133.245,30.03
X$5844 444 23 445 644 645 cell_1rw
* cell instance $5845 r0 *1 133.95,30.03
X$5845 446 23 447 644 645 cell_1rw
* cell instance $5846 r0 *1 134.655,30.03
X$5846 448 23 449 644 645 cell_1rw
* cell instance $5847 r0 *1 135.36,30.03
X$5847 450 23 451 644 645 cell_1rw
* cell instance $5848 r0 *1 136.065,30.03
X$5848 452 23 453 644 645 cell_1rw
* cell instance $5849 r0 *1 136.77,30.03
X$5849 454 23 455 644 645 cell_1rw
* cell instance $5850 r0 *1 137.475,30.03
X$5850 456 23 457 644 645 cell_1rw
* cell instance $5851 r0 *1 138.18,30.03
X$5851 458 23 459 644 645 cell_1rw
* cell instance $5852 r0 *1 138.885,30.03
X$5852 460 23 461 644 645 cell_1rw
* cell instance $5853 r0 *1 139.59,30.03
X$5853 462 23 463 644 645 cell_1rw
* cell instance $5854 r0 *1 140.295,30.03
X$5854 464 23 465 644 645 cell_1rw
* cell instance $5855 r0 *1 141,30.03
X$5855 466 23 467 644 645 cell_1rw
* cell instance $5856 r0 *1 141.705,30.03
X$5856 468 23 469 644 645 cell_1rw
* cell instance $5857 r0 *1 142.41,30.03
X$5857 470 23 471 644 645 cell_1rw
* cell instance $5858 r0 *1 143.115,30.03
X$5858 472 23 473 644 645 cell_1rw
* cell instance $5859 r0 *1 143.82,30.03
X$5859 474 23 475 644 645 cell_1rw
* cell instance $5860 r0 *1 144.525,30.03
X$5860 476 23 477 644 645 cell_1rw
* cell instance $5861 r0 *1 145.23,30.03
X$5861 478 23 479 644 645 cell_1rw
* cell instance $5862 r0 *1 145.935,30.03
X$5862 480 23 481 644 645 cell_1rw
* cell instance $5863 r0 *1 146.64,30.03
X$5863 482 23 483 644 645 cell_1rw
* cell instance $5864 r0 *1 147.345,30.03
X$5864 484 23 485 644 645 cell_1rw
* cell instance $5865 r0 *1 148.05,30.03
X$5865 486 23 487 644 645 cell_1rw
* cell instance $5866 r0 *1 148.755,30.03
X$5866 488 23 489 644 645 cell_1rw
* cell instance $5867 r0 *1 149.46,30.03
X$5867 490 23 491 644 645 cell_1rw
* cell instance $5868 r0 *1 150.165,30.03
X$5868 492 23 493 644 645 cell_1rw
* cell instance $5869 r0 *1 150.87,30.03
X$5869 494 23 495 644 645 cell_1rw
* cell instance $5870 r0 *1 151.575,30.03
X$5870 496 23 497 644 645 cell_1rw
* cell instance $5871 r0 *1 152.28,30.03
X$5871 498 23 499 644 645 cell_1rw
* cell instance $5872 r0 *1 152.985,30.03
X$5872 500 23 501 644 645 cell_1rw
* cell instance $5873 r0 *1 153.69,30.03
X$5873 502 23 503 644 645 cell_1rw
* cell instance $5874 r0 *1 154.395,30.03
X$5874 504 23 505 644 645 cell_1rw
* cell instance $5875 r0 *1 155.1,30.03
X$5875 506 23 507 644 645 cell_1rw
* cell instance $5876 r0 *1 155.805,30.03
X$5876 508 23 509 644 645 cell_1rw
* cell instance $5877 r0 *1 156.51,30.03
X$5877 510 23 511 644 645 cell_1rw
* cell instance $5878 r0 *1 157.215,30.03
X$5878 512 23 513 644 645 cell_1rw
* cell instance $5879 r0 *1 157.92,30.03
X$5879 514 23 515 644 645 cell_1rw
* cell instance $5880 r0 *1 158.625,30.03
X$5880 516 23 517 644 645 cell_1rw
* cell instance $5881 r0 *1 159.33,30.03
X$5881 518 23 519 644 645 cell_1rw
* cell instance $5882 r0 *1 160.035,30.03
X$5882 520 23 521 644 645 cell_1rw
* cell instance $5883 r0 *1 160.74,30.03
X$5883 522 23 523 644 645 cell_1rw
* cell instance $5884 r0 *1 161.445,30.03
X$5884 524 23 525 644 645 cell_1rw
* cell instance $5885 r0 *1 162.15,30.03
X$5885 526 23 527 644 645 cell_1rw
* cell instance $5886 r0 *1 162.855,30.03
X$5886 528 23 529 644 645 cell_1rw
* cell instance $5887 r0 *1 163.56,30.03
X$5887 530 23 531 644 645 cell_1rw
* cell instance $5888 r0 *1 164.265,30.03
X$5888 532 23 533 644 645 cell_1rw
* cell instance $5889 r0 *1 164.97,30.03
X$5889 534 23 535 644 645 cell_1rw
* cell instance $5890 r0 *1 165.675,30.03
X$5890 536 23 537 644 645 cell_1rw
* cell instance $5891 r0 *1 166.38,30.03
X$5891 538 23 539 644 645 cell_1rw
* cell instance $5892 r0 *1 167.085,30.03
X$5892 540 23 541 644 645 cell_1rw
* cell instance $5893 r0 *1 167.79,30.03
X$5893 542 23 543 644 645 cell_1rw
* cell instance $5894 r0 *1 168.495,30.03
X$5894 544 23 545 644 645 cell_1rw
* cell instance $5895 r0 *1 169.2,30.03
X$5895 546 23 547 644 645 cell_1rw
* cell instance $5896 r0 *1 169.905,30.03
X$5896 548 23 549 644 645 cell_1rw
* cell instance $5897 r0 *1 170.61,30.03
X$5897 550 23 551 644 645 cell_1rw
* cell instance $5898 r0 *1 171.315,30.03
X$5898 552 23 553 644 645 cell_1rw
* cell instance $5899 r0 *1 172.02,30.03
X$5899 554 23 555 644 645 cell_1rw
* cell instance $5900 r0 *1 172.725,30.03
X$5900 556 23 557 644 645 cell_1rw
* cell instance $5901 r0 *1 173.43,30.03
X$5901 558 23 559 644 645 cell_1rw
* cell instance $5902 r0 *1 174.135,30.03
X$5902 560 23 561 644 645 cell_1rw
* cell instance $5903 r0 *1 174.84,30.03
X$5903 562 23 563 644 645 cell_1rw
* cell instance $5904 r0 *1 175.545,30.03
X$5904 564 23 565 644 645 cell_1rw
* cell instance $5905 r0 *1 176.25,30.03
X$5905 566 23 567 644 645 cell_1rw
* cell instance $5906 r0 *1 176.955,30.03
X$5906 568 23 569 644 645 cell_1rw
* cell instance $5907 r0 *1 177.66,30.03
X$5907 570 23 571 644 645 cell_1rw
* cell instance $5908 r0 *1 178.365,30.03
X$5908 572 23 573 644 645 cell_1rw
* cell instance $5909 r0 *1 179.07,30.03
X$5909 574 23 575 644 645 cell_1rw
* cell instance $5910 r0 *1 179.775,30.03
X$5910 576 23 577 644 645 cell_1rw
* cell instance $5911 r0 *1 180.48,30.03
X$5911 578 23 579 644 645 cell_1rw
* cell instance $5912 m0 *1 0.705,32.76
X$5912 67 24 68 644 645 cell_1rw
* cell instance $5913 m0 *1 0,32.76
X$5913 65 24 66 644 645 cell_1rw
* cell instance $5914 m0 *1 1.41,32.76
X$5914 69 24 70 644 645 cell_1rw
* cell instance $5915 m0 *1 2.115,32.76
X$5915 71 24 72 644 645 cell_1rw
* cell instance $5916 m0 *1 2.82,32.76
X$5916 73 24 74 644 645 cell_1rw
* cell instance $5917 m0 *1 3.525,32.76
X$5917 75 24 76 644 645 cell_1rw
* cell instance $5918 m0 *1 4.23,32.76
X$5918 77 24 78 644 645 cell_1rw
* cell instance $5919 m0 *1 4.935,32.76
X$5919 79 24 80 644 645 cell_1rw
* cell instance $5920 m0 *1 5.64,32.76
X$5920 81 24 82 644 645 cell_1rw
* cell instance $5921 m0 *1 6.345,32.76
X$5921 83 24 84 644 645 cell_1rw
* cell instance $5922 m0 *1 7.05,32.76
X$5922 85 24 86 644 645 cell_1rw
* cell instance $5923 m0 *1 7.755,32.76
X$5923 87 24 88 644 645 cell_1rw
* cell instance $5924 m0 *1 8.46,32.76
X$5924 89 24 90 644 645 cell_1rw
* cell instance $5925 m0 *1 9.165,32.76
X$5925 91 24 92 644 645 cell_1rw
* cell instance $5926 m0 *1 9.87,32.76
X$5926 93 24 94 644 645 cell_1rw
* cell instance $5927 m0 *1 10.575,32.76
X$5927 95 24 96 644 645 cell_1rw
* cell instance $5928 m0 *1 11.28,32.76
X$5928 97 24 98 644 645 cell_1rw
* cell instance $5929 m0 *1 11.985,32.76
X$5929 99 24 100 644 645 cell_1rw
* cell instance $5930 m0 *1 12.69,32.76
X$5930 101 24 102 644 645 cell_1rw
* cell instance $5931 m0 *1 13.395,32.76
X$5931 103 24 104 644 645 cell_1rw
* cell instance $5932 m0 *1 14.1,32.76
X$5932 105 24 106 644 645 cell_1rw
* cell instance $5933 m0 *1 14.805,32.76
X$5933 107 24 108 644 645 cell_1rw
* cell instance $5934 m0 *1 15.51,32.76
X$5934 109 24 110 644 645 cell_1rw
* cell instance $5935 m0 *1 16.215,32.76
X$5935 111 24 112 644 645 cell_1rw
* cell instance $5936 m0 *1 16.92,32.76
X$5936 113 24 114 644 645 cell_1rw
* cell instance $5937 m0 *1 17.625,32.76
X$5937 115 24 116 644 645 cell_1rw
* cell instance $5938 m0 *1 18.33,32.76
X$5938 117 24 118 644 645 cell_1rw
* cell instance $5939 m0 *1 19.035,32.76
X$5939 119 24 120 644 645 cell_1rw
* cell instance $5940 m0 *1 19.74,32.76
X$5940 121 24 122 644 645 cell_1rw
* cell instance $5941 m0 *1 20.445,32.76
X$5941 123 24 124 644 645 cell_1rw
* cell instance $5942 m0 *1 21.15,32.76
X$5942 125 24 126 644 645 cell_1rw
* cell instance $5943 m0 *1 21.855,32.76
X$5943 127 24 128 644 645 cell_1rw
* cell instance $5944 m0 *1 22.56,32.76
X$5944 129 24 130 644 645 cell_1rw
* cell instance $5945 m0 *1 23.265,32.76
X$5945 131 24 132 644 645 cell_1rw
* cell instance $5946 m0 *1 23.97,32.76
X$5946 133 24 134 644 645 cell_1rw
* cell instance $5947 m0 *1 24.675,32.76
X$5947 135 24 136 644 645 cell_1rw
* cell instance $5948 m0 *1 25.38,32.76
X$5948 137 24 138 644 645 cell_1rw
* cell instance $5949 m0 *1 26.085,32.76
X$5949 139 24 140 644 645 cell_1rw
* cell instance $5950 m0 *1 26.79,32.76
X$5950 141 24 142 644 645 cell_1rw
* cell instance $5951 m0 *1 27.495,32.76
X$5951 143 24 144 644 645 cell_1rw
* cell instance $5952 m0 *1 28.2,32.76
X$5952 145 24 146 644 645 cell_1rw
* cell instance $5953 m0 *1 28.905,32.76
X$5953 147 24 148 644 645 cell_1rw
* cell instance $5954 m0 *1 29.61,32.76
X$5954 149 24 150 644 645 cell_1rw
* cell instance $5955 m0 *1 30.315,32.76
X$5955 151 24 152 644 645 cell_1rw
* cell instance $5956 m0 *1 31.02,32.76
X$5956 153 24 154 644 645 cell_1rw
* cell instance $5957 m0 *1 31.725,32.76
X$5957 155 24 156 644 645 cell_1rw
* cell instance $5958 m0 *1 32.43,32.76
X$5958 157 24 158 644 645 cell_1rw
* cell instance $5959 m0 *1 33.135,32.76
X$5959 159 24 160 644 645 cell_1rw
* cell instance $5960 m0 *1 33.84,32.76
X$5960 161 24 162 644 645 cell_1rw
* cell instance $5961 m0 *1 34.545,32.76
X$5961 163 24 164 644 645 cell_1rw
* cell instance $5962 m0 *1 35.25,32.76
X$5962 165 24 166 644 645 cell_1rw
* cell instance $5963 m0 *1 35.955,32.76
X$5963 167 24 168 644 645 cell_1rw
* cell instance $5964 m0 *1 36.66,32.76
X$5964 169 24 170 644 645 cell_1rw
* cell instance $5965 m0 *1 37.365,32.76
X$5965 171 24 172 644 645 cell_1rw
* cell instance $5966 m0 *1 38.07,32.76
X$5966 173 24 174 644 645 cell_1rw
* cell instance $5967 m0 *1 38.775,32.76
X$5967 175 24 176 644 645 cell_1rw
* cell instance $5968 m0 *1 39.48,32.76
X$5968 177 24 178 644 645 cell_1rw
* cell instance $5969 m0 *1 40.185,32.76
X$5969 179 24 180 644 645 cell_1rw
* cell instance $5970 m0 *1 40.89,32.76
X$5970 181 24 182 644 645 cell_1rw
* cell instance $5971 m0 *1 41.595,32.76
X$5971 183 24 184 644 645 cell_1rw
* cell instance $5972 m0 *1 42.3,32.76
X$5972 185 24 186 644 645 cell_1rw
* cell instance $5973 m0 *1 43.005,32.76
X$5973 187 24 188 644 645 cell_1rw
* cell instance $5974 m0 *1 43.71,32.76
X$5974 189 24 190 644 645 cell_1rw
* cell instance $5975 m0 *1 44.415,32.76
X$5975 191 24 192 644 645 cell_1rw
* cell instance $5976 m0 *1 45.12,32.76
X$5976 193 24 194 644 645 cell_1rw
* cell instance $5977 m0 *1 45.825,32.76
X$5977 195 24 196 644 645 cell_1rw
* cell instance $5978 m0 *1 46.53,32.76
X$5978 197 24 198 644 645 cell_1rw
* cell instance $5979 m0 *1 47.235,32.76
X$5979 199 24 200 644 645 cell_1rw
* cell instance $5980 m0 *1 47.94,32.76
X$5980 201 24 202 644 645 cell_1rw
* cell instance $5981 m0 *1 48.645,32.76
X$5981 203 24 204 644 645 cell_1rw
* cell instance $5982 m0 *1 49.35,32.76
X$5982 205 24 206 644 645 cell_1rw
* cell instance $5983 m0 *1 50.055,32.76
X$5983 207 24 208 644 645 cell_1rw
* cell instance $5984 m0 *1 50.76,32.76
X$5984 209 24 210 644 645 cell_1rw
* cell instance $5985 m0 *1 51.465,32.76
X$5985 211 24 212 644 645 cell_1rw
* cell instance $5986 m0 *1 52.17,32.76
X$5986 213 24 214 644 645 cell_1rw
* cell instance $5987 m0 *1 52.875,32.76
X$5987 215 24 216 644 645 cell_1rw
* cell instance $5988 m0 *1 53.58,32.76
X$5988 217 24 218 644 645 cell_1rw
* cell instance $5989 m0 *1 54.285,32.76
X$5989 219 24 220 644 645 cell_1rw
* cell instance $5990 m0 *1 54.99,32.76
X$5990 221 24 222 644 645 cell_1rw
* cell instance $5991 m0 *1 55.695,32.76
X$5991 223 24 224 644 645 cell_1rw
* cell instance $5992 m0 *1 56.4,32.76
X$5992 225 24 226 644 645 cell_1rw
* cell instance $5993 m0 *1 57.105,32.76
X$5993 227 24 228 644 645 cell_1rw
* cell instance $5994 m0 *1 57.81,32.76
X$5994 229 24 230 644 645 cell_1rw
* cell instance $5995 m0 *1 58.515,32.76
X$5995 231 24 232 644 645 cell_1rw
* cell instance $5996 m0 *1 59.22,32.76
X$5996 233 24 234 644 645 cell_1rw
* cell instance $5997 m0 *1 59.925,32.76
X$5997 235 24 236 644 645 cell_1rw
* cell instance $5998 m0 *1 60.63,32.76
X$5998 237 24 238 644 645 cell_1rw
* cell instance $5999 m0 *1 61.335,32.76
X$5999 239 24 240 644 645 cell_1rw
* cell instance $6000 m0 *1 62.04,32.76
X$6000 241 24 242 644 645 cell_1rw
* cell instance $6001 m0 *1 62.745,32.76
X$6001 243 24 244 644 645 cell_1rw
* cell instance $6002 m0 *1 63.45,32.76
X$6002 245 24 246 644 645 cell_1rw
* cell instance $6003 m0 *1 64.155,32.76
X$6003 247 24 248 644 645 cell_1rw
* cell instance $6004 m0 *1 64.86,32.76
X$6004 249 24 250 644 645 cell_1rw
* cell instance $6005 m0 *1 65.565,32.76
X$6005 251 24 252 644 645 cell_1rw
* cell instance $6006 m0 *1 66.27,32.76
X$6006 253 24 254 644 645 cell_1rw
* cell instance $6007 m0 *1 66.975,32.76
X$6007 255 24 256 644 645 cell_1rw
* cell instance $6008 m0 *1 67.68,32.76
X$6008 257 24 258 644 645 cell_1rw
* cell instance $6009 m0 *1 68.385,32.76
X$6009 259 24 260 644 645 cell_1rw
* cell instance $6010 m0 *1 69.09,32.76
X$6010 261 24 262 644 645 cell_1rw
* cell instance $6011 m0 *1 69.795,32.76
X$6011 263 24 264 644 645 cell_1rw
* cell instance $6012 m0 *1 70.5,32.76
X$6012 265 24 266 644 645 cell_1rw
* cell instance $6013 m0 *1 71.205,32.76
X$6013 267 24 268 644 645 cell_1rw
* cell instance $6014 m0 *1 71.91,32.76
X$6014 269 24 270 644 645 cell_1rw
* cell instance $6015 m0 *1 72.615,32.76
X$6015 271 24 272 644 645 cell_1rw
* cell instance $6016 m0 *1 73.32,32.76
X$6016 273 24 274 644 645 cell_1rw
* cell instance $6017 m0 *1 74.025,32.76
X$6017 275 24 276 644 645 cell_1rw
* cell instance $6018 m0 *1 74.73,32.76
X$6018 277 24 278 644 645 cell_1rw
* cell instance $6019 m0 *1 75.435,32.76
X$6019 279 24 280 644 645 cell_1rw
* cell instance $6020 m0 *1 76.14,32.76
X$6020 281 24 282 644 645 cell_1rw
* cell instance $6021 m0 *1 76.845,32.76
X$6021 283 24 284 644 645 cell_1rw
* cell instance $6022 m0 *1 77.55,32.76
X$6022 285 24 286 644 645 cell_1rw
* cell instance $6023 m0 *1 78.255,32.76
X$6023 287 24 288 644 645 cell_1rw
* cell instance $6024 m0 *1 78.96,32.76
X$6024 289 24 290 644 645 cell_1rw
* cell instance $6025 m0 *1 79.665,32.76
X$6025 291 24 292 644 645 cell_1rw
* cell instance $6026 m0 *1 80.37,32.76
X$6026 293 24 294 644 645 cell_1rw
* cell instance $6027 m0 *1 81.075,32.76
X$6027 295 24 296 644 645 cell_1rw
* cell instance $6028 m0 *1 81.78,32.76
X$6028 297 24 298 644 645 cell_1rw
* cell instance $6029 m0 *1 82.485,32.76
X$6029 299 24 300 644 645 cell_1rw
* cell instance $6030 m0 *1 83.19,32.76
X$6030 301 24 302 644 645 cell_1rw
* cell instance $6031 m0 *1 83.895,32.76
X$6031 303 24 304 644 645 cell_1rw
* cell instance $6032 m0 *1 84.6,32.76
X$6032 305 24 306 644 645 cell_1rw
* cell instance $6033 m0 *1 85.305,32.76
X$6033 307 24 308 644 645 cell_1rw
* cell instance $6034 m0 *1 86.01,32.76
X$6034 309 24 310 644 645 cell_1rw
* cell instance $6035 m0 *1 86.715,32.76
X$6035 311 24 312 644 645 cell_1rw
* cell instance $6036 m0 *1 87.42,32.76
X$6036 313 24 314 644 645 cell_1rw
* cell instance $6037 m0 *1 88.125,32.76
X$6037 315 24 316 644 645 cell_1rw
* cell instance $6038 m0 *1 88.83,32.76
X$6038 317 24 318 644 645 cell_1rw
* cell instance $6039 m0 *1 89.535,32.76
X$6039 319 24 320 644 645 cell_1rw
* cell instance $6040 m0 *1 90.24,32.76
X$6040 321 24 323 644 645 cell_1rw
* cell instance $6041 m0 *1 90.945,32.76
X$6041 324 24 325 644 645 cell_1rw
* cell instance $6042 m0 *1 91.65,32.76
X$6042 326 24 327 644 645 cell_1rw
* cell instance $6043 m0 *1 92.355,32.76
X$6043 328 24 329 644 645 cell_1rw
* cell instance $6044 m0 *1 93.06,32.76
X$6044 330 24 331 644 645 cell_1rw
* cell instance $6045 m0 *1 93.765,32.76
X$6045 332 24 333 644 645 cell_1rw
* cell instance $6046 m0 *1 94.47,32.76
X$6046 334 24 335 644 645 cell_1rw
* cell instance $6047 m0 *1 95.175,32.76
X$6047 336 24 337 644 645 cell_1rw
* cell instance $6048 m0 *1 95.88,32.76
X$6048 338 24 339 644 645 cell_1rw
* cell instance $6049 m0 *1 96.585,32.76
X$6049 340 24 341 644 645 cell_1rw
* cell instance $6050 m0 *1 97.29,32.76
X$6050 342 24 343 644 645 cell_1rw
* cell instance $6051 m0 *1 97.995,32.76
X$6051 344 24 345 644 645 cell_1rw
* cell instance $6052 m0 *1 98.7,32.76
X$6052 346 24 347 644 645 cell_1rw
* cell instance $6053 m0 *1 99.405,32.76
X$6053 348 24 349 644 645 cell_1rw
* cell instance $6054 m0 *1 100.11,32.76
X$6054 350 24 351 644 645 cell_1rw
* cell instance $6055 m0 *1 100.815,32.76
X$6055 352 24 353 644 645 cell_1rw
* cell instance $6056 m0 *1 101.52,32.76
X$6056 354 24 355 644 645 cell_1rw
* cell instance $6057 m0 *1 102.225,32.76
X$6057 356 24 357 644 645 cell_1rw
* cell instance $6058 m0 *1 102.93,32.76
X$6058 358 24 359 644 645 cell_1rw
* cell instance $6059 m0 *1 103.635,32.76
X$6059 360 24 361 644 645 cell_1rw
* cell instance $6060 m0 *1 104.34,32.76
X$6060 362 24 363 644 645 cell_1rw
* cell instance $6061 m0 *1 105.045,32.76
X$6061 364 24 365 644 645 cell_1rw
* cell instance $6062 m0 *1 105.75,32.76
X$6062 366 24 367 644 645 cell_1rw
* cell instance $6063 m0 *1 106.455,32.76
X$6063 368 24 369 644 645 cell_1rw
* cell instance $6064 m0 *1 107.16,32.76
X$6064 370 24 371 644 645 cell_1rw
* cell instance $6065 m0 *1 107.865,32.76
X$6065 372 24 373 644 645 cell_1rw
* cell instance $6066 m0 *1 108.57,32.76
X$6066 374 24 375 644 645 cell_1rw
* cell instance $6067 m0 *1 109.275,32.76
X$6067 376 24 377 644 645 cell_1rw
* cell instance $6068 m0 *1 109.98,32.76
X$6068 378 24 379 644 645 cell_1rw
* cell instance $6069 m0 *1 110.685,32.76
X$6069 380 24 381 644 645 cell_1rw
* cell instance $6070 m0 *1 111.39,32.76
X$6070 382 24 383 644 645 cell_1rw
* cell instance $6071 m0 *1 112.095,32.76
X$6071 384 24 385 644 645 cell_1rw
* cell instance $6072 m0 *1 112.8,32.76
X$6072 386 24 387 644 645 cell_1rw
* cell instance $6073 m0 *1 113.505,32.76
X$6073 388 24 389 644 645 cell_1rw
* cell instance $6074 m0 *1 114.21,32.76
X$6074 390 24 391 644 645 cell_1rw
* cell instance $6075 m0 *1 114.915,32.76
X$6075 392 24 393 644 645 cell_1rw
* cell instance $6076 m0 *1 115.62,32.76
X$6076 394 24 395 644 645 cell_1rw
* cell instance $6077 m0 *1 116.325,32.76
X$6077 396 24 397 644 645 cell_1rw
* cell instance $6078 m0 *1 117.03,32.76
X$6078 398 24 399 644 645 cell_1rw
* cell instance $6079 m0 *1 117.735,32.76
X$6079 400 24 401 644 645 cell_1rw
* cell instance $6080 m0 *1 118.44,32.76
X$6080 402 24 403 644 645 cell_1rw
* cell instance $6081 m0 *1 119.145,32.76
X$6081 404 24 405 644 645 cell_1rw
* cell instance $6082 m0 *1 119.85,32.76
X$6082 406 24 407 644 645 cell_1rw
* cell instance $6083 m0 *1 120.555,32.76
X$6083 408 24 409 644 645 cell_1rw
* cell instance $6084 m0 *1 121.26,32.76
X$6084 410 24 411 644 645 cell_1rw
* cell instance $6085 m0 *1 121.965,32.76
X$6085 412 24 413 644 645 cell_1rw
* cell instance $6086 m0 *1 122.67,32.76
X$6086 414 24 415 644 645 cell_1rw
* cell instance $6087 m0 *1 123.375,32.76
X$6087 416 24 417 644 645 cell_1rw
* cell instance $6088 m0 *1 124.08,32.76
X$6088 418 24 419 644 645 cell_1rw
* cell instance $6089 m0 *1 124.785,32.76
X$6089 420 24 421 644 645 cell_1rw
* cell instance $6090 m0 *1 125.49,32.76
X$6090 422 24 423 644 645 cell_1rw
* cell instance $6091 m0 *1 126.195,32.76
X$6091 424 24 425 644 645 cell_1rw
* cell instance $6092 m0 *1 126.9,32.76
X$6092 426 24 427 644 645 cell_1rw
* cell instance $6093 m0 *1 127.605,32.76
X$6093 428 24 429 644 645 cell_1rw
* cell instance $6094 m0 *1 128.31,32.76
X$6094 430 24 431 644 645 cell_1rw
* cell instance $6095 m0 *1 129.015,32.76
X$6095 432 24 433 644 645 cell_1rw
* cell instance $6096 m0 *1 129.72,32.76
X$6096 434 24 435 644 645 cell_1rw
* cell instance $6097 m0 *1 130.425,32.76
X$6097 436 24 437 644 645 cell_1rw
* cell instance $6098 m0 *1 131.13,32.76
X$6098 438 24 439 644 645 cell_1rw
* cell instance $6099 m0 *1 131.835,32.76
X$6099 440 24 441 644 645 cell_1rw
* cell instance $6100 m0 *1 132.54,32.76
X$6100 442 24 443 644 645 cell_1rw
* cell instance $6101 m0 *1 133.245,32.76
X$6101 444 24 445 644 645 cell_1rw
* cell instance $6102 m0 *1 133.95,32.76
X$6102 446 24 447 644 645 cell_1rw
* cell instance $6103 m0 *1 134.655,32.76
X$6103 448 24 449 644 645 cell_1rw
* cell instance $6104 m0 *1 135.36,32.76
X$6104 450 24 451 644 645 cell_1rw
* cell instance $6105 m0 *1 136.065,32.76
X$6105 452 24 453 644 645 cell_1rw
* cell instance $6106 m0 *1 136.77,32.76
X$6106 454 24 455 644 645 cell_1rw
* cell instance $6107 m0 *1 137.475,32.76
X$6107 456 24 457 644 645 cell_1rw
* cell instance $6108 m0 *1 138.18,32.76
X$6108 458 24 459 644 645 cell_1rw
* cell instance $6109 m0 *1 138.885,32.76
X$6109 460 24 461 644 645 cell_1rw
* cell instance $6110 m0 *1 139.59,32.76
X$6110 462 24 463 644 645 cell_1rw
* cell instance $6111 m0 *1 140.295,32.76
X$6111 464 24 465 644 645 cell_1rw
* cell instance $6112 m0 *1 141,32.76
X$6112 466 24 467 644 645 cell_1rw
* cell instance $6113 m0 *1 141.705,32.76
X$6113 468 24 469 644 645 cell_1rw
* cell instance $6114 m0 *1 142.41,32.76
X$6114 470 24 471 644 645 cell_1rw
* cell instance $6115 m0 *1 143.115,32.76
X$6115 472 24 473 644 645 cell_1rw
* cell instance $6116 m0 *1 143.82,32.76
X$6116 474 24 475 644 645 cell_1rw
* cell instance $6117 m0 *1 144.525,32.76
X$6117 476 24 477 644 645 cell_1rw
* cell instance $6118 m0 *1 145.23,32.76
X$6118 478 24 479 644 645 cell_1rw
* cell instance $6119 m0 *1 145.935,32.76
X$6119 480 24 481 644 645 cell_1rw
* cell instance $6120 m0 *1 146.64,32.76
X$6120 482 24 483 644 645 cell_1rw
* cell instance $6121 m0 *1 147.345,32.76
X$6121 484 24 485 644 645 cell_1rw
* cell instance $6122 m0 *1 148.05,32.76
X$6122 486 24 487 644 645 cell_1rw
* cell instance $6123 m0 *1 148.755,32.76
X$6123 488 24 489 644 645 cell_1rw
* cell instance $6124 m0 *1 149.46,32.76
X$6124 490 24 491 644 645 cell_1rw
* cell instance $6125 m0 *1 150.165,32.76
X$6125 492 24 493 644 645 cell_1rw
* cell instance $6126 m0 *1 150.87,32.76
X$6126 494 24 495 644 645 cell_1rw
* cell instance $6127 m0 *1 151.575,32.76
X$6127 496 24 497 644 645 cell_1rw
* cell instance $6128 m0 *1 152.28,32.76
X$6128 498 24 499 644 645 cell_1rw
* cell instance $6129 m0 *1 152.985,32.76
X$6129 500 24 501 644 645 cell_1rw
* cell instance $6130 m0 *1 153.69,32.76
X$6130 502 24 503 644 645 cell_1rw
* cell instance $6131 m0 *1 154.395,32.76
X$6131 504 24 505 644 645 cell_1rw
* cell instance $6132 m0 *1 155.1,32.76
X$6132 506 24 507 644 645 cell_1rw
* cell instance $6133 m0 *1 155.805,32.76
X$6133 508 24 509 644 645 cell_1rw
* cell instance $6134 m0 *1 156.51,32.76
X$6134 510 24 511 644 645 cell_1rw
* cell instance $6135 m0 *1 157.215,32.76
X$6135 512 24 513 644 645 cell_1rw
* cell instance $6136 m0 *1 157.92,32.76
X$6136 514 24 515 644 645 cell_1rw
* cell instance $6137 m0 *1 158.625,32.76
X$6137 516 24 517 644 645 cell_1rw
* cell instance $6138 m0 *1 159.33,32.76
X$6138 518 24 519 644 645 cell_1rw
* cell instance $6139 m0 *1 160.035,32.76
X$6139 520 24 521 644 645 cell_1rw
* cell instance $6140 m0 *1 160.74,32.76
X$6140 522 24 523 644 645 cell_1rw
* cell instance $6141 m0 *1 161.445,32.76
X$6141 524 24 525 644 645 cell_1rw
* cell instance $6142 m0 *1 162.15,32.76
X$6142 526 24 527 644 645 cell_1rw
* cell instance $6143 m0 *1 162.855,32.76
X$6143 528 24 529 644 645 cell_1rw
* cell instance $6144 m0 *1 163.56,32.76
X$6144 530 24 531 644 645 cell_1rw
* cell instance $6145 m0 *1 164.265,32.76
X$6145 532 24 533 644 645 cell_1rw
* cell instance $6146 m0 *1 164.97,32.76
X$6146 534 24 535 644 645 cell_1rw
* cell instance $6147 m0 *1 165.675,32.76
X$6147 536 24 537 644 645 cell_1rw
* cell instance $6148 m0 *1 166.38,32.76
X$6148 538 24 539 644 645 cell_1rw
* cell instance $6149 m0 *1 167.085,32.76
X$6149 540 24 541 644 645 cell_1rw
* cell instance $6150 m0 *1 167.79,32.76
X$6150 542 24 543 644 645 cell_1rw
* cell instance $6151 m0 *1 168.495,32.76
X$6151 544 24 545 644 645 cell_1rw
* cell instance $6152 m0 *1 169.2,32.76
X$6152 546 24 547 644 645 cell_1rw
* cell instance $6153 m0 *1 169.905,32.76
X$6153 548 24 549 644 645 cell_1rw
* cell instance $6154 m0 *1 170.61,32.76
X$6154 550 24 551 644 645 cell_1rw
* cell instance $6155 m0 *1 171.315,32.76
X$6155 552 24 553 644 645 cell_1rw
* cell instance $6156 m0 *1 172.02,32.76
X$6156 554 24 555 644 645 cell_1rw
* cell instance $6157 m0 *1 172.725,32.76
X$6157 556 24 557 644 645 cell_1rw
* cell instance $6158 m0 *1 173.43,32.76
X$6158 558 24 559 644 645 cell_1rw
* cell instance $6159 m0 *1 174.135,32.76
X$6159 560 24 561 644 645 cell_1rw
* cell instance $6160 m0 *1 174.84,32.76
X$6160 562 24 563 644 645 cell_1rw
* cell instance $6161 m0 *1 175.545,32.76
X$6161 564 24 565 644 645 cell_1rw
* cell instance $6162 m0 *1 176.25,32.76
X$6162 566 24 567 644 645 cell_1rw
* cell instance $6163 m0 *1 176.955,32.76
X$6163 568 24 569 644 645 cell_1rw
* cell instance $6164 m0 *1 177.66,32.76
X$6164 570 24 571 644 645 cell_1rw
* cell instance $6165 m0 *1 178.365,32.76
X$6165 572 24 573 644 645 cell_1rw
* cell instance $6166 m0 *1 179.07,32.76
X$6166 574 24 575 644 645 cell_1rw
* cell instance $6167 m0 *1 179.775,32.76
X$6167 576 24 577 644 645 cell_1rw
* cell instance $6168 m0 *1 180.48,32.76
X$6168 578 24 579 644 645 cell_1rw
* cell instance $6169 m0 *1 0.705,35.49
X$6169 67 25 68 644 645 cell_1rw
* cell instance $6170 m0 *1 0,35.49
X$6170 65 25 66 644 645 cell_1rw
* cell instance $6171 m0 *1 1.41,35.49
X$6171 69 25 70 644 645 cell_1rw
* cell instance $6172 m0 *1 2.115,35.49
X$6172 71 25 72 644 645 cell_1rw
* cell instance $6173 m0 *1 2.82,35.49
X$6173 73 25 74 644 645 cell_1rw
* cell instance $6174 m0 *1 3.525,35.49
X$6174 75 25 76 644 645 cell_1rw
* cell instance $6175 m0 *1 4.23,35.49
X$6175 77 25 78 644 645 cell_1rw
* cell instance $6176 m0 *1 4.935,35.49
X$6176 79 25 80 644 645 cell_1rw
* cell instance $6177 m0 *1 5.64,35.49
X$6177 81 25 82 644 645 cell_1rw
* cell instance $6178 m0 *1 6.345,35.49
X$6178 83 25 84 644 645 cell_1rw
* cell instance $6179 m0 *1 7.05,35.49
X$6179 85 25 86 644 645 cell_1rw
* cell instance $6180 m0 *1 7.755,35.49
X$6180 87 25 88 644 645 cell_1rw
* cell instance $6181 m0 *1 8.46,35.49
X$6181 89 25 90 644 645 cell_1rw
* cell instance $6182 m0 *1 9.165,35.49
X$6182 91 25 92 644 645 cell_1rw
* cell instance $6183 m0 *1 9.87,35.49
X$6183 93 25 94 644 645 cell_1rw
* cell instance $6184 m0 *1 10.575,35.49
X$6184 95 25 96 644 645 cell_1rw
* cell instance $6185 m0 *1 11.28,35.49
X$6185 97 25 98 644 645 cell_1rw
* cell instance $6186 m0 *1 11.985,35.49
X$6186 99 25 100 644 645 cell_1rw
* cell instance $6187 m0 *1 12.69,35.49
X$6187 101 25 102 644 645 cell_1rw
* cell instance $6188 m0 *1 13.395,35.49
X$6188 103 25 104 644 645 cell_1rw
* cell instance $6189 m0 *1 14.1,35.49
X$6189 105 25 106 644 645 cell_1rw
* cell instance $6190 m0 *1 14.805,35.49
X$6190 107 25 108 644 645 cell_1rw
* cell instance $6191 m0 *1 15.51,35.49
X$6191 109 25 110 644 645 cell_1rw
* cell instance $6192 m0 *1 16.215,35.49
X$6192 111 25 112 644 645 cell_1rw
* cell instance $6193 m0 *1 16.92,35.49
X$6193 113 25 114 644 645 cell_1rw
* cell instance $6194 m0 *1 17.625,35.49
X$6194 115 25 116 644 645 cell_1rw
* cell instance $6195 m0 *1 18.33,35.49
X$6195 117 25 118 644 645 cell_1rw
* cell instance $6196 m0 *1 19.035,35.49
X$6196 119 25 120 644 645 cell_1rw
* cell instance $6197 m0 *1 19.74,35.49
X$6197 121 25 122 644 645 cell_1rw
* cell instance $6198 m0 *1 20.445,35.49
X$6198 123 25 124 644 645 cell_1rw
* cell instance $6199 m0 *1 21.15,35.49
X$6199 125 25 126 644 645 cell_1rw
* cell instance $6200 m0 *1 21.855,35.49
X$6200 127 25 128 644 645 cell_1rw
* cell instance $6201 m0 *1 22.56,35.49
X$6201 129 25 130 644 645 cell_1rw
* cell instance $6202 m0 *1 23.265,35.49
X$6202 131 25 132 644 645 cell_1rw
* cell instance $6203 m0 *1 23.97,35.49
X$6203 133 25 134 644 645 cell_1rw
* cell instance $6204 m0 *1 24.675,35.49
X$6204 135 25 136 644 645 cell_1rw
* cell instance $6205 m0 *1 25.38,35.49
X$6205 137 25 138 644 645 cell_1rw
* cell instance $6206 m0 *1 26.085,35.49
X$6206 139 25 140 644 645 cell_1rw
* cell instance $6207 m0 *1 26.79,35.49
X$6207 141 25 142 644 645 cell_1rw
* cell instance $6208 m0 *1 27.495,35.49
X$6208 143 25 144 644 645 cell_1rw
* cell instance $6209 m0 *1 28.2,35.49
X$6209 145 25 146 644 645 cell_1rw
* cell instance $6210 m0 *1 28.905,35.49
X$6210 147 25 148 644 645 cell_1rw
* cell instance $6211 m0 *1 29.61,35.49
X$6211 149 25 150 644 645 cell_1rw
* cell instance $6212 m0 *1 30.315,35.49
X$6212 151 25 152 644 645 cell_1rw
* cell instance $6213 m0 *1 31.02,35.49
X$6213 153 25 154 644 645 cell_1rw
* cell instance $6214 m0 *1 31.725,35.49
X$6214 155 25 156 644 645 cell_1rw
* cell instance $6215 m0 *1 32.43,35.49
X$6215 157 25 158 644 645 cell_1rw
* cell instance $6216 m0 *1 33.135,35.49
X$6216 159 25 160 644 645 cell_1rw
* cell instance $6217 m0 *1 33.84,35.49
X$6217 161 25 162 644 645 cell_1rw
* cell instance $6218 m0 *1 34.545,35.49
X$6218 163 25 164 644 645 cell_1rw
* cell instance $6219 m0 *1 35.25,35.49
X$6219 165 25 166 644 645 cell_1rw
* cell instance $6220 m0 *1 35.955,35.49
X$6220 167 25 168 644 645 cell_1rw
* cell instance $6221 m0 *1 36.66,35.49
X$6221 169 25 170 644 645 cell_1rw
* cell instance $6222 m0 *1 37.365,35.49
X$6222 171 25 172 644 645 cell_1rw
* cell instance $6223 m0 *1 38.07,35.49
X$6223 173 25 174 644 645 cell_1rw
* cell instance $6224 m0 *1 38.775,35.49
X$6224 175 25 176 644 645 cell_1rw
* cell instance $6225 m0 *1 39.48,35.49
X$6225 177 25 178 644 645 cell_1rw
* cell instance $6226 m0 *1 40.185,35.49
X$6226 179 25 180 644 645 cell_1rw
* cell instance $6227 m0 *1 40.89,35.49
X$6227 181 25 182 644 645 cell_1rw
* cell instance $6228 m0 *1 41.595,35.49
X$6228 183 25 184 644 645 cell_1rw
* cell instance $6229 m0 *1 42.3,35.49
X$6229 185 25 186 644 645 cell_1rw
* cell instance $6230 m0 *1 43.005,35.49
X$6230 187 25 188 644 645 cell_1rw
* cell instance $6231 m0 *1 43.71,35.49
X$6231 189 25 190 644 645 cell_1rw
* cell instance $6232 m0 *1 44.415,35.49
X$6232 191 25 192 644 645 cell_1rw
* cell instance $6233 m0 *1 45.12,35.49
X$6233 193 25 194 644 645 cell_1rw
* cell instance $6234 m0 *1 45.825,35.49
X$6234 195 25 196 644 645 cell_1rw
* cell instance $6235 m0 *1 46.53,35.49
X$6235 197 25 198 644 645 cell_1rw
* cell instance $6236 m0 *1 47.235,35.49
X$6236 199 25 200 644 645 cell_1rw
* cell instance $6237 m0 *1 47.94,35.49
X$6237 201 25 202 644 645 cell_1rw
* cell instance $6238 m0 *1 48.645,35.49
X$6238 203 25 204 644 645 cell_1rw
* cell instance $6239 m0 *1 49.35,35.49
X$6239 205 25 206 644 645 cell_1rw
* cell instance $6240 m0 *1 50.055,35.49
X$6240 207 25 208 644 645 cell_1rw
* cell instance $6241 m0 *1 50.76,35.49
X$6241 209 25 210 644 645 cell_1rw
* cell instance $6242 m0 *1 51.465,35.49
X$6242 211 25 212 644 645 cell_1rw
* cell instance $6243 m0 *1 52.17,35.49
X$6243 213 25 214 644 645 cell_1rw
* cell instance $6244 m0 *1 52.875,35.49
X$6244 215 25 216 644 645 cell_1rw
* cell instance $6245 m0 *1 53.58,35.49
X$6245 217 25 218 644 645 cell_1rw
* cell instance $6246 m0 *1 54.285,35.49
X$6246 219 25 220 644 645 cell_1rw
* cell instance $6247 m0 *1 54.99,35.49
X$6247 221 25 222 644 645 cell_1rw
* cell instance $6248 m0 *1 55.695,35.49
X$6248 223 25 224 644 645 cell_1rw
* cell instance $6249 m0 *1 56.4,35.49
X$6249 225 25 226 644 645 cell_1rw
* cell instance $6250 m0 *1 57.105,35.49
X$6250 227 25 228 644 645 cell_1rw
* cell instance $6251 m0 *1 57.81,35.49
X$6251 229 25 230 644 645 cell_1rw
* cell instance $6252 m0 *1 58.515,35.49
X$6252 231 25 232 644 645 cell_1rw
* cell instance $6253 m0 *1 59.22,35.49
X$6253 233 25 234 644 645 cell_1rw
* cell instance $6254 m0 *1 59.925,35.49
X$6254 235 25 236 644 645 cell_1rw
* cell instance $6255 m0 *1 60.63,35.49
X$6255 237 25 238 644 645 cell_1rw
* cell instance $6256 m0 *1 61.335,35.49
X$6256 239 25 240 644 645 cell_1rw
* cell instance $6257 m0 *1 62.04,35.49
X$6257 241 25 242 644 645 cell_1rw
* cell instance $6258 m0 *1 62.745,35.49
X$6258 243 25 244 644 645 cell_1rw
* cell instance $6259 m0 *1 63.45,35.49
X$6259 245 25 246 644 645 cell_1rw
* cell instance $6260 m0 *1 64.155,35.49
X$6260 247 25 248 644 645 cell_1rw
* cell instance $6261 m0 *1 64.86,35.49
X$6261 249 25 250 644 645 cell_1rw
* cell instance $6262 m0 *1 65.565,35.49
X$6262 251 25 252 644 645 cell_1rw
* cell instance $6263 m0 *1 66.27,35.49
X$6263 253 25 254 644 645 cell_1rw
* cell instance $6264 m0 *1 66.975,35.49
X$6264 255 25 256 644 645 cell_1rw
* cell instance $6265 m0 *1 67.68,35.49
X$6265 257 25 258 644 645 cell_1rw
* cell instance $6266 m0 *1 68.385,35.49
X$6266 259 25 260 644 645 cell_1rw
* cell instance $6267 m0 *1 69.09,35.49
X$6267 261 25 262 644 645 cell_1rw
* cell instance $6268 m0 *1 69.795,35.49
X$6268 263 25 264 644 645 cell_1rw
* cell instance $6269 m0 *1 70.5,35.49
X$6269 265 25 266 644 645 cell_1rw
* cell instance $6270 m0 *1 71.205,35.49
X$6270 267 25 268 644 645 cell_1rw
* cell instance $6271 m0 *1 71.91,35.49
X$6271 269 25 270 644 645 cell_1rw
* cell instance $6272 m0 *1 72.615,35.49
X$6272 271 25 272 644 645 cell_1rw
* cell instance $6273 m0 *1 73.32,35.49
X$6273 273 25 274 644 645 cell_1rw
* cell instance $6274 m0 *1 74.025,35.49
X$6274 275 25 276 644 645 cell_1rw
* cell instance $6275 m0 *1 74.73,35.49
X$6275 277 25 278 644 645 cell_1rw
* cell instance $6276 m0 *1 75.435,35.49
X$6276 279 25 280 644 645 cell_1rw
* cell instance $6277 m0 *1 76.14,35.49
X$6277 281 25 282 644 645 cell_1rw
* cell instance $6278 m0 *1 76.845,35.49
X$6278 283 25 284 644 645 cell_1rw
* cell instance $6279 m0 *1 77.55,35.49
X$6279 285 25 286 644 645 cell_1rw
* cell instance $6280 m0 *1 78.255,35.49
X$6280 287 25 288 644 645 cell_1rw
* cell instance $6281 m0 *1 78.96,35.49
X$6281 289 25 290 644 645 cell_1rw
* cell instance $6282 m0 *1 79.665,35.49
X$6282 291 25 292 644 645 cell_1rw
* cell instance $6283 m0 *1 80.37,35.49
X$6283 293 25 294 644 645 cell_1rw
* cell instance $6284 m0 *1 81.075,35.49
X$6284 295 25 296 644 645 cell_1rw
* cell instance $6285 m0 *1 81.78,35.49
X$6285 297 25 298 644 645 cell_1rw
* cell instance $6286 m0 *1 82.485,35.49
X$6286 299 25 300 644 645 cell_1rw
* cell instance $6287 m0 *1 83.19,35.49
X$6287 301 25 302 644 645 cell_1rw
* cell instance $6288 m0 *1 83.895,35.49
X$6288 303 25 304 644 645 cell_1rw
* cell instance $6289 m0 *1 84.6,35.49
X$6289 305 25 306 644 645 cell_1rw
* cell instance $6290 m0 *1 85.305,35.49
X$6290 307 25 308 644 645 cell_1rw
* cell instance $6291 m0 *1 86.01,35.49
X$6291 309 25 310 644 645 cell_1rw
* cell instance $6292 m0 *1 86.715,35.49
X$6292 311 25 312 644 645 cell_1rw
* cell instance $6293 m0 *1 87.42,35.49
X$6293 313 25 314 644 645 cell_1rw
* cell instance $6294 m0 *1 88.125,35.49
X$6294 315 25 316 644 645 cell_1rw
* cell instance $6295 m0 *1 88.83,35.49
X$6295 317 25 318 644 645 cell_1rw
* cell instance $6296 m0 *1 89.535,35.49
X$6296 319 25 320 644 645 cell_1rw
* cell instance $6297 m0 *1 90.24,35.49
X$6297 321 25 323 644 645 cell_1rw
* cell instance $6298 m0 *1 90.945,35.49
X$6298 324 25 325 644 645 cell_1rw
* cell instance $6299 m0 *1 91.65,35.49
X$6299 326 25 327 644 645 cell_1rw
* cell instance $6300 m0 *1 92.355,35.49
X$6300 328 25 329 644 645 cell_1rw
* cell instance $6301 m0 *1 93.06,35.49
X$6301 330 25 331 644 645 cell_1rw
* cell instance $6302 m0 *1 93.765,35.49
X$6302 332 25 333 644 645 cell_1rw
* cell instance $6303 m0 *1 94.47,35.49
X$6303 334 25 335 644 645 cell_1rw
* cell instance $6304 m0 *1 95.175,35.49
X$6304 336 25 337 644 645 cell_1rw
* cell instance $6305 m0 *1 95.88,35.49
X$6305 338 25 339 644 645 cell_1rw
* cell instance $6306 m0 *1 96.585,35.49
X$6306 340 25 341 644 645 cell_1rw
* cell instance $6307 m0 *1 97.29,35.49
X$6307 342 25 343 644 645 cell_1rw
* cell instance $6308 m0 *1 97.995,35.49
X$6308 344 25 345 644 645 cell_1rw
* cell instance $6309 m0 *1 98.7,35.49
X$6309 346 25 347 644 645 cell_1rw
* cell instance $6310 m0 *1 99.405,35.49
X$6310 348 25 349 644 645 cell_1rw
* cell instance $6311 m0 *1 100.11,35.49
X$6311 350 25 351 644 645 cell_1rw
* cell instance $6312 m0 *1 100.815,35.49
X$6312 352 25 353 644 645 cell_1rw
* cell instance $6313 m0 *1 101.52,35.49
X$6313 354 25 355 644 645 cell_1rw
* cell instance $6314 m0 *1 102.225,35.49
X$6314 356 25 357 644 645 cell_1rw
* cell instance $6315 m0 *1 102.93,35.49
X$6315 358 25 359 644 645 cell_1rw
* cell instance $6316 m0 *1 103.635,35.49
X$6316 360 25 361 644 645 cell_1rw
* cell instance $6317 m0 *1 104.34,35.49
X$6317 362 25 363 644 645 cell_1rw
* cell instance $6318 m0 *1 105.045,35.49
X$6318 364 25 365 644 645 cell_1rw
* cell instance $6319 m0 *1 105.75,35.49
X$6319 366 25 367 644 645 cell_1rw
* cell instance $6320 m0 *1 106.455,35.49
X$6320 368 25 369 644 645 cell_1rw
* cell instance $6321 m0 *1 107.16,35.49
X$6321 370 25 371 644 645 cell_1rw
* cell instance $6322 m0 *1 107.865,35.49
X$6322 372 25 373 644 645 cell_1rw
* cell instance $6323 m0 *1 108.57,35.49
X$6323 374 25 375 644 645 cell_1rw
* cell instance $6324 m0 *1 109.275,35.49
X$6324 376 25 377 644 645 cell_1rw
* cell instance $6325 m0 *1 109.98,35.49
X$6325 378 25 379 644 645 cell_1rw
* cell instance $6326 m0 *1 110.685,35.49
X$6326 380 25 381 644 645 cell_1rw
* cell instance $6327 m0 *1 111.39,35.49
X$6327 382 25 383 644 645 cell_1rw
* cell instance $6328 m0 *1 112.095,35.49
X$6328 384 25 385 644 645 cell_1rw
* cell instance $6329 m0 *1 112.8,35.49
X$6329 386 25 387 644 645 cell_1rw
* cell instance $6330 m0 *1 113.505,35.49
X$6330 388 25 389 644 645 cell_1rw
* cell instance $6331 m0 *1 114.21,35.49
X$6331 390 25 391 644 645 cell_1rw
* cell instance $6332 m0 *1 114.915,35.49
X$6332 392 25 393 644 645 cell_1rw
* cell instance $6333 m0 *1 115.62,35.49
X$6333 394 25 395 644 645 cell_1rw
* cell instance $6334 m0 *1 116.325,35.49
X$6334 396 25 397 644 645 cell_1rw
* cell instance $6335 m0 *1 117.03,35.49
X$6335 398 25 399 644 645 cell_1rw
* cell instance $6336 m0 *1 117.735,35.49
X$6336 400 25 401 644 645 cell_1rw
* cell instance $6337 m0 *1 118.44,35.49
X$6337 402 25 403 644 645 cell_1rw
* cell instance $6338 m0 *1 119.145,35.49
X$6338 404 25 405 644 645 cell_1rw
* cell instance $6339 m0 *1 119.85,35.49
X$6339 406 25 407 644 645 cell_1rw
* cell instance $6340 m0 *1 120.555,35.49
X$6340 408 25 409 644 645 cell_1rw
* cell instance $6341 m0 *1 121.26,35.49
X$6341 410 25 411 644 645 cell_1rw
* cell instance $6342 m0 *1 121.965,35.49
X$6342 412 25 413 644 645 cell_1rw
* cell instance $6343 m0 *1 122.67,35.49
X$6343 414 25 415 644 645 cell_1rw
* cell instance $6344 m0 *1 123.375,35.49
X$6344 416 25 417 644 645 cell_1rw
* cell instance $6345 m0 *1 124.08,35.49
X$6345 418 25 419 644 645 cell_1rw
* cell instance $6346 m0 *1 124.785,35.49
X$6346 420 25 421 644 645 cell_1rw
* cell instance $6347 m0 *1 125.49,35.49
X$6347 422 25 423 644 645 cell_1rw
* cell instance $6348 m0 *1 126.195,35.49
X$6348 424 25 425 644 645 cell_1rw
* cell instance $6349 m0 *1 126.9,35.49
X$6349 426 25 427 644 645 cell_1rw
* cell instance $6350 m0 *1 127.605,35.49
X$6350 428 25 429 644 645 cell_1rw
* cell instance $6351 m0 *1 128.31,35.49
X$6351 430 25 431 644 645 cell_1rw
* cell instance $6352 m0 *1 129.015,35.49
X$6352 432 25 433 644 645 cell_1rw
* cell instance $6353 m0 *1 129.72,35.49
X$6353 434 25 435 644 645 cell_1rw
* cell instance $6354 m0 *1 130.425,35.49
X$6354 436 25 437 644 645 cell_1rw
* cell instance $6355 m0 *1 131.13,35.49
X$6355 438 25 439 644 645 cell_1rw
* cell instance $6356 m0 *1 131.835,35.49
X$6356 440 25 441 644 645 cell_1rw
* cell instance $6357 m0 *1 132.54,35.49
X$6357 442 25 443 644 645 cell_1rw
* cell instance $6358 m0 *1 133.245,35.49
X$6358 444 25 445 644 645 cell_1rw
* cell instance $6359 m0 *1 133.95,35.49
X$6359 446 25 447 644 645 cell_1rw
* cell instance $6360 m0 *1 134.655,35.49
X$6360 448 25 449 644 645 cell_1rw
* cell instance $6361 m0 *1 135.36,35.49
X$6361 450 25 451 644 645 cell_1rw
* cell instance $6362 m0 *1 136.065,35.49
X$6362 452 25 453 644 645 cell_1rw
* cell instance $6363 m0 *1 136.77,35.49
X$6363 454 25 455 644 645 cell_1rw
* cell instance $6364 m0 *1 137.475,35.49
X$6364 456 25 457 644 645 cell_1rw
* cell instance $6365 m0 *1 138.18,35.49
X$6365 458 25 459 644 645 cell_1rw
* cell instance $6366 m0 *1 138.885,35.49
X$6366 460 25 461 644 645 cell_1rw
* cell instance $6367 m0 *1 139.59,35.49
X$6367 462 25 463 644 645 cell_1rw
* cell instance $6368 m0 *1 140.295,35.49
X$6368 464 25 465 644 645 cell_1rw
* cell instance $6369 m0 *1 141,35.49
X$6369 466 25 467 644 645 cell_1rw
* cell instance $6370 m0 *1 141.705,35.49
X$6370 468 25 469 644 645 cell_1rw
* cell instance $6371 m0 *1 142.41,35.49
X$6371 470 25 471 644 645 cell_1rw
* cell instance $6372 m0 *1 143.115,35.49
X$6372 472 25 473 644 645 cell_1rw
* cell instance $6373 m0 *1 143.82,35.49
X$6373 474 25 475 644 645 cell_1rw
* cell instance $6374 m0 *1 144.525,35.49
X$6374 476 25 477 644 645 cell_1rw
* cell instance $6375 m0 *1 145.23,35.49
X$6375 478 25 479 644 645 cell_1rw
* cell instance $6376 m0 *1 145.935,35.49
X$6376 480 25 481 644 645 cell_1rw
* cell instance $6377 m0 *1 146.64,35.49
X$6377 482 25 483 644 645 cell_1rw
* cell instance $6378 m0 *1 147.345,35.49
X$6378 484 25 485 644 645 cell_1rw
* cell instance $6379 m0 *1 148.05,35.49
X$6379 486 25 487 644 645 cell_1rw
* cell instance $6380 m0 *1 148.755,35.49
X$6380 488 25 489 644 645 cell_1rw
* cell instance $6381 m0 *1 149.46,35.49
X$6381 490 25 491 644 645 cell_1rw
* cell instance $6382 m0 *1 150.165,35.49
X$6382 492 25 493 644 645 cell_1rw
* cell instance $6383 m0 *1 150.87,35.49
X$6383 494 25 495 644 645 cell_1rw
* cell instance $6384 m0 *1 151.575,35.49
X$6384 496 25 497 644 645 cell_1rw
* cell instance $6385 m0 *1 152.28,35.49
X$6385 498 25 499 644 645 cell_1rw
* cell instance $6386 m0 *1 152.985,35.49
X$6386 500 25 501 644 645 cell_1rw
* cell instance $6387 m0 *1 153.69,35.49
X$6387 502 25 503 644 645 cell_1rw
* cell instance $6388 m0 *1 154.395,35.49
X$6388 504 25 505 644 645 cell_1rw
* cell instance $6389 m0 *1 155.1,35.49
X$6389 506 25 507 644 645 cell_1rw
* cell instance $6390 m0 *1 155.805,35.49
X$6390 508 25 509 644 645 cell_1rw
* cell instance $6391 m0 *1 156.51,35.49
X$6391 510 25 511 644 645 cell_1rw
* cell instance $6392 m0 *1 157.215,35.49
X$6392 512 25 513 644 645 cell_1rw
* cell instance $6393 m0 *1 157.92,35.49
X$6393 514 25 515 644 645 cell_1rw
* cell instance $6394 m0 *1 158.625,35.49
X$6394 516 25 517 644 645 cell_1rw
* cell instance $6395 m0 *1 159.33,35.49
X$6395 518 25 519 644 645 cell_1rw
* cell instance $6396 m0 *1 160.035,35.49
X$6396 520 25 521 644 645 cell_1rw
* cell instance $6397 m0 *1 160.74,35.49
X$6397 522 25 523 644 645 cell_1rw
* cell instance $6398 m0 *1 161.445,35.49
X$6398 524 25 525 644 645 cell_1rw
* cell instance $6399 m0 *1 162.15,35.49
X$6399 526 25 527 644 645 cell_1rw
* cell instance $6400 m0 *1 162.855,35.49
X$6400 528 25 529 644 645 cell_1rw
* cell instance $6401 m0 *1 163.56,35.49
X$6401 530 25 531 644 645 cell_1rw
* cell instance $6402 m0 *1 164.265,35.49
X$6402 532 25 533 644 645 cell_1rw
* cell instance $6403 m0 *1 164.97,35.49
X$6403 534 25 535 644 645 cell_1rw
* cell instance $6404 m0 *1 165.675,35.49
X$6404 536 25 537 644 645 cell_1rw
* cell instance $6405 m0 *1 166.38,35.49
X$6405 538 25 539 644 645 cell_1rw
* cell instance $6406 m0 *1 167.085,35.49
X$6406 540 25 541 644 645 cell_1rw
* cell instance $6407 m0 *1 167.79,35.49
X$6407 542 25 543 644 645 cell_1rw
* cell instance $6408 m0 *1 168.495,35.49
X$6408 544 25 545 644 645 cell_1rw
* cell instance $6409 m0 *1 169.2,35.49
X$6409 546 25 547 644 645 cell_1rw
* cell instance $6410 m0 *1 169.905,35.49
X$6410 548 25 549 644 645 cell_1rw
* cell instance $6411 m0 *1 170.61,35.49
X$6411 550 25 551 644 645 cell_1rw
* cell instance $6412 m0 *1 171.315,35.49
X$6412 552 25 553 644 645 cell_1rw
* cell instance $6413 m0 *1 172.02,35.49
X$6413 554 25 555 644 645 cell_1rw
* cell instance $6414 m0 *1 172.725,35.49
X$6414 556 25 557 644 645 cell_1rw
* cell instance $6415 m0 *1 173.43,35.49
X$6415 558 25 559 644 645 cell_1rw
* cell instance $6416 m0 *1 174.135,35.49
X$6416 560 25 561 644 645 cell_1rw
* cell instance $6417 m0 *1 174.84,35.49
X$6417 562 25 563 644 645 cell_1rw
* cell instance $6418 m0 *1 175.545,35.49
X$6418 564 25 565 644 645 cell_1rw
* cell instance $6419 m0 *1 176.25,35.49
X$6419 566 25 567 644 645 cell_1rw
* cell instance $6420 m0 *1 176.955,35.49
X$6420 568 25 569 644 645 cell_1rw
* cell instance $6421 m0 *1 177.66,35.49
X$6421 570 25 571 644 645 cell_1rw
* cell instance $6422 m0 *1 178.365,35.49
X$6422 572 25 573 644 645 cell_1rw
* cell instance $6423 m0 *1 179.07,35.49
X$6423 574 25 575 644 645 cell_1rw
* cell instance $6424 m0 *1 179.775,35.49
X$6424 576 25 577 644 645 cell_1rw
* cell instance $6425 m0 *1 180.48,35.49
X$6425 578 25 579 644 645 cell_1rw
* cell instance $6426 r0 *1 0.705,32.76
X$6426 67 26 68 644 645 cell_1rw
* cell instance $6427 r0 *1 0,32.76
X$6427 65 26 66 644 645 cell_1rw
* cell instance $6428 r0 *1 1.41,32.76
X$6428 69 26 70 644 645 cell_1rw
* cell instance $6429 r0 *1 2.115,32.76
X$6429 71 26 72 644 645 cell_1rw
* cell instance $6430 r0 *1 2.82,32.76
X$6430 73 26 74 644 645 cell_1rw
* cell instance $6431 r0 *1 3.525,32.76
X$6431 75 26 76 644 645 cell_1rw
* cell instance $6432 r0 *1 4.23,32.76
X$6432 77 26 78 644 645 cell_1rw
* cell instance $6433 r0 *1 4.935,32.76
X$6433 79 26 80 644 645 cell_1rw
* cell instance $6434 r0 *1 5.64,32.76
X$6434 81 26 82 644 645 cell_1rw
* cell instance $6435 r0 *1 6.345,32.76
X$6435 83 26 84 644 645 cell_1rw
* cell instance $6436 r0 *1 7.05,32.76
X$6436 85 26 86 644 645 cell_1rw
* cell instance $6437 r0 *1 7.755,32.76
X$6437 87 26 88 644 645 cell_1rw
* cell instance $6438 r0 *1 8.46,32.76
X$6438 89 26 90 644 645 cell_1rw
* cell instance $6439 r0 *1 9.165,32.76
X$6439 91 26 92 644 645 cell_1rw
* cell instance $6440 r0 *1 9.87,32.76
X$6440 93 26 94 644 645 cell_1rw
* cell instance $6441 r0 *1 10.575,32.76
X$6441 95 26 96 644 645 cell_1rw
* cell instance $6442 r0 *1 11.28,32.76
X$6442 97 26 98 644 645 cell_1rw
* cell instance $6443 r0 *1 11.985,32.76
X$6443 99 26 100 644 645 cell_1rw
* cell instance $6444 r0 *1 12.69,32.76
X$6444 101 26 102 644 645 cell_1rw
* cell instance $6445 r0 *1 13.395,32.76
X$6445 103 26 104 644 645 cell_1rw
* cell instance $6446 r0 *1 14.1,32.76
X$6446 105 26 106 644 645 cell_1rw
* cell instance $6447 r0 *1 14.805,32.76
X$6447 107 26 108 644 645 cell_1rw
* cell instance $6448 r0 *1 15.51,32.76
X$6448 109 26 110 644 645 cell_1rw
* cell instance $6449 r0 *1 16.215,32.76
X$6449 111 26 112 644 645 cell_1rw
* cell instance $6450 r0 *1 16.92,32.76
X$6450 113 26 114 644 645 cell_1rw
* cell instance $6451 r0 *1 17.625,32.76
X$6451 115 26 116 644 645 cell_1rw
* cell instance $6452 r0 *1 18.33,32.76
X$6452 117 26 118 644 645 cell_1rw
* cell instance $6453 r0 *1 19.035,32.76
X$6453 119 26 120 644 645 cell_1rw
* cell instance $6454 r0 *1 19.74,32.76
X$6454 121 26 122 644 645 cell_1rw
* cell instance $6455 r0 *1 20.445,32.76
X$6455 123 26 124 644 645 cell_1rw
* cell instance $6456 r0 *1 21.15,32.76
X$6456 125 26 126 644 645 cell_1rw
* cell instance $6457 r0 *1 21.855,32.76
X$6457 127 26 128 644 645 cell_1rw
* cell instance $6458 r0 *1 22.56,32.76
X$6458 129 26 130 644 645 cell_1rw
* cell instance $6459 r0 *1 23.265,32.76
X$6459 131 26 132 644 645 cell_1rw
* cell instance $6460 r0 *1 23.97,32.76
X$6460 133 26 134 644 645 cell_1rw
* cell instance $6461 r0 *1 24.675,32.76
X$6461 135 26 136 644 645 cell_1rw
* cell instance $6462 r0 *1 25.38,32.76
X$6462 137 26 138 644 645 cell_1rw
* cell instance $6463 r0 *1 26.085,32.76
X$6463 139 26 140 644 645 cell_1rw
* cell instance $6464 r0 *1 26.79,32.76
X$6464 141 26 142 644 645 cell_1rw
* cell instance $6465 r0 *1 27.495,32.76
X$6465 143 26 144 644 645 cell_1rw
* cell instance $6466 r0 *1 28.2,32.76
X$6466 145 26 146 644 645 cell_1rw
* cell instance $6467 r0 *1 28.905,32.76
X$6467 147 26 148 644 645 cell_1rw
* cell instance $6468 r0 *1 29.61,32.76
X$6468 149 26 150 644 645 cell_1rw
* cell instance $6469 r0 *1 30.315,32.76
X$6469 151 26 152 644 645 cell_1rw
* cell instance $6470 r0 *1 31.02,32.76
X$6470 153 26 154 644 645 cell_1rw
* cell instance $6471 r0 *1 31.725,32.76
X$6471 155 26 156 644 645 cell_1rw
* cell instance $6472 r0 *1 32.43,32.76
X$6472 157 26 158 644 645 cell_1rw
* cell instance $6473 r0 *1 33.135,32.76
X$6473 159 26 160 644 645 cell_1rw
* cell instance $6474 r0 *1 33.84,32.76
X$6474 161 26 162 644 645 cell_1rw
* cell instance $6475 r0 *1 34.545,32.76
X$6475 163 26 164 644 645 cell_1rw
* cell instance $6476 r0 *1 35.25,32.76
X$6476 165 26 166 644 645 cell_1rw
* cell instance $6477 r0 *1 35.955,32.76
X$6477 167 26 168 644 645 cell_1rw
* cell instance $6478 r0 *1 36.66,32.76
X$6478 169 26 170 644 645 cell_1rw
* cell instance $6479 r0 *1 37.365,32.76
X$6479 171 26 172 644 645 cell_1rw
* cell instance $6480 r0 *1 38.07,32.76
X$6480 173 26 174 644 645 cell_1rw
* cell instance $6481 r0 *1 38.775,32.76
X$6481 175 26 176 644 645 cell_1rw
* cell instance $6482 r0 *1 39.48,32.76
X$6482 177 26 178 644 645 cell_1rw
* cell instance $6483 r0 *1 40.185,32.76
X$6483 179 26 180 644 645 cell_1rw
* cell instance $6484 r0 *1 40.89,32.76
X$6484 181 26 182 644 645 cell_1rw
* cell instance $6485 r0 *1 41.595,32.76
X$6485 183 26 184 644 645 cell_1rw
* cell instance $6486 r0 *1 42.3,32.76
X$6486 185 26 186 644 645 cell_1rw
* cell instance $6487 r0 *1 43.005,32.76
X$6487 187 26 188 644 645 cell_1rw
* cell instance $6488 r0 *1 43.71,32.76
X$6488 189 26 190 644 645 cell_1rw
* cell instance $6489 r0 *1 44.415,32.76
X$6489 191 26 192 644 645 cell_1rw
* cell instance $6490 r0 *1 45.12,32.76
X$6490 193 26 194 644 645 cell_1rw
* cell instance $6491 r0 *1 45.825,32.76
X$6491 195 26 196 644 645 cell_1rw
* cell instance $6492 r0 *1 46.53,32.76
X$6492 197 26 198 644 645 cell_1rw
* cell instance $6493 r0 *1 47.235,32.76
X$6493 199 26 200 644 645 cell_1rw
* cell instance $6494 r0 *1 47.94,32.76
X$6494 201 26 202 644 645 cell_1rw
* cell instance $6495 r0 *1 48.645,32.76
X$6495 203 26 204 644 645 cell_1rw
* cell instance $6496 r0 *1 49.35,32.76
X$6496 205 26 206 644 645 cell_1rw
* cell instance $6497 r0 *1 50.055,32.76
X$6497 207 26 208 644 645 cell_1rw
* cell instance $6498 r0 *1 50.76,32.76
X$6498 209 26 210 644 645 cell_1rw
* cell instance $6499 r0 *1 51.465,32.76
X$6499 211 26 212 644 645 cell_1rw
* cell instance $6500 r0 *1 52.17,32.76
X$6500 213 26 214 644 645 cell_1rw
* cell instance $6501 r0 *1 52.875,32.76
X$6501 215 26 216 644 645 cell_1rw
* cell instance $6502 r0 *1 53.58,32.76
X$6502 217 26 218 644 645 cell_1rw
* cell instance $6503 r0 *1 54.285,32.76
X$6503 219 26 220 644 645 cell_1rw
* cell instance $6504 r0 *1 54.99,32.76
X$6504 221 26 222 644 645 cell_1rw
* cell instance $6505 r0 *1 55.695,32.76
X$6505 223 26 224 644 645 cell_1rw
* cell instance $6506 r0 *1 56.4,32.76
X$6506 225 26 226 644 645 cell_1rw
* cell instance $6507 r0 *1 57.105,32.76
X$6507 227 26 228 644 645 cell_1rw
* cell instance $6508 r0 *1 57.81,32.76
X$6508 229 26 230 644 645 cell_1rw
* cell instance $6509 r0 *1 58.515,32.76
X$6509 231 26 232 644 645 cell_1rw
* cell instance $6510 r0 *1 59.22,32.76
X$6510 233 26 234 644 645 cell_1rw
* cell instance $6511 r0 *1 59.925,32.76
X$6511 235 26 236 644 645 cell_1rw
* cell instance $6512 r0 *1 60.63,32.76
X$6512 237 26 238 644 645 cell_1rw
* cell instance $6513 r0 *1 61.335,32.76
X$6513 239 26 240 644 645 cell_1rw
* cell instance $6514 r0 *1 62.04,32.76
X$6514 241 26 242 644 645 cell_1rw
* cell instance $6515 r0 *1 62.745,32.76
X$6515 243 26 244 644 645 cell_1rw
* cell instance $6516 r0 *1 63.45,32.76
X$6516 245 26 246 644 645 cell_1rw
* cell instance $6517 r0 *1 64.155,32.76
X$6517 247 26 248 644 645 cell_1rw
* cell instance $6518 r0 *1 64.86,32.76
X$6518 249 26 250 644 645 cell_1rw
* cell instance $6519 r0 *1 65.565,32.76
X$6519 251 26 252 644 645 cell_1rw
* cell instance $6520 r0 *1 66.27,32.76
X$6520 253 26 254 644 645 cell_1rw
* cell instance $6521 r0 *1 66.975,32.76
X$6521 255 26 256 644 645 cell_1rw
* cell instance $6522 r0 *1 67.68,32.76
X$6522 257 26 258 644 645 cell_1rw
* cell instance $6523 r0 *1 68.385,32.76
X$6523 259 26 260 644 645 cell_1rw
* cell instance $6524 r0 *1 69.09,32.76
X$6524 261 26 262 644 645 cell_1rw
* cell instance $6525 r0 *1 69.795,32.76
X$6525 263 26 264 644 645 cell_1rw
* cell instance $6526 r0 *1 70.5,32.76
X$6526 265 26 266 644 645 cell_1rw
* cell instance $6527 r0 *1 71.205,32.76
X$6527 267 26 268 644 645 cell_1rw
* cell instance $6528 r0 *1 71.91,32.76
X$6528 269 26 270 644 645 cell_1rw
* cell instance $6529 r0 *1 72.615,32.76
X$6529 271 26 272 644 645 cell_1rw
* cell instance $6530 r0 *1 73.32,32.76
X$6530 273 26 274 644 645 cell_1rw
* cell instance $6531 r0 *1 74.025,32.76
X$6531 275 26 276 644 645 cell_1rw
* cell instance $6532 r0 *1 74.73,32.76
X$6532 277 26 278 644 645 cell_1rw
* cell instance $6533 r0 *1 75.435,32.76
X$6533 279 26 280 644 645 cell_1rw
* cell instance $6534 r0 *1 76.14,32.76
X$6534 281 26 282 644 645 cell_1rw
* cell instance $6535 r0 *1 76.845,32.76
X$6535 283 26 284 644 645 cell_1rw
* cell instance $6536 r0 *1 77.55,32.76
X$6536 285 26 286 644 645 cell_1rw
* cell instance $6537 r0 *1 78.255,32.76
X$6537 287 26 288 644 645 cell_1rw
* cell instance $6538 r0 *1 78.96,32.76
X$6538 289 26 290 644 645 cell_1rw
* cell instance $6539 r0 *1 79.665,32.76
X$6539 291 26 292 644 645 cell_1rw
* cell instance $6540 r0 *1 80.37,32.76
X$6540 293 26 294 644 645 cell_1rw
* cell instance $6541 r0 *1 81.075,32.76
X$6541 295 26 296 644 645 cell_1rw
* cell instance $6542 r0 *1 81.78,32.76
X$6542 297 26 298 644 645 cell_1rw
* cell instance $6543 r0 *1 82.485,32.76
X$6543 299 26 300 644 645 cell_1rw
* cell instance $6544 r0 *1 83.19,32.76
X$6544 301 26 302 644 645 cell_1rw
* cell instance $6545 r0 *1 83.895,32.76
X$6545 303 26 304 644 645 cell_1rw
* cell instance $6546 r0 *1 84.6,32.76
X$6546 305 26 306 644 645 cell_1rw
* cell instance $6547 r0 *1 85.305,32.76
X$6547 307 26 308 644 645 cell_1rw
* cell instance $6548 r0 *1 86.01,32.76
X$6548 309 26 310 644 645 cell_1rw
* cell instance $6549 r0 *1 86.715,32.76
X$6549 311 26 312 644 645 cell_1rw
* cell instance $6550 r0 *1 87.42,32.76
X$6550 313 26 314 644 645 cell_1rw
* cell instance $6551 r0 *1 88.125,32.76
X$6551 315 26 316 644 645 cell_1rw
* cell instance $6552 r0 *1 88.83,32.76
X$6552 317 26 318 644 645 cell_1rw
* cell instance $6553 r0 *1 89.535,32.76
X$6553 319 26 320 644 645 cell_1rw
* cell instance $6554 r0 *1 90.24,32.76
X$6554 321 26 323 644 645 cell_1rw
* cell instance $6555 r0 *1 90.945,32.76
X$6555 324 26 325 644 645 cell_1rw
* cell instance $6556 r0 *1 91.65,32.76
X$6556 326 26 327 644 645 cell_1rw
* cell instance $6557 r0 *1 92.355,32.76
X$6557 328 26 329 644 645 cell_1rw
* cell instance $6558 r0 *1 93.06,32.76
X$6558 330 26 331 644 645 cell_1rw
* cell instance $6559 r0 *1 93.765,32.76
X$6559 332 26 333 644 645 cell_1rw
* cell instance $6560 r0 *1 94.47,32.76
X$6560 334 26 335 644 645 cell_1rw
* cell instance $6561 r0 *1 95.175,32.76
X$6561 336 26 337 644 645 cell_1rw
* cell instance $6562 r0 *1 95.88,32.76
X$6562 338 26 339 644 645 cell_1rw
* cell instance $6563 r0 *1 96.585,32.76
X$6563 340 26 341 644 645 cell_1rw
* cell instance $6564 r0 *1 97.29,32.76
X$6564 342 26 343 644 645 cell_1rw
* cell instance $6565 r0 *1 97.995,32.76
X$6565 344 26 345 644 645 cell_1rw
* cell instance $6566 r0 *1 98.7,32.76
X$6566 346 26 347 644 645 cell_1rw
* cell instance $6567 r0 *1 99.405,32.76
X$6567 348 26 349 644 645 cell_1rw
* cell instance $6568 r0 *1 100.11,32.76
X$6568 350 26 351 644 645 cell_1rw
* cell instance $6569 r0 *1 100.815,32.76
X$6569 352 26 353 644 645 cell_1rw
* cell instance $6570 r0 *1 101.52,32.76
X$6570 354 26 355 644 645 cell_1rw
* cell instance $6571 r0 *1 102.225,32.76
X$6571 356 26 357 644 645 cell_1rw
* cell instance $6572 r0 *1 102.93,32.76
X$6572 358 26 359 644 645 cell_1rw
* cell instance $6573 r0 *1 103.635,32.76
X$6573 360 26 361 644 645 cell_1rw
* cell instance $6574 r0 *1 104.34,32.76
X$6574 362 26 363 644 645 cell_1rw
* cell instance $6575 r0 *1 105.045,32.76
X$6575 364 26 365 644 645 cell_1rw
* cell instance $6576 r0 *1 105.75,32.76
X$6576 366 26 367 644 645 cell_1rw
* cell instance $6577 r0 *1 106.455,32.76
X$6577 368 26 369 644 645 cell_1rw
* cell instance $6578 r0 *1 107.16,32.76
X$6578 370 26 371 644 645 cell_1rw
* cell instance $6579 r0 *1 107.865,32.76
X$6579 372 26 373 644 645 cell_1rw
* cell instance $6580 r0 *1 108.57,32.76
X$6580 374 26 375 644 645 cell_1rw
* cell instance $6581 r0 *1 109.275,32.76
X$6581 376 26 377 644 645 cell_1rw
* cell instance $6582 r0 *1 109.98,32.76
X$6582 378 26 379 644 645 cell_1rw
* cell instance $6583 r0 *1 110.685,32.76
X$6583 380 26 381 644 645 cell_1rw
* cell instance $6584 r0 *1 111.39,32.76
X$6584 382 26 383 644 645 cell_1rw
* cell instance $6585 r0 *1 112.095,32.76
X$6585 384 26 385 644 645 cell_1rw
* cell instance $6586 r0 *1 112.8,32.76
X$6586 386 26 387 644 645 cell_1rw
* cell instance $6587 r0 *1 113.505,32.76
X$6587 388 26 389 644 645 cell_1rw
* cell instance $6588 r0 *1 114.21,32.76
X$6588 390 26 391 644 645 cell_1rw
* cell instance $6589 r0 *1 114.915,32.76
X$6589 392 26 393 644 645 cell_1rw
* cell instance $6590 r0 *1 115.62,32.76
X$6590 394 26 395 644 645 cell_1rw
* cell instance $6591 r0 *1 116.325,32.76
X$6591 396 26 397 644 645 cell_1rw
* cell instance $6592 r0 *1 117.03,32.76
X$6592 398 26 399 644 645 cell_1rw
* cell instance $6593 r0 *1 117.735,32.76
X$6593 400 26 401 644 645 cell_1rw
* cell instance $6594 r0 *1 118.44,32.76
X$6594 402 26 403 644 645 cell_1rw
* cell instance $6595 r0 *1 119.145,32.76
X$6595 404 26 405 644 645 cell_1rw
* cell instance $6596 r0 *1 119.85,32.76
X$6596 406 26 407 644 645 cell_1rw
* cell instance $6597 r0 *1 120.555,32.76
X$6597 408 26 409 644 645 cell_1rw
* cell instance $6598 r0 *1 121.26,32.76
X$6598 410 26 411 644 645 cell_1rw
* cell instance $6599 r0 *1 121.965,32.76
X$6599 412 26 413 644 645 cell_1rw
* cell instance $6600 r0 *1 122.67,32.76
X$6600 414 26 415 644 645 cell_1rw
* cell instance $6601 r0 *1 123.375,32.76
X$6601 416 26 417 644 645 cell_1rw
* cell instance $6602 r0 *1 124.08,32.76
X$6602 418 26 419 644 645 cell_1rw
* cell instance $6603 r0 *1 124.785,32.76
X$6603 420 26 421 644 645 cell_1rw
* cell instance $6604 r0 *1 125.49,32.76
X$6604 422 26 423 644 645 cell_1rw
* cell instance $6605 r0 *1 126.195,32.76
X$6605 424 26 425 644 645 cell_1rw
* cell instance $6606 r0 *1 126.9,32.76
X$6606 426 26 427 644 645 cell_1rw
* cell instance $6607 r0 *1 127.605,32.76
X$6607 428 26 429 644 645 cell_1rw
* cell instance $6608 r0 *1 128.31,32.76
X$6608 430 26 431 644 645 cell_1rw
* cell instance $6609 r0 *1 129.015,32.76
X$6609 432 26 433 644 645 cell_1rw
* cell instance $6610 r0 *1 129.72,32.76
X$6610 434 26 435 644 645 cell_1rw
* cell instance $6611 r0 *1 130.425,32.76
X$6611 436 26 437 644 645 cell_1rw
* cell instance $6612 r0 *1 131.13,32.76
X$6612 438 26 439 644 645 cell_1rw
* cell instance $6613 r0 *1 131.835,32.76
X$6613 440 26 441 644 645 cell_1rw
* cell instance $6614 r0 *1 132.54,32.76
X$6614 442 26 443 644 645 cell_1rw
* cell instance $6615 r0 *1 133.245,32.76
X$6615 444 26 445 644 645 cell_1rw
* cell instance $6616 r0 *1 133.95,32.76
X$6616 446 26 447 644 645 cell_1rw
* cell instance $6617 r0 *1 134.655,32.76
X$6617 448 26 449 644 645 cell_1rw
* cell instance $6618 r0 *1 135.36,32.76
X$6618 450 26 451 644 645 cell_1rw
* cell instance $6619 r0 *1 136.065,32.76
X$6619 452 26 453 644 645 cell_1rw
* cell instance $6620 r0 *1 136.77,32.76
X$6620 454 26 455 644 645 cell_1rw
* cell instance $6621 r0 *1 137.475,32.76
X$6621 456 26 457 644 645 cell_1rw
* cell instance $6622 r0 *1 138.18,32.76
X$6622 458 26 459 644 645 cell_1rw
* cell instance $6623 r0 *1 138.885,32.76
X$6623 460 26 461 644 645 cell_1rw
* cell instance $6624 r0 *1 139.59,32.76
X$6624 462 26 463 644 645 cell_1rw
* cell instance $6625 r0 *1 140.295,32.76
X$6625 464 26 465 644 645 cell_1rw
* cell instance $6626 r0 *1 141,32.76
X$6626 466 26 467 644 645 cell_1rw
* cell instance $6627 r0 *1 141.705,32.76
X$6627 468 26 469 644 645 cell_1rw
* cell instance $6628 r0 *1 142.41,32.76
X$6628 470 26 471 644 645 cell_1rw
* cell instance $6629 r0 *1 143.115,32.76
X$6629 472 26 473 644 645 cell_1rw
* cell instance $6630 r0 *1 143.82,32.76
X$6630 474 26 475 644 645 cell_1rw
* cell instance $6631 r0 *1 144.525,32.76
X$6631 476 26 477 644 645 cell_1rw
* cell instance $6632 r0 *1 145.23,32.76
X$6632 478 26 479 644 645 cell_1rw
* cell instance $6633 r0 *1 145.935,32.76
X$6633 480 26 481 644 645 cell_1rw
* cell instance $6634 r0 *1 146.64,32.76
X$6634 482 26 483 644 645 cell_1rw
* cell instance $6635 r0 *1 147.345,32.76
X$6635 484 26 485 644 645 cell_1rw
* cell instance $6636 r0 *1 148.05,32.76
X$6636 486 26 487 644 645 cell_1rw
* cell instance $6637 r0 *1 148.755,32.76
X$6637 488 26 489 644 645 cell_1rw
* cell instance $6638 r0 *1 149.46,32.76
X$6638 490 26 491 644 645 cell_1rw
* cell instance $6639 r0 *1 150.165,32.76
X$6639 492 26 493 644 645 cell_1rw
* cell instance $6640 r0 *1 150.87,32.76
X$6640 494 26 495 644 645 cell_1rw
* cell instance $6641 r0 *1 151.575,32.76
X$6641 496 26 497 644 645 cell_1rw
* cell instance $6642 r0 *1 152.28,32.76
X$6642 498 26 499 644 645 cell_1rw
* cell instance $6643 r0 *1 152.985,32.76
X$6643 500 26 501 644 645 cell_1rw
* cell instance $6644 r0 *1 153.69,32.76
X$6644 502 26 503 644 645 cell_1rw
* cell instance $6645 r0 *1 154.395,32.76
X$6645 504 26 505 644 645 cell_1rw
* cell instance $6646 r0 *1 155.1,32.76
X$6646 506 26 507 644 645 cell_1rw
* cell instance $6647 r0 *1 155.805,32.76
X$6647 508 26 509 644 645 cell_1rw
* cell instance $6648 r0 *1 156.51,32.76
X$6648 510 26 511 644 645 cell_1rw
* cell instance $6649 r0 *1 157.215,32.76
X$6649 512 26 513 644 645 cell_1rw
* cell instance $6650 r0 *1 157.92,32.76
X$6650 514 26 515 644 645 cell_1rw
* cell instance $6651 r0 *1 158.625,32.76
X$6651 516 26 517 644 645 cell_1rw
* cell instance $6652 r0 *1 159.33,32.76
X$6652 518 26 519 644 645 cell_1rw
* cell instance $6653 r0 *1 160.035,32.76
X$6653 520 26 521 644 645 cell_1rw
* cell instance $6654 r0 *1 160.74,32.76
X$6654 522 26 523 644 645 cell_1rw
* cell instance $6655 r0 *1 161.445,32.76
X$6655 524 26 525 644 645 cell_1rw
* cell instance $6656 r0 *1 162.15,32.76
X$6656 526 26 527 644 645 cell_1rw
* cell instance $6657 r0 *1 162.855,32.76
X$6657 528 26 529 644 645 cell_1rw
* cell instance $6658 r0 *1 163.56,32.76
X$6658 530 26 531 644 645 cell_1rw
* cell instance $6659 r0 *1 164.265,32.76
X$6659 532 26 533 644 645 cell_1rw
* cell instance $6660 r0 *1 164.97,32.76
X$6660 534 26 535 644 645 cell_1rw
* cell instance $6661 r0 *1 165.675,32.76
X$6661 536 26 537 644 645 cell_1rw
* cell instance $6662 r0 *1 166.38,32.76
X$6662 538 26 539 644 645 cell_1rw
* cell instance $6663 r0 *1 167.085,32.76
X$6663 540 26 541 644 645 cell_1rw
* cell instance $6664 r0 *1 167.79,32.76
X$6664 542 26 543 644 645 cell_1rw
* cell instance $6665 r0 *1 168.495,32.76
X$6665 544 26 545 644 645 cell_1rw
* cell instance $6666 r0 *1 169.2,32.76
X$6666 546 26 547 644 645 cell_1rw
* cell instance $6667 r0 *1 169.905,32.76
X$6667 548 26 549 644 645 cell_1rw
* cell instance $6668 r0 *1 170.61,32.76
X$6668 550 26 551 644 645 cell_1rw
* cell instance $6669 r0 *1 171.315,32.76
X$6669 552 26 553 644 645 cell_1rw
* cell instance $6670 r0 *1 172.02,32.76
X$6670 554 26 555 644 645 cell_1rw
* cell instance $6671 r0 *1 172.725,32.76
X$6671 556 26 557 644 645 cell_1rw
* cell instance $6672 r0 *1 173.43,32.76
X$6672 558 26 559 644 645 cell_1rw
* cell instance $6673 r0 *1 174.135,32.76
X$6673 560 26 561 644 645 cell_1rw
* cell instance $6674 r0 *1 174.84,32.76
X$6674 562 26 563 644 645 cell_1rw
* cell instance $6675 r0 *1 175.545,32.76
X$6675 564 26 565 644 645 cell_1rw
* cell instance $6676 r0 *1 176.25,32.76
X$6676 566 26 567 644 645 cell_1rw
* cell instance $6677 r0 *1 176.955,32.76
X$6677 568 26 569 644 645 cell_1rw
* cell instance $6678 r0 *1 177.66,32.76
X$6678 570 26 571 644 645 cell_1rw
* cell instance $6679 r0 *1 178.365,32.76
X$6679 572 26 573 644 645 cell_1rw
* cell instance $6680 r0 *1 179.07,32.76
X$6680 574 26 575 644 645 cell_1rw
* cell instance $6681 r0 *1 179.775,32.76
X$6681 576 26 577 644 645 cell_1rw
* cell instance $6682 r0 *1 180.48,32.76
X$6682 578 26 579 644 645 cell_1rw
* cell instance $6683 r0 *1 0.705,35.49
X$6683 67 27 68 644 645 cell_1rw
* cell instance $6684 r0 *1 0,35.49
X$6684 65 27 66 644 645 cell_1rw
* cell instance $6685 r0 *1 1.41,35.49
X$6685 69 27 70 644 645 cell_1rw
* cell instance $6686 r0 *1 2.115,35.49
X$6686 71 27 72 644 645 cell_1rw
* cell instance $6687 r0 *1 2.82,35.49
X$6687 73 27 74 644 645 cell_1rw
* cell instance $6688 r0 *1 3.525,35.49
X$6688 75 27 76 644 645 cell_1rw
* cell instance $6689 r0 *1 4.23,35.49
X$6689 77 27 78 644 645 cell_1rw
* cell instance $6690 r0 *1 4.935,35.49
X$6690 79 27 80 644 645 cell_1rw
* cell instance $6691 r0 *1 5.64,35.49
X$6691 81 27 82 644 645 cell_1rw
* cell instance $6692 r0 *1 6.345,35.49
X$6692 83 27 84 644 645 cell_1rw
* cell instance $6693 r0 *1 7.05,35.49
X$6693 85 27 86 644 645 cell_1rw
* cell instance $6694 r0 *1 7.755,35.49
X$6694 87 27 88 644 645 cell_1rw
* cell instance $6695 r0 *1 8.46,35.49
X$6695 89 27 90 644 645 cell_1rw
* cell instance $6696 r0 *1 9.165,35.49
X$6696 91 27 92 644 645 cell_1rw
* cell instance $6697 r0 *1 9.87,35.49
X$6697 93 27 94 644 645 cell_1rw
* cell instance $6698 r0 *1 10.575,35.49
X$6698 95 27 96 644 645 cell_1rw
* cell instance $6699 r0 *1 11.28,35.49
X$6699 97 27 98 644 645 cell_1rw
* cell instance $6700 r0 *1 11.985,35.49
X$6700 99 27 100 644 645 cell_1rw
* cell instance $6701 r0 *1 12.69,35.49
X$6701 101 27 102 644 645 cell_1rw
* cell instance $6702 r0 *1 13.395,35.49
X$6702 103 27 104 644 645 cell_1rw
* cell instance $6703 r0 *1 14.1,35.49
X$6703 105 27 106 644 645 cell_1rw
* cell instance $6704 r0 *1 14.805,35.49
X$6704 107 27 108 644 645 cell_1rw
* cell instance $6705 r0 *1 15.51,35.49
X$6705 109 27 110 644 645 cell_1rw
* cell instance $6706 r0 *1 16.215,35.49
X$6706 111 27 112 644 645 cell_1rw
* cell instance $6707 r0 *1 16.92,35.49
X$6707 113 27 114 644 645 cell_1rw
* cell instance $6708 r0 *1 17.625,35.49
X$6708 115 27 116 644 645 cell_1rw
* cell instance $6709 r0 *1 18.33,35.49
X$6709 117 27 118 644 645 cell_1rw
* cell instance $6710 r0 *1 19.035,35.49
X$6710 119 27 120 644 645 cell_1rw
* cell instance $6711 r0 *1 19.74,35.49
X$6711 121 27 122 644 645 cell_1rw
* cell instance $6712 r0 *1 20.445,35.49
X$6712 123 27 124 644 645 cell_1rw
* cell instance $6713 r0 *1 21.15,35.49
X$6713 125 27 126 644 645 cell_1rw
* cell instance $6714 r0 *1 21.855,35.49
X$6714 127 27 128 644 645 cell_1rw
* cell instance $6715 r0 *1 22.56,35.49
X$6715 129 27 130 644 645 cell_1rw
* cell instance $6716 r0 *1 23.265,35.49
X$6716 131 27 132 644 645 cell_1rw
* cell instance $6717 r0 *1 23.97,35.49
X$6717 133 27 134 644 645 cell_1rw
* cell instance $6718 r0 *1 24.675,35.49
X$6718 135 27 136 644 645 cell_1rw
* cell instance $6719 r0 *1 25.38,35.49
X$6719 137 27 138 644 645 cell_1rw
* cell instance $6720 r0 *1 26.085,35.49
X$6720 139 27 140 644 645 cell_1rw
* cell instance $6721 r0 *1 26.79,35.49
X$6721 141 27 142 644 645 cell_1rw
* cell instance $6722 r0 *1 27.495,35.49
X$6722 143 27 144 644 645 cell_1rw
* cell instance $6723 r0 *1 28.2,35.49
X$6723 145 27 146 644 645 cell_1rw
* cell instance $6724 r0 *1 28.905,35.49
X$6724 147 27 148 644 645 cell_1rw
* cell instance $6725 r0 *1 29.61,35.49
X$6725 149 27 150 644 645 cell_1rw
* cell instance $6726 r0 *1 30.315,35.49
X$6726 151 27 152 644 645 cell_1rw
* cell instance $6727 r0 *1 31.02,35.49
X$6727 153 27 154 644 645 cell_1rw
* cell instance $6728 r0 *1 31.725,35.49
X$6728 155 27 156 644 645 cell_1rw
* cell instance $6729 r0 *1 32.43,35.49
X$6729 157 27 158 644 645 cell_1rw
* cell instance $6730 r0 *1 33.135,35.49
X$6730 159 27 160 644 645 cell_1rw
* cell instance $6731 r0 *1 33.84,35.49
X$6731 161 27 162 644 645 cell_1rw
* cell instance $6732 r0 *1 34.545,35.49
X$6732 163 27 164 644 645 cell_1rw
* cell instance $6733 r0 *1 35.25,35.49
X$6733 165 27 166 644 645 cell_1rw
* cell instance $6734 r0 *1 35.955,35.49
X$6734 167 27 168 644 645 cell_1rw
* cell instance $6735 r0 *1 36.66,35.49
X$6735 169 27 170 644 645 cell_1rw
* cell instance $6736 r0 *1 37.365,35.49
X$6736 171 27 172 644 645 cell_1rw
* cell instance $6737 r0 *1 38.07,35.49
X$6737 173 27 174 644 645 cell_1rw
* cell instance $6738 r0 *1 38.775,35.49
X$6738 175 27 176 644 645 cell_1rw
* cell instance $6739 r0 *1 39.48,35.49
X$6739 177 27 178 644 645 cell_1rw
* cell instance $6740 r0 *1 40.185,35.49
X$6740 179 27 180 644 645 cell_1rw
* cell instance $6741 r0 *1 40.89,35.49
X$6741 181 27 182 644 645 cell_1rw
* cell instance $6742 r0 *1 41.595,35.49
X$6742 183 27 184 644 645 cell_1rw
* cell instance $6743 r0 *1 42.3,35.49
X$6743 185 27 186 644 645 cell_1rw
* cell instance $6744 r0 *1 43.005,35.49
X$6744 187 27 188 644 645 cell_1rw
* cell instance $6745 r0 *1 43.71,35.49
X$6745 189 27 190 644 645 cell_1rw
* cell instance $6746 r0 *1 44.415,35.49
X$6746 191 27 192 644 645 cell_1rw
* cell instance $6747 r0 *1 45.12,35.49
X$6747 193 27 194 644 645 cell_1rw
* cell instance $6748 r0 *1 45.825,35.49
X$6748 195 27 196 644 645 cell_1rw
* cell instance $6749 r0 *1 46.53,35.49
X$6749 197 27 198 644 645 cell_1rw
* cell instance $6750 r0 *1 47.235,35.49
X$6750 199 27 200 644 645 cell_1rw
* cell instance $6751 r0 *1 47.94,35.49
X$6751 201 27 202 644 645 cell_1rw
* cell instance $6752 r0 *1 48.645,35.49
X$6752 203 27 204 644 645 cell_1rw
* cell instance $6753 r0 *1 49.35,35.49
X$6753 205 27 206 644 645 cell_1rw
* cell instance $6754 r0 *1 50.055,35.49
X$6754 207 27 208 644 645 cell_1rw
* cell instance $6755 r0 *1 50.76,35.49
X$6755 209 27 210 644 645 cell_1rw
* cell instance $6756 r0 *1 51.465,35.49
X$6756 211 27 212 644 645 cell_1rw
* cell instance $6757 r0 *1 52.17,35.49
X$6757 213 27 214 644 645 cell_1rw
* cell instance $6758 r0 *1 52.875,35.49
X$6758 215 27 216 644 645 cell_1rw
* cell instance $6759 r0 *1 53.58,35.49
X$6759 217 27 218 644 645 cell_1rw
* cell instance $6760 r0 *1 54.285,35.49
X$6760 219 27 220 644 645 cell_1rw
* cell instance $6761 r0 *1 54.99,35.49
X$6761 221 27 222 644 645 cell_1rw
* cell instance $6762 r0 *1 55.695,35.49
X$6762 223 27 224 644 645 cell_1rw
* cell instance $6763 r0 *1 56.4,35.49
X$6763 225 27 226 644 645 cell_1rw
* cell instance $6764 r0 *1 57.105,35.49
X$6764 227 27 228 644 645 cell_1rw
* cell instance $6765 r0 *1 57.81,35.49
X$6765 229 27 230 644 645 cell_1rw
* cell instance $6766 r0 *1 58.515,35.49
X$6766 231 27 232 644 645 cell_1rw
* cell instance $6767 r0 *1 59.22,35.49
X$6767 233 27 234 644 645 cell_1rw
* cell instance $6768 r0 *1 59.925,35.49
X$6768 235 27 236 644 645 cell_1rw
* cell instance $6769 r0 *1 60.63,35.49
X$6769 237 27 238 644 645 cell_1rw
* cell instance $6770 r0 *1 61.335,35.49
X$6770 239 27 240 644 645 cell_1rw
* cell instance $6771 r0 *1 62.04,35.49
X$6771 241 27 242 644 645 cell_1rw
* cell instance $6772 r0 *1 62.745,35.49
X$6772 243 27 244 644 645 cell_1rw
* cell instance $6773 r0 *1 63.45,35.49
X$6773 245 27 246 644 645 cell_1rw
* cell instance $6774 r0 *1 64.155,35.49
X$6774 247 27 248 644 645 cell_1rw
* cell instance $6775 r0 *1 64.86,35.49
X$6775 249 27 250 644 645 cell_1rw
* cell instance $6776 r0 *1 65.565,35.49
X$6776 251 27 252 644 645 cell_1rw
* cell instance $6777 r0 *1 66.27,35.49
X$6777 253 27 254 644 645 cell_1rw
* cell instance $6778 r0 *1 66.975,35.49
X$6778 255 27 256 644 645 cell_1rw
* cell instance $6779 r0 *1 67.68,35.49
X$6779 257 27 258 644 645 cell_1rw
* cell instance $6780 r0 *1 68.385,35.49
X$6780 259 27 260 644 645 cell_1rw
* cell instance $6781 r0 *1 69.09,35.49
X$6781 261 27 262 644 645 cell_1rw
* cell instance $6782 r0 *1 69.795,35.49
X$6782 263 27 264 644 645 cell_1rw
* cell instance $6783 r0 *1 70.5,35.49
X$6783 265 27 266 644 645 cell_1rw
* cell instance $6784 r0 *1 71.205,35.49
X$6784 267 27 268 644 645 cell_1rw
* cell instance $6785 r0 *1 71.91,35.49
X$6785 269 27 270 644 645 cell_1rw
* cell instance $6786 r0 *1 72.615,35.49
X$6786 271 27 272 644 645 cell_1rw
* cell instance $6787 r0 *1 73.32,35.49
X$6787 273 27 274 644 645 cell_1rw
* cell instance $6788 r0 *1 74.025,35.49
X$6788 275 27 276 644 645 cell_1rw
* cell instance $6789 r0 *1 74.73,35.49
X$6789 277 27 278 644 645 cell_1rw
* cell instance $6790 r0 *1 75.435,35.49
X$6790 279 27 280 644 645 cell_1rw
* cell instance $6791 r0 *1 76.14,35.49
X$6791 281 27 282 644 645 cell_1rw
* cell instance $6792 r0 *1 76.845,35.49
X$6792 283 27 284 644 645 cell_1rw
* cell instance $6793 r0 *1 77.55,35.49
X$6793 285 27 286 644 645 cell_1rw
* cell instance $6794 r0 *1 78.255,35.49
X$6794 287 27 288 644 645 cell_1rw
* cell instance $6795 r0 *1 78.96,35.49
X$6795 289 27 290 644 645 cell_1rw
* cell instance $6796 r0 *1 79.665,35.49
X$6796 291 27 292 644 645 cell_1rw
* cell instance $6797 r0 *1 80.37,35.49
X$6797 293 27 294 644 645 cell_1rw
* cell instance $6798 r0 *1 81.075,35.49
X$6798 295 27 296 644 645 cell_1rw
* cell instance $6799 r0 *1 81.78,35.49
X$6799 297 27 298 644 645 cell_1rw
* cell instance $6800 r0 *1 82.485,35.49
X$6800 299 27 300 644 645 cell_1rw
* cell instance $6801 r0 *1 83.19,35.49
X$6801 301 27 302 644 645 cell_1rw
* cell instance $6802 r0 *1 83.895,35.49
X$6802 303 27 304 644 645 cell_1rw
* cell instance $6803 r0 *1 84.6,35.49
X$6803 305 27 306 644 645 cell_1rw
* cell instance $6804 r0 *1 85.305,35.49
X$6804 307 27 308 644 645 cell_1rw
* cell instance $6805 r0 *1 86.01,35.49
X$6805 309 27 310 644 645 cell_1rw
* cell instance $6806 r0 *1 86.715,35.49
X$6806 311 27 312 644 645 cell_1rw
* cell instance $6807 r0 *1 87.42,35.49
X$6807 313 27 314 644 645 cell_1rw
* cell instance $6808 r0 *1 88.125,35.49
X$6808 315 27 316 644 645 cell_1rw
* cell instance $6809 r0 *1 88.83,35.49
X$6809 317 27 318 644 645 cell_1rw
* cell instance $6810 r0 *1 89.535,35.49
X$6810 319 27 320 644 645 cell_1rw
* cell instance $6811 r0 *1 90.24,35.49
X$6811 321 27 323 644 645 cell_1rw
* cell instance $6812 r0 *1 90.945,35.49
X$6812 324 27 325 644 645 cell_1rw
* cell instance $6813 r0 *1 91.65,35.49
X$6813 326 27 327 644 645 cell_1rw
* cell instance $6814 r0 *1 92.355,35.49
X$6814 328 27 329 644 645 cell_1rw
* cell instance $6815 r0 *1 93.06,35.49
X$6815 330 27 331 644 645 cell_1rw
* cell instance $6816 r0 *1 93.765,35.49
X$6816 332 27 333 644 645 cell_1rw
* cell instance $6817 r0 *1 94.47,35.49
X$6817 334 27 335 644 645 cell_1rw
* cell instance $6818 r0 *1 95.175,35.49
X$6818 336 27 337 644 645 cell_1rw
* cell instance $6819 r0 *1 95.88,35.49
X$6819 338 27 339 644 645 cell_1rw
* cell instance $6820 r0 *1 96.585,35.49
X$6820 340 27 341 644 645 cell_1rw
* cell instance $6821 r0 *1 97.29,35.49
X$6821 342 27 343 644 645 cell_1rw
* cell instance $6822 r0 *1 97.995,35.49
X$6822 344 27 345 644 645 cell_1rw
* cell instance $6823 r0 *1 98.7,35.49
X$6823 346 27 347 644 645 cell_1rw
* cell instance $6824 r0 *1 99.405,35.49
X$6824 348 27 349 644 645 cell_1rw
* cell instance $6825 r0 *1 100.11,35.49
X$6825 350 27 351 644 645 cell_1rw
* cell instance $6826 r0 *1 100.815,35.49
X$6826 352 27 353 644 645 cell_1rw
* cell instance $6827 r0 *1 101.52,35.49
X$6827 354 27 355 644 645 cell_1rw
* cell instance $6828 r0 *1 102.225,35.49
X$6828 356 27 357 644 645 cell_1rw
* cell instance $6829 r0 *1 102.93,35.49
X$6829 358 27 359 644 645 cell_1rw
* cell instance $6830 r0 *1 103.635,35.49
X$6830 360 27 361 644 645 cell_1rw
* cell instance $6831 r0 *1 104.34,35.49
X$6831 362 27 363 644 645 cell_1rw
* cell instance $6832 r0 *1 105.045,35.49
X$6832 364 27 365 644 645 cell_1rw
* cell instance $6833 r0 *1 105.75,35.49
X$6833 366 27 367 644 645 cell_1rw
* cell instance $6834 r0 *1 106.455,35.49
X$6834 368 27 369 644 645 cell_1rw
* cell instance $6835 r0 *1 107.16,35.49
X$6835 370 27 371 644 645 cell_1rw
* cell instance $6836 r0 *1 107.865,35.49
X$6836 372 27 373 644 645 cell_1rw
* cell instance $6837 r0 *1 108.57,35.49
X$6837 374 27 375 644 645 cell_1rw
* cell instance $6838 r0 *1 109.275,35.49
X$6838 376 27 377 644 645 cell_1rw
* cell instance $6839 r0 *1 109.98,35.49
X$6839 378 27 379 644 645 cell_1rw
* cell instance $6840 r0 *1 110.685,35.49
X$6840 380 27 381 644 645 cell_1rw
* cell instance $6841 r0 *1 111.39,35.49
X$6841 382 27 383 644 645 cell_1rw
* cell instance $6842 r0 *1 112.095,35.49
X$6842 384 27 385 644 645 cell_1rw
* cell instance $6843 r0 *1 112.8,35.49
X$6843 386 27 387 644 645 cell_1rw
* cell instance $6844 r0 *1 113.505,35.49
X$6844 388 27 389 644 645 cell_1rw
* cell instance $6845 r0 *1 114.21,35.49
X$6845 390 27 391 644 645 cell_1rw
* cell instance $6846 r0 *1 114.915,35.49
X$6846 392 27 393 644 645 cell_1rw
* cell instance $6847 r0 *1 115.62,35.49
X$6847 394 27 395 644 645 cell_1rw
* cell instance $6848 r0 *1 116.325,35.49
X$6848 396 27 397 644 645 cell_1rw
* cell instance $6849 r0 *1 117.03,35.49
X$6849 398 27 399 644 645 cell_1rw
* cell instance $6850 r0 *1 117.735,35.49
X$6850 400 27 401 644 645 cell_1rw
* cell instance $6851 r0 *1 118.44,35.49
X$6851 402 27 403 644 645 cell_1rw
* cell instance $6852 r0 *1 119.145,35.49
X$6852 404 27 405 644 645 cell_1rw
* cell instance $6853 r0 *1 119.85,35.49
X$6853 406 27 407 644 645 cell_1rw
* cell instance $6854 r0 *1 120.555,35.49
X$6854 408 27 409 644 645 cell_1rw
* cell instance $6855 r0 *1 121.26,35.49
X$6855 410 27 411 644 645 cell_1rw
* cell instance $6856 r0 *1 121.965,35.49
X$6856 412 27 413 644 645 cell_1rw
* cell instance $6857 r0 *1 122.67,35.49
X$6857 414 27 415 644 645 cell_1rw
* cell instance $6858 r0 *1 123.375,35.49
X$6858 416 27 417 644 645 cell_1rw
* cell instance $6859 r0 *1 124.08,35.49
X$6859 418 27 419 644 645 cell_1rw
* cell instance $6860 r0 *1 124.785,35.49
X$6860 420 27 421 644 645 cell_1rw
* cell instance $6861 r0 *1 125.49,35.49
X$6861 422 27 423 644 645 cell_1rw
* cell instance $6862 r0 *1 126.195,35.49
X$6862 424 27 425 644 645 cell_1rw
* cell instance $6863 r0 *1 126.9,35.49
X$6863 426 27 427 644 645 cell_1rw
* cell instance $6864 r0 *1 127.605,35.49
X$6864 428 27 429 644 645 cell_1rw
* cell instance $6865 r0 *1 128.31,35.49
X$6865 430 27 431 644 645 cell_1rw
* cell instance $6866 r0 *1 129.015,35.49
X$6866 432 27 433 644 645 cell_1rw
* cell instance $6867 r0 *1 129.72,35.49
X$6867 434 27 435 644 645 cell_1rw
* cell instance $6868 r0 *1 130.425,35.49
X$6868 436 27 437 644 645 cell_1rw
* cell instance $6869 r0 *1 131.13,35.49
X$6869 438 27 439 644 645 cell_1rw
* cell instance $6870 r0 *1 131.835,35.49
X$6870 440 27 441 644 645 cell_1rw
* cell instance $6871 r0 *1 132.54,35.49
X$6871 442 27 443 644 645 cell_1rw
* cell instance $6872 r0 *1 133.245,35.49
X$6872 444 27 445 644 645 cell_1rw
* cell instance $6873 r0 *1 133.95,35.49
X$6873 446 27 447 644 645 cell_1rw
* cell instance $6874 r0 *1 134.655,35.49
X$6874 448 27 449 644 645 cell_1rw
* cell instance $6875 r0 *1 135.36,35.49
X$6875 450 27 451 644 645 cell_1rw
* cell instance $6876 r0 *1 136.065,35.49
X$6876 452 27 453 644 645 cell_1rw
* cell instance $6877 r0 *1 136.77,35.49
X$6877 454 27 455 644 645 cell_1rw
* cell instance $6878 r0 *1 137.475,35.49
X$6878 456 27 457 644 645 cell_1rw
* cell instance $6879 r0 *1 138.18,35.49
X$6879 458 27 459 644 645 cell_1rw
* cell instance $6880 r0 *1 138.885,35.49
X$6880 460 27 461 644 645 cell_1rw
* cell instance $6881 r0 *1 139.59,35.49
X$6881 462 27 463 644 645 cell_1rw
* cell instance $6882 r0 *1 140.295,35.49
X$6882 464 27 465 644 645 cell_1rw
* cell instance $6883 r0 *1 141,35.49
X$6883 466 27 467 644 645 cell_1rw
* cell instance $6884 r0 *1 141.705,35.49
X$6884 468 27 469 644 645 cell_1rw
* cell instance $6885 r0 *1 142.41,35.49
X$6885 470 27 471 644 645 cell_1rw
* cell instance $6886 r0 *1 143.115,35.49
X$6886 472 27 473 644 645 cell_1rw
* cell instance $6887 r0 *1 143.82,35.49
X$6887 474 27 475 644 645 cell_1rw
* cell instance $6888 r0 *1 144.525,35.49
X$6888 476 27 477 644 645 cell_1rw
* cell instance $6889 r0 *1 145.23,35.49
X$6889 478 27 479 644 645 cell_1rw
* cell instance $6890 r0 *1 145.935,35.49
X$6890 480 27 481 644 645 cell_1rw
* cell instance $6891 r0 *1 146.64,35.49
X$6891 482 27 483 644 645 cell_1rw
* cell instance $6892 r0 *1 147.345,35.49
X$6892 484 27 485 644 645 cell_1rw
* cell instance $6893 r0 *1 148.05,35.49
X$6893 486 27 487 644 645 cell_1rw
* cell instance $6894 r0 *1 148.755,35.49
X$6894 488 27 489 644 645 cell_1rw
* cell instance $6895 r0 *1 149.46,35.49
X$6895 490 27 491 644 645 cell_1rw
* cell instance $6896 r0 *1 150.165,35.49
X$6896 492 27 493 644 645 cell_1rw
* cell instance $6897 r0 *1 150.87,35.49
X$6897 494 27 495 644 645 cell_1rw
* cell instance $6898 r0 *1 151.575,35.49
X$6898 496 27 497 644 645 cell_1rw
* cell instance $6899 r0 *1 152.28,35.49
X$6899 498 27 499 644 645 cell_1rw
* cell instance $6900 r0 *1 152.985,35.49
X$6900 500 27 501 644 645 cell_1rw
* cell instance $6901 r0 *1 153.69,35.49
X$6901 502 27 503 644 645 cell_1rw
* cell instance $6902 r0 *1 154.395,35.49
X$6902 504 27 505 644 645 cell_1rw
* cell instance $6903 r0 *1 155.1,35.49
X$6903 506 27 507 644 645 cell_1rw
* cell instance $6904 r0 *1 155.805,35.49
X$6904 508 27 509 644 645 cell_1rw
* cell instance $6905 r0 *1 156.51,35.49
X$6905 510 27 511 644 645 cell_1rw
* cell instance $6906 r0 *1 157.215,35.49
X$6906 512 27 513 644 645 cell_1rw
* cell instance $6907 r0 *1 157.92,35.49
X$6907 514 27 515 644 645 cell_1rw
* cell instance $6908 r0 *1 158.625,35.49
X$6908 516 27 517 644 645 cell_1rw
* cell instance $6909 r0 *1 159.33,35.49
X$6909 518 27 519 644 645 cell_1rw
* cell instance $6910 r0 *1 160.035,35.49
X$6910 520 27 521 644 645 cell_1rw
* cell instance $6911 r0 *1 160.74,35.49
X$6911 522 27 523 644 645 cell_1rw
* cell instance $6912 r0 *1 161.445,35.49
X$6912 524 27 525 644 645 cell_1rw
* cell instance $6913 r0 *1 162.15,35.49
X$6913 526 27 527 644 645 cell_1rw
* cell instance $6914 r0 *1 162.855,35.49
X$6914 528 27 529 644 645 cell_1rw
* cell instance $6915 r0 *1 163.56,35.49
X$6915 530 27 531 644 645 cell_1rw
* cell instance $6916 r0 *1 164.265,35.49
X$6916 532 27 533 644 645 cell_1rw
* cell instance $6917 r0 *1 164.97,35.49
X$6917 534 27 535 644 645 cell_1rw
* cell instance $6918 r0 *1 165.675,35.49
X$6918 536 27 537 644 645 cell_1rw
* cell instance $6919 r0 *1 166.38,35.49
X$6919 538 27 539 644 645 cell_1rw
* cell instance $6920 r0 *1 167.085,35.49
X$6920 540 27 541 644 645 cell_1rw
* cell instance $6921 r0 *1 167.79,35.49
X$6921 542 27 543 644 645 cell_1rw
* cell instance $6922 r0 *1 168.495,35.49
X$6922 544 27 545 644 645 cell_1rw
* cell instance $6923 r0 *1 169.2,35.49
X$6923 546 27 547 644 645 cell_1rw
* cell instance $6924 r0 *1 169.905,35.49
X$6924 548 27 549 644 645 cell_1rw
* cell instance $6925 r0 *1 170.61,35.49
X$6925 550 27 551 644 645 cell_1rw
* cell instance $6926 r0 *1 171.315,35.49
X$6926 552 27 553 644 645 cell_1rw
* cell instance $6927 r0 *1 172.02,35.49
X$6927 554 27 555 644 645 cell_1rw
* cell instance $6928 r0 *1 172.725,35.49
X$6928 556 27 557 644 645 cell_1rw
* cell instance $6929 r0 *1 173.43,35.49
X$6929 558 27 559 644 645 cell_1rw
* cell instance $6930 r0 *1 174.135,35.49
X$6930 560 27 561 644 645 cell_1rw
* cell instance $6931 r0 *1 174.84,35.49
X$6931 562 27 563 644 645 cell_1rw
* cell instance $6932 r0 *1 175.545,35.49
X$6932 564 27 565 644 645 cell_1rw
* cell instance $6933 r0 *1 176.25,35.49
X$6933 566 27 567 644 645 cell_1rw
* cell instance $6934 r0 *1 176.955,35.49
X$6934 568 27 569 644 645 cell_1rw
* cell instance $6935 r0 *1 177.66,35.49
X$6935 570 27 571 644 645 cell_1rw
* cell instance $6936 r0 *1 178.365,35.49
X$6936 572 27 573 644 645 cell_1rw
* cell instance $6937 r0 *1 179.07,35.49
X$6937 574 27 575 644 645 cell_1rw
* cell instance $6938 r0 *1 179.775,35.49
X$6938 576 27 577 644 645 cell_1rw
* cell instance $6939 r0 *1 180.48,35.49
X$6939 578 27 579 644 645 cell_1rw
* cell instance $6940 m0 *1 0.705,38.22
X$6940 67 28 68 644 645 cell_1rw
* cell instance $6941 m0 *1 0,38.22
X$6941 65 28 66 644 645 cell_1rw
* cell instance $6942 m0 *1 1.41,38.22
X$6942 69 28 70 644 645 cell_1rw
* cell instance $6943 m0 *1 2.115,38.22
X$6943 71 28 72 644 645 cell_1rw
* cell instance $6944 m0 *1 2.82,38.22
X$6944 73 28 74 644 645 cell_1rw
* cell instance $6945 m0 *1 3.525,38.22
X$6945 75 28 76 644 645 cell_1rw
* cell instance $6946 m0 *1 4.23,38.22
X$6946 77 28 78 644 645 cell_1rw
* cell instance $6947 m0 *1 4.935,38.22
X$6947 79 28 80 644 645 cell_1rw
* cell instance $6948 m0 *1 5.64,38.22
X$6948 81 28 82 644 645 cell_1rw
* cell instance $6949 m0 *1 6.345,38.22
X$6949 83 28 84 644 645 cell_1rw
* cell instance $6950 m0 *1 7.05,38.22
X$6950 85 28 86 644 645 cell_1rw
* cell instance $6951 m0 *1 7.755,38.22
X$6951 87 28 88 644 645 cell_1rw
* cell instance $6952 m0 *1 8.46,38.22
X$6952 89 28 90 644 645 cell_1rw
* cell instance $6953 m0 *1 9.165,38.22
X$6953 91 28 92 644 645 cell_1rw
* cell instance $6954 m0 *1 9.87,38.22
X$6954 93 28 94 644 645 cell_1rw
* cell instance $6955 m0 *1 10.575,38.22
X$6955 95 28 96 644 645 cell_1rw
* cell instance $6956 m0 *1 11.28,38.22
X$6956 97 28 98 644 645 cell_1rw
* cell instance $6957 m0 *1 11.985,38.22
X$6957 99 28 100 644 645 cell_1rw
* cell instance $6958 m0 *1 12.69,38.22
X$6958 101 28 102 644 645 cell_1rw
* cell instance $6959 m0 *1 13.395,38.22
X$6959 103 28 104 644 645 cell_1rw
* cell instance $6960 m0 *1 14.1,38.22
X$6960 105 28 106 644 645 cell_1rw
* cell instance $6961 m0 *1 14.805,38.22
X$6961 107 28 108 644 645 cell_1rw
* cell instance $6962 m0 *1 15.51,38.22
X$6962 109 28 110 644 645 cell_1rw
* cell instance $6963 m0 *1 16.215,38.22
X$6963 111 28 112 644 645 cell_1rw
* cell instance $6964 m0 *1 16.92,38.22
X$6964 113 28 114 644 645 cell_1rw
* cell instance $6965 m0 *1 17.625,38.22
X$6965 115 28 116 644 645 cell_1rw
* cell instance $6966 m0 *1 18.33,38.22
X$6966 117 28 118 644 645 cell_1rw
* cell instance $6967 m0 *1 19.035,38.22
X$6967 119 28 120 644 645 cell_1rw
* cell instance $6968 m0 *1 19.74,38.22
X$6968 121 28 122 644 645 cell_1rw
* cell instance $6969 m0 *1 20.445,38.22
X$6969 123 28 124 644 645 cell_1rw
* cell instance $6970 m0 *1 21.15,38.22
X$6970 125 28 126 644 645 cell_1rw
* cell instance $6971 m0 *1 21.855,38.22
X$6971 127 28 128 644 645 cell_1rw
* cell instance $6972 m0 *1 22.56,38.22
X$6972 129 28 130 644 645 cell_1rw
* cell instance $6973 m0 *1 23.265,38.22
X$6973 131 28 132 644 645 cell_1rw
* cell instance $6974 m0 *1 23.97,38.22
X$6974 133 28 134 644 645 cell_1rw
* cell instance $6975 m0 *1 24.675,38.22
X$6975 135 28 136 644 645 cell_1rw
* cell instance $6976 m0 *1 25.38,38.22
X$6976 137 28 138 644 645 cell_1rw
* cell instance $6977 m0 *1 26.085,38.22
X$6977 139 28 140 644 645 cell_1rw
* cell instance $6978 m0 *1 26.79,38.22
X$6978 141 28 142 644 645 cell_1rw
* cell instance $6979 m0 *1 27.495,38.22
X$6979 143 28 144 644 645 cell_1rw
* cell instance $6980 m0 *1 28.2,38.22
X$6980 145 28 146 644 645 cell_1rw
* cell instance $6981 m0 *1 28.905,38.22
X$6981 147 28 148 644 645 cell_1rw
* cell instance $6982 m0 *1 29.61,38.22
X$6982 149 28 150 644 645 cell_1rw
* cell instance $6983 m0 *1 30.315,38.22
X$6983 151 28 152 644 645 cell_1rw
* cell instance $6984 m0 *1 31.02,38.22
X$6984 153 28 154 644 645 cell_1rw
* cell instance $6985 m0 *1 31.725,38.22
X$6985 155 28 156 644 645 cell_1rw
* cell instance $6986 m0 *1 32.43,38.22
X$6986 157 28 158 644 645 cell_1rw
* cell instance $6987 m0 *1 33.135,38.22
X$6987 159 28 160 644 645 cell_1rw
* cell instance $6988 m0 *1 33.84,38.22
X$6988 161 28 162 644 645 cell_1rw
* cell instance $6989 m0 *1 34.545,38.22
X$6989 163 28 164 644 645 cell_1rw
* cell instance $6990 m0 *1 35.25,38.22
X$6990 165 28 166 644 645 cell_1rw
* cell instance $6991 m0 *1 35.955,38.22
X$6991 167 28 168 644 645 cell_1rw
* cell instance $6992 m0 *1 36.66,38.22
X$6992 169 28 170 644 645 cell_1rw
* cell instance $6993 m0 *1 37.365,38.22
X$6993 171 28 172 644 645 cell_1rw
* cell instance $6994 m0 *1 38.07,38.22
X$6994 173 28 174 644 645 cell_1rw
* cell instance $6995 m0 *1 38.775,38.22
X$6995 175 28 176 644 645 cell_1rw
* cell instance $6996 m0 *1 39.48,38.22
X$6996 177 28 178 644 645 cell_1rw
* cell instance $6997 m0 *1 40.185,38.22
X$6997 179 28 180 644 645 cell_1rw
* cell instance $6998 m0 *1 40.89,38.22
X$6998 181 28 182 644 645 cell_1rw
* cell instance $6999 m0 *1 41.595,38.22
X$6999 183 28 184 644 645 cell_1rw
* cell instance $7000 m0 *1 42.3,38.22
X$7000 185 28 186 644 645 cell_1rw
* cell instance $7001 m0 *1 43.005,38.22
X$7001 187 28 188 644 645 cell_1rw
* cell instance $7002 m0 *1 43.71,38.22
X$7002 189 28 190 644 645 cell_1rw
* cell instance $7003 m0 *1 44.415,38.22
X$7003 191 28 192 644 645 cell_1rw
* cell instance $7004 m0 *1 45.12,38.22
X$7004 193 28 194 644 645 cell_1rw
* cell instance $7005 m0 *1 45.825,38.22
X$7005 195 28 196 644 645 cell_1rw
* cell instance $7006 m0 *1 46.53,38.22
X$7006 197 28 198 644 645 cell_1rw
* cell instance $7007 m0 *1 47.235,38.22
X$7007 199 28 200 644 645 cell_1rw
* cell instance $7008 m0 *1 47.94,38.22
X$7008 201 28 202 644 645 cell_1rw
* cell instance $7009 m0 *1 48.645,38.22
X$7009 203 28 204 644 645 cell_1rw
* cell instance $7010 m0 *1 49.35,38.22
X$7010 205 28 206 644 645 cell_1rw
* cell instance $7011 m0 *1 50.055,38.22
X$7011 207 28 208 644 645 cell_1rw
* cell instance $7012 m0 *1 50.76,38.22
X$7012 209 28 210 644 645 cell_1rw
* cell instance $7013 m0 *1 51.465,38.22
X$7013 211 28 212 644 645 cell_1rw
* cell instance $7014 m0 *1 52.17,38.22
X$7014 213 28 214 644 645 cell_1rw
* cell instance $7015 m0 *1 52.875,38.22
X$7015 215 28 216 644 645 cell_1rw
* cell instance $7016 m0 *1 53.58,38.22
X$7016 217 28 218 644 645 cell_1rw
* cell instance $7017 m0 *1 54.285,38.22
X$7017 219 28 220 644 645 cell_1rw
* cell instance $7018 m0 *1 54.99,38.22
X$7018 221 28 222 644 645 cell_1rw
* cell instance $7019 m0 *1 55.695,38.22
X$7019 223 28 224 644 645 cell_1rw
* cell instance $7020 m0 *1 56.4,38.22
X$7020 225 28 226 644 645 cell_1rw
* cell instance $7021 m0 *1 57.105,38.22
X$7021 227 28 228 644 645 cell_1rw
* cell instance $7022 m0 *1 57.81,38.22
X$7022 229 28 230 644 645 cell_1rw
* cell instance $7023 m0 *1 58.515,38.22
X$7023 231 28 232 644 645 cell_1rw
* cell instance $7024 m0 *1 59.22,38.22
X$7024 233 28 234 644 645 cell_1rw
* cell instance $7025 m0 *1 59.925,38.22
X$7025 235 28 236 644 645 cell_1rw
* cell instance $7026 m0 *1 60.63,38.22
X$7026 237 28 238 644 645 cell_1rw
* cell instance $7027 m0 *1 61.335,38.22
X$7027 239 28 240 644 645 cell_1rw
* cell instance $7028 m0 *1 62.04,38.22
X$7028 241 28 242 644 645 cell_1rw
* cell instance $7029 m0 *1 62.745,38.22
X$7029 243 28 244 644 645 cell_1rw
* cell instance $7030 m0 *1 63.45,38.22
X$7030 245 28 246 644 645 cell_1rw
* cell instance $7031 m0 *1 64.155,38.22
X$7031 247 28 248 644 645 cell_1rw
* cell instance $7032 m0 *1 64.86,38.22
X$7032 249 28 250 644 645 cell_1rw
* cell instance $7033 m0 *1 65.565,38.22
X$7033 251 28 252 644 645 cell_1rw
* cell instance $7034 m0 *1 66.27,38.22
X$7034 253 28 254 644 645 cell_1rw
* cell instance $7035 m0 *1 66.975,38.22
X$7035 255 28 256 644 645 cell_1rw
* cell instance $7036 m0 *1 67.68,38.22
X$7036 257 28 258 644 645 cell_1rw
* cell instance $7037 m0 *1 68.385,38.22
X$7037 259 28 260 644 645 cell_1rw
* cell instance $7038 m0 *1 69.09,38.22
X$7038 261 28 262 644 645 cell_1rw
* cell instance $7039 m0 *1 69.795,38.22
X$7039 263 28 264 644 645 cell_1rw
* cell instance $7040 m0 *1 70.5,38.22
X$7040 265 28 266 644 645 cell_1rw
* cell instance $7041 m0 *1 71.205,38.22
X$7041 267 28 268 644 645 cell_1rw
* cell instance $7042 m0 *1 71.91,38.22
X$7042 269 28 270 644 645 cell_1rw
* cell instance $7043 m0 *1 72.615,38.22
X$7043 271 28 272 644 645 cell_1rw
* cell instance $7044 m0 *1 73.32,38.22
X$7044 273 28 274 644 645 cell_1rw
* cell instance $7045 m0 *1 74.025,38.22
X$7045 275 28 276 644 645 cell_1rw
* cell instance $7046 m0 *1 74.73,38.22
X$7046 277 28 278 644 645 cell_1rw
* cell instance $7047 m0 *1 75.435,38.22
X$7047 279 28 280 644 645 cell_1rw
* cell instance $7048 m0 *1 76.14,38.22
X$7048 281 28 282 644 645 cell_1rw
* cell instance $7049 m0 *1 76.845,38.22
X$7049 283 28 284 644 645 cell_1rw
* cell instance $7050 m0 *1 77.55,38.22
X$7050 285 28 286 644 645 cell_1rw
* cell instance $7051 m0 *1 78.255,38.22
X$7051 287 28 288 644 645 cell_1rw
* cell instance $7052 m0 *1 78.96,38.22
X$7052 289 28 290 644 645 cell_1rw
* cell instance $7053 m0 *1 79.665,38.22
X$7053 291 28 292 644 645 cell_1rw
* cell instance $7054 m0 *1 80.37,38.22
X$7054 293 28 294 644 645 cell_1rw
* cell instance $7055 m0 *1 81.075,38.22
X$7055 295 28 296 644 645 cell_1rw
* cell instance $7056 m0 *1 81.78,38.22
X$7056 297 28 298 644 645 cell_1rw
* cell instance $7057 m0 *1 82.485,38.22
X$7057 299 28 300 644 645 cell_1rw
* cell instance $7058 m0 *1 83.19,38.22
X$7058 301 28 302 644 645 cell_1rw
* cell instance $7059 m0 *1 83.895,38.22
X$7059 303 28 304 644 645 cell_1rw
* cell instance $7060 m0 *1 84.6,38.22
X$7060 305 28 306 644 645 cell_1rw
* cell instance $7061 m0 *1 85.305,38.22
X$7061 307 28 308 644 645 cell_1rw
* cell instance $7062 m0 *1 86.01,38.22
X$7062 309 28 310 644 645 cell_1rw
* cell instance $7063 m0 *1 86.715,38.22
X$7063 311 28 312 644 645 cell_1rw
* cell instance $7064 m0 *1 87.42,38.22
X$7064 313 28 314 644 645 cell_1rw
* cell instance $7065 m0 *1 88.125,38.22
X$7065 315 28 316 644 645 cell_1rw
* cell instance $7066 m0 *1 88.83,38.22
X$7066 317 28 318 644 645 cell_1rw
* cell instance $7067 m0 *1 89.535,38.22
X$7067 319 28 320 644 645 cell_1rw
* cell instance $7068 m0 *1 90.24,38.22
X$7068 321 28 323 644 645 cell_1rw
* cell instance $7069 m0 *1 90.945,38.22
X$7069 324 28 325 644 645 cell_1rw
* cell instance $7070 m0 *1 91.65,38.22
X$7070 326 28 327 644 645 cell_1rw
* cell instance $7071 m0 *1 92.355,38.22
X$7071 328 28 329 644 645 cell_1rw
* cell instance $7072 m0 *1 93.06,38.22
X$7072 330 28 331 644 645 cell_1rw
* cell instance $7073 m0 *1 93.765,38.22
X$7073 332 28 333 644 645 cell_1rw
* cell instance $7074 m0 *1 94.47,38.22
X$7074 334 28 335 644 645 cell_1rw
* cell instance $7075 m0 *1 95.175,38.22
X$7075 336 28 337 644 645 cell_1rw
* cell instance $7076 m0 *1 95.88,38.22
X$7076 338 28 339 644 645 cell_1rw
* cell instance $7077 m0 *1 96.585,38.22
X$7077 340 28 341 644 645 cell_1rw
* cell instance $7078 m0 *1 97.29,38.22
X$7078 342 28 343 644 645 cell_1rw
* cell instance $7079 m0 *1 97.995,38.22
X$7079 344 28 345 644 645 cell_1rw
* cell instance $7080 m0 *1 98.7,38.22
X$7080 346 28 347 644 645 cell_1rw
* cell instance $7081 m0 *1 99.405,38.22
X$7081 348 28 349 644 645 cell_1rw
* cell instance $7082 m0 *1 100.11,38.22
X$7082 350 28 351 644 645 cell_1rw
* cell instance $7083 m0 *1 100.815,38.22
X$7083 352 28 353 644 645 cell_1rw
* cell instance $7084 m0 *1 101.52,38.22
X$7084 354 28 355 644 645 cell_1rw
* cell instance $7085 m0 *1 102.225,38.22
X$7085 356 28 357 644 645 cell_1rw
* cell instance $7086 m0 *1 102.93,38.22
X$7086 358 28 359 644 645 cell_1rw
* cell instance $7087 m0 *1 103.635,38.22
X$7087 360 28 361 644 645 cell_1rw
* cell instance $7088 m0 *1 104.34,38.22
X$7088 362 28 363 644 645 cell_1rw
* cell instance $7089 m0 *1 105.045,38.22
X$7089 364 28 365 644 645 cell_1rw
* cell instance $7090 m0 *1 105.75,38.22
X$7090 366 28 367 644 645 cell_1rw
* cell instance $7091 m0 *1 106.455,38.22
X$7091 368 28 369 644 645 cell_1rw
* cell instance $7092 m0 *1 107.16,38.22
X$7092 370 28 371 644 645 cell_1rw
* cell instance $7093 m0 *1 107.865,38.22
X$7093 372 28 373 644 645 cell_1rw
* cell instance $7094 m0 *1 108.57,38.22
X$7094 374 28 375 644 645 cell_1rw
* cell instance $7095 m0 *1 109.275,38.22
X$7095 376 28 377 644 645 cell_1rw
* cell instance $7096 m0 *1 109.98,38.22
X$7096 378 28 379 644 645 cell_1rw
* cell instance $7097 m0 *1 110.685,38.22
X$7097 380 28 381 644 645 cell_1rw
* cell instance $7098 m0 *1 111.39,38.22
X$7098 382 28 383 644 645 cell_1rw
* cell instance $7099 m0 *1 112.095,38.22
X$7099 384 28 385 644 645 cell_1rw
* cell instance $7100 m0 *1 112.8,38.22
X$7100 386 28 387 644 645 cell_1rw
* cell instance $7101 m0 *1 113.505,38.22
X$7101 388 28 389 644 645 cell_1rw
* cell instance $7102 m0 *1 114.21,38.22
X$7102 390 28 391 644 645 cell_1rw
* cell instance $7103 m0 *1 114.915,38.22
X$7103 392 28 393 644 645 cell_1rw
* cell instance $7104 m0 *1 115.62,38.22
X$7104 394 28 395 644 645 cell_1rw
* cell instance $7105 m0 *1 116.325,38.22
X$7105 396 28 397 644 645 cell_1rw
* cell instance $7106 m0 *1 117.03,38.22
X$7106 398 28 399 644 645 cell_1rw
* cell instance $7107 m0 *1 117.735,38.22
X$7107 400 28 401 644 645 cell_1rw
* cell instance $7108 m0 *1 118.44,38.22
X$7108 402 28 403 644 645 cell_1rw
* cell instance $7109 m0 *1 119.145,38.22
X$7109 404 28 405 644 645 cell_1rw
* cell instance $7110 m0 *1 119.85,38.22
X$7110 406 28 407 644 645 cell_1rw
* cell instance $7111 m0 *1 120.555,38.22
X$7111 408 28 409 644 645 cell_1rw
* cell instance $7112 m0 *1 121.26,38.22
X$7112 410 28 411 644 645 cell_1rw
* cell instance $7113 m0 *1 121.965,38.22
X$7113 412 28 413 644 645 cell_1rw
* cell instance $7114 m0 *1 122.67,38.22
X$7114 414 28 415 644 645 cell_1rw
* cell instance $7115 m0 *1 123.375,38.22
X$7115 416 28 417 644 645 cell_1rw
* cell instance $7116 m0 *1 124.08,38.22
X$7116 418 28 419 644 645 cell_1rw
* cell instance $7117 m0 *1 124.785,38.22
X$7117 420 28 421 644 645 cell_1rw
* cell instance $7118 m0 *1 125.49,38.22
X$7118 422 28 423 644 645 cell_1rw
* cell instance $7119 m0 *1 126.195,38.22
X$7119 424 28 425 644 645 cell_1rw
* cell instance $7120 m0 *1 126.9,38.22
X$7120 426 28 427 644 645 cell_1rw
* cell instance $7121 m0 *1 127.605,38.22
X$7121 428 28 429 644 645 cell_1rw
* cell instance $7122 m0 *1 128.31,38.22
X$7122 430 28 431 644 645 cell_1rw
* cell instance $7123 m0 *1 129.015,38.22
X$7123 432 28 433 644 645 cell_1rw
* cell instance $7124 m0 *1 129.72,38.22
X$7124 434 28 435 644 645 cell_1rw
* cell instance $7125 m0 *1 130.425,38.22
X$7125 436 28 437 644 645 cell_1rw
* cell instance $7126 m0 *1 131.13,38.22
X$7126 438 28 439 644 645 cell_1rw
* cell instance $7127 m0 *1 131.835,38.22
X$7127 440 28 441 644 645 cell_1rw
* cell instance $7128 m0 *1 132.54,38.22
X$7128 442 28 443 644 645 cell_1rw
* cell instance $7129 m0 *1 133.245,38.22
X$7129 444 28 445 644 645 cell_1rw
* cell instance $7130 m0 *1 133.95,38.22
X$7130 446 28 447 644 645 cell_1rw
* cell instance $7131 m0 *1 134.655,38.22
X$7131 448 28 449 644 645 cell_1rw
* cell instance $7132 m0 *1 135.36,38.22
X$7132 450 28 451 644 645 cell_1rw
* cell instance $7133 m0 *1 136.065,38.22
X$7133 452 28 453 644 645 cell_1rw
* cell instance $7134 m0 *1 136.77,38.22
X$7134 454 28 455 644 645 cell_1rw
* cell instance $7135 m0 *1 137.475,38.22
X$7135 456 28 457 644 645 cell_1rw
* cell instance $7136 m0 *1 138.18,38.22
X$7136 458 28 459 644 645 cell_1rw
* cell instance $7137 m0 *1 138.885,38.22
X$7137 460 28 461 644 645 cell_1rw
* cell instance $7138 m0 *1 139.59,38.22
X$7138 462 28 463 644 645 cell_1rw
* cell instance $7139 m0 *1 140.295,38.22
X$7139 464 28 465 644 645 cell_1rw
* cell instance $7140 m0 *1 141,38.22
X$7140 466 28 467 644 645 cell_1rw
* cell instance $7141 m0 *1 141.705,38.22
X$7141 468 28 469 644 645 cell_1rw
* cell instance $7142 m0 *1 142.41,38.22
X$7142 470 28 471 644 645 cell_1rw
* cell instance $7143 m0 *1 143.115,38.22
X$7143 472 28 473 644 645 cell_1rw
* cell instance $7144 m0 *1 143.82,38.22
X$7144 474 28 475 644 645 cell_1rw
* cell instance $7145 m0 *1 144.525,38.22
X$7145 476 28 477 644 645 cell_1rw
* cell instance $7146 m0 *1 145.23,38.22
X$7146 478 28 479 644 645 cell_1rw
* cell instance $7147 m0 *1 145.935,38.22
X$7147 480 28 481 644 645 cell_1rw
* cell instance $7148 m0 *1 146.64,38.22
X$7148 482 28 483 644 645 cell_1rw
* cell instance $7149 m0 *1 147.345,38.22
X$7149 484 28 485 644 645 cell_1rw
* cell instance $7150 m0 *1 148.05,38.22
X$7150 486 28 487 644 645 cell_1rw
* cell instance $7151 m0 *1 148.755,38.22
X$7151 488 28 489 644 645 cell_1rw
* cell instance $7152 m0 *1 149.46,38.22
X$7152 490 28 491 644 645 cell_1rw
* cell instance $7153 m0 *1 150.165,38.22
X$7153 492 28 493 644 645 cell_1rw
* cell instance $7154 m0 *1 150.87,38.22
X$7154 494 28 495 644 645 cell_1rw
* cell instance $7155 m0 *1 151.575,38.22
X$7155 496 28 497 644 645 cell_1rw
* cell instance $7156 m0 *1 152.28,38.22
X$7156 498 28 499 644 645 cell_1rw
* cell instance $7157 m0 *1 152.985,38.22
X$7157 500 28 501 644 645 cell_1rw
* cell instance $7158 m0 *1 153.69,38.22
X$7158 502 28 503 644 645 cell_1rw
* cell instance $7159 m0 *1 154.395,38.22
X$7159 504 28 505 644 645 cell_1rw
* cell instance $7160 m0 *1 155.1,38.22
X$7160 506 28 507 644 645 cell_1rw
* cell instance $7161 m0 *1 155.805,38.22
X$7161 508 28 509 644 645 cell_1rw
* cell instance $7162 m0 *1 156.51,38.22
X$7162 510 28 511 644 645 cell_1rw
* cell instance $7163 m0 *1 157.215,38.22
X$7163 512 28 513 644 645 cell_1rw
* cell instance $7164 m0 *1 157.92,38.22
X$7164 514 28 515 644 645 cell_1rw
* cell instance $7165 m0 *1 158.625,38.22
X$7165 516 28 517 644 645 cell_1rw
* cell instance $7166 m0 *1 159.33,38.22
X$7166 518 28 519 644 645 cell_1rw
* cell instance $7167 m0 *1 160.035,38.22
X$7167 520 28 521 644 645 cell_1rw
* cell instance $7168 m0 *1 160.74,38.22
X$7168 522 28 523 644 645 cell_1rw
* cell instance $7169 m0 *1 161.445,38.22
X$7169 524 28 525 644 645 cell_1rw
* cell instance $7170 m0 *1 162.15,38.22
X$7170 526 28 527 644 645 cell_1rw
* cell instance $7171 m0 *1 162.855,38.22
X$7171 528 28 529 644 645 cell_1rw
* cell instance $7172 m0 *1 163.56,38.22
X$7172 530 28 531 644 645 cell_1rw
* cell instance $7173 m0 *1 164.265,38.22
X$7173 532 28 533 644 645 cell_1rw
* cell instance $7174 m0 *1 164.97,38.22
X$7174 534 28 535 644 645 cell_1rw
* cell instance $7175 m0 *1 165.675,38.22
X$7175 536 28 537 644 645 cell_1rw
* cell instance $7176 m0 *1 166.38,38.22
X$7176 538 28 539 644 645 cell_1rw
* cell instance $7177 m0 *1 167.085,38.22
X$7177 540 28 541 644 645 cell_1rw
* cell instance $7178 m0 *1 167.79,38.22
X$7178 542 28 543 644 645 cell_1rw
* cell instance $7179 m0 *1 168.495,38.22
X$7179 544 28 545 644 645 cell_1rw
* cell instance $7180 m0 *1 169.2,38.22
X$7180 546 28 547 644 645 cell_1rw
* cell instance $7181 m0 *1 169.905,38.22
X$7181 548 28 549 644 645 cell_1rw
* cell instance $7182 m0 *1 170.61,38.22
X$7182 550 28 551 644 645 cell_1rw
* cell instance $7183 m0 *1 171.315,38.22
X$7183 552 28 553 644 645 cell_1rw
* cell instance $7184 m0 *1 172.02,38.22
X$7184 554 28 555 644 645 cell_1rw
* cell instance $7185 m0 *1 172.725,38.22
X$7185 556 28 557 644 645 cell_1rw
* cell instance $7186 m0 *1 173.43,38.22
X$7186 558 28 559 644 645 cell_1rw
* cell instance $7187 m0 *1 174.135,38.22
X$7187 560 28 561 644 645 cell_1rw
* cell instance $7188 m0 *1 174.84,38.22
X$7188 562 28 563 644 645 cell_1rw
* cell instance $7189 m0 *1 175.545,38.22
X$7189 564 28 565 644 645 cell_1rw
* cell instance $7190 m0 *1 176.25,38.22
X$7190 566 28 567 644 645 cell_1rw
* cell instance $7191 m0 *1 176.955,38.22
X$7191 568 28 569 644 645 cell_1rw
* cell instance $7192 m0 *1 177.66,38.22
X$7192 570 28 571 644 645 cell_1rw
* cell instance $7193 m0 *1 178.365,38.22
X$7193 572 28 573 644 645 cell_1rw
* cell instance $7194 m0 *1 179.07,38.22
X$7194 574 28 575 644 645 cell_1rw
* cell instance $7195 m0 *1 179.775,38.22
X$7195 576 28 577 644 645 cell_1rw
* cell instance $7196 m0 *1 180.48,38.22
X$7196 578 28 579 644 645 cell_1rw
* cell instance $7197 r0 *1 0.705,38.22
X$7197 67 29 68 644 645 cell_1rw
* cell instance $7198 r0 *1 0,38.22
X$7198 65 29 66 644 645 cell_1rw
* cell instance $7199 r0 *1 1.41,38.22
X$7199 69 29 70 644 645 cell_1rw
* cell instance $7200 r0 *1 2.115,38.22
X$7200 71 29 72 644 645 cell_1rw
* cell instance $7201 r0 *1 2.82,38.22
X$7201 73 29 74 644 645 cell_1rw
* cell instance $7202 r0 *1 3.525,38.22
X$7202 75 29 76 644 645 cell_1rw
* cell instance $7203 r0 *1 4.23,38.22
X$7203 77 29 78 644 645 cell_1rw
* cell instance $7204 r0 *1 4.935,38.22
X$7204 79 29 80 644 645 cell_1rw
* cell instance $7205 r0 *1 5.64,38.22
X$7205 81 29 82 644 645 cell_1rw
* cell instance $7206 r0 *1 6.345,38.22
X$7206 83 29 84 644 645 cell_1rw
* cell instance $7207 r0 *1 7.05,38.22
X$7207 85 29 86 644 645 cell_1rw
* cell instance $7208 r0 *1 7.755,38.22
X$7208 87 29 88 644 645 cell_1rw
* cell instance $7209 r0 *1 8.46,38.22
X$7209 89 29 90 644 645 cell_1rw
* cell instance $7210 r0 *1 9.165,38.22
X$7210 91 29 92 644 645 cell_1rw
* cell instance $7211 r0 *1 9.87,38.22
X$7211 93 29 94 644 645 cell_1rw
* cell instance $7212 r0 *1 10.575,38.22
X$7212 95 29 96 644 645 cell_1rw
* cell instance $7213 r0 *1 11.28,38.22
X$7213 97 29 98 644 645 cell_1rw
* cell instance $7214 r0 *1 11.985,38.22
X$7214 99 29 100 644 645 cell_1rw
* cell instance $7215 r0 *1 12.69,38.22
X$7215 101 29 102 644 645 cell_1rw
* cell instance $7216 r0 *1 13.395,38.22
X$7216 103 29 104 644 645 cell_1rw
* cell instance $7217 r0 *1 14.1,38.22
X$7217 105 29 106 644 645 cell_1rw
* cell instance $7218 r0 *1 14.805,38.22
X$7218 107 29 108 644 645 cell_1rw
* cell instance $7219 r0 *1 15.51,38.22
X$7219 109 29 110 644 645 cell_1rw
* cell instance $7220 r0 *1 16.215,38.22
X$7220 111 29 112 644 645 cell_1rw
* cell instance $7221 r0 *1 16.92,38.22
X$7221 113 29 114 644 645 cell_1rw
* cell instance $7222 r0 *1 17.625,38.22
X$7222 115 29 116 644 645 cell_1rw
* cell instance $7223 r0 *1 18.33,38.22
X$7223 117 29 118 644 645 cell_1rw
* cell instance $7224 r0 *1 19.035,38.22
X$7224 119 29 120 644 645 cell_1rw
* cell instance $7225 r0 *1 19.74,38.22
X$7225 121 29 122 644 645 cell_1rw
* cell instance $7226 r0 *1 20.445,38.22
X$7226 123 29 124 644 645 cell_1rw
* cell instance $7227 r0 *1 21.15,38.22
X$7227 125 29 126 644 645 cell_1rw
* cell instance $7228 r0 *1 21.855,38.22
X$7228 127 29 128 644 645 cell_1rw
* cell instance $7229 r0 *1 22.56,38.22
X$7229 129 29 130 644 645 cell_1rw
* cell instance $7230 r0 *1 23.265,38.22
X$7230 131 29 132 644 645 cell_1rw
* cell instance $7231 r0 *1 23.97,38.22
X$7231 133 29 134 644 645 cell_1rw
* cell instance $7232 r0 *1 24.675,38.22
X$7232 135 29 136 644 645 cell_1rw
* cell instance $7233 r0 *1 25.38,38.22
X$7233 137 29 138 644 645 cell_1rw
* cell instance $7234 r0 *1 26.085,38.22
X$7234 139 29 140 644 645 cell_1rw
* cell instance $7235 r0 *1 26.79,38.22
X$7235 141 29 142 644 645 cell_1rw
* cell instance $7236 r0 *1 27.495,38.22
X$7236 143 29 144 644 645 cell_1rw
* cell instance $7237 r0 *1 28.2,38.22
X$7237 145 29 146 644 645 cell_1rw
* cell instance $7238 r0 *1 28.905,38.22
X$7238 147 29 148 644 645 cell_1rw
* cell instance $7239 r0 *1 29.61,38.22
X$7239 149 29 150 644 645 cell_1rw
* cell instance $7240 r0 *1 30.315,38.22
X$7240 151 29 152 644 645 cell_1rw
* cell instance $7241 r0 *1 31.02,38.22
X$7241 153 29 154 644 645 cell_1rw
* cell instance $7242 r0 *1 31.725,38.22
X$7242 155 29 156 644 645 cell_1rw
* cell instance $7243 r0 *1 32.43,38.22
X$7243 157 29 158 644 645 cell_1rw
* cell instance $7244 r0 *1 33.135,38.22
X$7244 159 29 160 644 645 cell_1rw
* cell instance $7245 r0 *1 33.84,38.22
X$7245 161 29 162 644 645 cell_1rw
* cell instance $7246 r0 *1 34.545,38.22
X$7246 163 29 164 644 645 cell_1rw
* cell instance $7247 r0 *1 35.25,38.22
X$7247 165 29 166 644 645 cell_1rw
* cell instance $7248 r0 *1 35.955,38.22
X$7248 167 29 168 644 645 cell_1rw
* cell instance $7249 r0 *1 36.66,38.22
X$7249 169 29 170 644 645 cell_1rw
* cell instance $7250 r0 *1 37.365,38.22
X$7250 171 29 172 644 645 cell_1rw
* cell instance $7251 r0 *1 38.07,38.22
X$7251 173 29 174 644 645 cell_1rw
* cell instance $7252 r0 *1 38.775,38.22
X$7252 175 29 176 644 645 cell_1rw
* cell instance $7253 r0 *1 39.48,38.22
X$7253 177 29 178 644 645 cell_1rw
* cell instance $7254 r0 *1 40.185,38.22
X$7254 179 29 180 644 645 cell_1rw
* cell instance $7255 r0 *1 40.89,38.22
X$7255 181 29 182 644 645 cell_1rw
* cell instance $7256 r0 *1 41.595,38.22
X$7256 183 29 184 644 645 cell_1rw
* cell instance $7257 r0 *1 42.3,38.22
X$7257 185 29 186 644 645 cell_1rw
* cell instance $7258 r0 *1 43.005,38.22
X$7258 187 29 188 644 645 cell_1rw
* cell instance $7259 r0 *1 43.71,38.22
X$7259 189 29 190 644 645 cell_1rw
* cell instance $7260 r0 *1 44.415,38.22
X$7260 191 29 192 644 645 cell_1rw
* cell instance $7261 r0 *1 45.12,38.22
X$7261 193 29 194 644 645 cell_1rw
* cell instance $7262 r0 *1 45.825,38.22
X$7262 195 29 196 644 645 cell_1rw
* cell instance $7263 r0 *1 46.53,38.22
X$7263 197 29 198 644 645 cell_1rw
* cell instance $7264 r0 *1 47.235,38.22
X$7264 199 29 200 644 645 cell_1rw
* cell instance $7265 r0 *1 47.94,38.22
X$7265 201 29 202 644 645 cell_1rw
* cell instance $7266 r0 *1 48.645,38.22
X$7266 203 29 204 644 645 cell_1rw
* cell instance $7267 r0 *1 49.35,38.22
X$7267 205 29 206 644 645 cell_1rw
* cell instance $7268 r0 *1 50.055,38.22
X$7268 207 29 208 644 645 cell_1rw
* cell instance $7269 r0 *1 50.76,38.22
X$7269 209 29 210 644 645 cell_1rw
* cell instance $7270 r0 *1 51.465,38.22
X$7270 211 29 212 644 645 cell_1rw
* cell instance $7271 r0 *1 52.17,38.22
X$7271 213 29 214 644 645 cell_1rw
* cell instance $7272 r0 *1 52.875,38.22
X$7272 215 29 216 644 645 cell_1rw
* cell instance $7273 r0 *1 53.58,38.22
X$7273 217 29 218 644 645 cell_1rw
* cell instance $7274 r0 *1 54.285,38.22
X$7274 219 29 220 644 645 cell_1rw
* cell instance $7275 r0 *1 54.99,38.22
X$7275 221 29 222 644 645 cell_1rw
* cell instance $7276 r0 *1 55.695,38.22
X$7276 223 29 224 644 645 cell_1rw
* cell instance $7277 r0 *1 56.4,38.22
X$7277 225 29 226 644 645 cell_1rw
* cell instance $7278 r0 *1 57.105,38.22
X$7278 227 29 228 644 645 cell_1rw
* cell instance $7279 r0 *1 57.81,38.22
X$7279 229 29 230 644 645 cell_1rw
* cell instance $7280 r0 *1 58.515,38.22
X$7280 231 29 232 644 645 cell_1rw
* cell instance $7281 r0 *1 59.22,38.22
X$7281 233 29 234 644 645 cell_1rw
* cell instance $7282 r0 *1 59.925,38.22
X$7282 235 29 236 644 645 cell_1rw
* cell instance $7283 r0 *1 60.63,38.22
X$7283 237 29 238 644 645 cell_1rw
* cell instance $7284 r0 *1 61.335,38.22
X$7284 239 29 240 644 645 cell_1rw
* cell instance $7285 r0 *1 62.04,38.22
X$7285 241 29 242 644 645 cell_1rw
* cell instance $7286 r0 *1 62.745,38.22
X$7286 243 29 244 644 645 cell_1rw
* cell instance $7287 r0 *1 63.45,38.22
X$7287 245 29 246 644 645 cell_1rw
* cell instance $7288 r0 *1 64.155,38.22
X$7288 247 29 248 644 645 cell_1rw
* cell instance $7289 r0 *1 64.86,38.22
X$7289 249 29 250 644 645 cell_1rw
* cell instance $7290 r0 *1 65.565,38.22
X$7290 251 29 252 644 645 cell_1rw
* cell instance $7291 r0 *1 66.27,38.22
X$7291 253 29 254 644 645 cell_1rw
* cell instance $7292 r0 *1 66.975,38.22
X$7292 255 29 256 644 645 cell_1rw
* cell instance $7293 r0 *1 67.68,38.22
X$7293 257 29 258 644 645 cell_1rw
* cell instance $7294 r0 *1 68.385,38.22
X$7294 259 29 260 644 645 cell_1rw
* cell instance $7295 r0 *1 69.09,38.22
X$7295 261 29 262 644 645 cell_1rw
* cell instance $7296 r0 *1 69.795,38.22
X$7296 263 29 264 644 645 cell_1rw
* cell instance $7297 r0 *1 70.5,38.22
X$7297 265 29 266 644 645 cell_1rw
* cell instance $7298 r0 *1 71.205,38.22
X$7298 267 29 268 644 645 cell_1rw
* cell instance $7299 r0 *1 71.91,38.22
X$7299 269 29 270 644 645 cell_1rw
* cell instance $7300 r0 *1 72.615,38.22
X$7300 271 29 272 644 645 cell_1rw
* cell instance $7301 r0 *1 73.32,38.22
X$7301 273 29 274 644 645 cell_1rw
* cell instance $7302 r0 *1 74.025,38.22
X$7302 275 29 276 644 645 cell_1rw
* cell instance $7303 r0 *1 74.73,38.22
X$7303 277 29 278 644 645 cell_1rw
* cell instance $7304 r0 *1 75.435,38.22
X$7304 279 29 280 644 645 cell_1rw
* cell instance $7305 r0 *1 76.14,38.22
X$7305 281 29 282 644 645 cell_1rw
* cell instance $7306 r0 *1 76.845,38.22
X$7306 283 29 284 644 645 cell_1rw
* cell instance $7307 r0 *1 77.55,38.22
X$7307 285 29 286 644 645 cell_1rw
* cell instance $7308 r0 *1 78.255,38.22
X$7308 287 29 288 644 645 cell_1rw
* cell instance $7309 r0 *1 78.96,38.22
X$7309 289 29 290 644 645 cell_1rw
* cell instance $7310 r0 *1 79.665,38.22
X$7310 291 29 292 644 645 cell_1rw
* cell instance $7311 r0 *1 80.37,38.22
X$7311 293 29 294 644 645 cell_1rw
* cell instance $7312 r0 *1 81.075,38.22
X$7312 295 29 296 644 645 cell_1rw
* cell instance $7313 r0 *1 81.78,38.22
X$7313 297 29 298 644 645 cell_1rw
* cell instance $7314 r0 *1 82.485,38.22
X$7314 299 29 300 644 645 cell_1rw
* cell instance $7315 r0 *1 83.19,38.22
X$7315 301 29 302 644 645 cell_1rw
* cell instance $7316 r0 *1 83.895,38.22
X$7316 303 29 304 644 645 cell_1rw
* cell instance $7317 r0 *1 84.6,38.22
X$7317 305 29 306 644 645 cell_1rw
* cell instance $7318 r0 *1 85.305,38.22
X$7318 307 29 308 644 645 cell_1rw
* cell instance $7319 r0 *1 86.01,38.22
X$7319 309 29 310 644 645 cell_1rw
* cell instance $7320 r0 *1 86.715,38.22
X$7320 311 29 312 644 645 cell_1rw
* cell instance $7321 r0 *1 87.42,38.22
X$7321 313 29 314 644 645 cell_1rw
* cell instance $7322 r0 *1 88.125,38.22
X$7322 315 29 316 644 645 cell_1rw
* cell instance $7323 r0 *1 88.83,38.22
X$7323 317 29 318 644 645 cell_1rw
* cell instance $7324 r0 *1 89.535,38.22
X$7324 319 29 320 644 645 cell_1rw
* cell instance $7325 r0 *1 90.24,38.22
X$7325 321 29 323 644 645 cell_1rw
* cell instance $7326 r0 *1 90.945,38.22
X$7326 324 29 325 644 645 cell_1rw
* cell instance $7327 r0 *1 91.65,38.22
X$7327 326 29 327 644 645 cell_1rw
* cell instance $7328 r0 *1 92.355,38.22
X$7328 328 29 329 644 645 cell_1rw
* cell instance $7329 r0 *1 93.06,38.22
X$7329 330 29 331 644 645 cell_1rw
* cell instance $7330 r0 *1 93.765,38.22
X$7330 332 29 333 644 645 cell_1rw
* cell instance $7331 r0 *1 94.47,38.22
X$7331 334 29 335 644 645 cell_1rw
* cell instance $7332 r0 *1 95.175,38.22
X$7332 336 29 337 644 645 cell_1rw
* cell instance $7333 r0 *1 95.88,38.22
X$7333 338 29 339 644 645 cell_1rw
* cell instance $7334 r0 *1 96.585,38.22
X$7334 340 29 341 644 645 cell_1rw
* cell instance $7335 r0 *1 97.29,38.22
X$7335 342 29 343 644 645 cell_1rw
* cell instance $7336 r0 *1 97.995,38.22
X$7336 344 29 345 644 645 cell_1rw
* cell instance $7337 r0 *1 98.7,38.22
X$7337 346 29 347 644 645 cell_1rw
* cell instance $7338 r0 *1 99.405,38.22
X$7338 348 29 349 644 645 cell_1rw
* cell instance $7339 r0 *1 100.11,38.22
X$7339 350 29 351 644 645 cell_1rw
* cell instance $7340 r0 *1 100.815,38.22
X$7340 352 29 353 644 645 cell_1rw
* cell instance $7341 r0 *1 101.52,38.22
X$7341 354 29 355 644 645 cell_1rw
* cell instance $7342 r0 *1 102.225,38.22
X$7342 356 29 357 644 645 cell_1rw
* cell instance $7343 r0 *1 102.93,38.22
X$7343 358 29 359 644 645 cell_1rw
* cell instance $7344 r0 *1 103.635,38.22
X$7344 360 29 361 644 645 cell_1rw
* cell instance $7345 r0 *1 104.34,38.22
X$7345 362 29 363 644 645 cell_1rw
* cell instance $7346 r0 *1 105.045,38.22
X$7346 364 29 365 644 645 cell_1rw
* cell instance $7347 r0 *1 105.75,38.22
X$7347 366 29 367 644 645 cell_1rw
* cell instance $7348 r0 *1 106.455,38.22
X$7348 368 29 369 644 645 cell_1rw
* cell instance $7349 r0 *1 107.16,38.22
X$7349 370 29 371 644 645 cell_1rw
* cell instance $7350 r0 *1 107.865,38.22
X$7350 372 29 373 644 645 cell_1rw
* cell instance $7351 r0 *1 108.57,38.22
X$7351 374 29 375 644 645 cell_1rw
* cell instance $7352 r0 *1 109.275,38.22
X$7352 376 29 377 644 645 cell_1rw
* cell instance $7353 r0 *1 109.98,38.22
X$7353 378 29 379 644 645 cell_1rw
* cell instance $7354 r0 *1 110.685,38.22
X$7354 380 29 381 644 645 cell_1rw
* cell instance $7355 r0 *1 111.39,38.22
X$7355 382 29 383 644 645 cell_1rw
* cell instance $7356 r0 *1 112.095,38.22
X$7356 384 29 385 644 645 cell_1rw
* cell instance $7357 r0 *1 112.8,38.22
X$7357 386 29 387 644 645 cell_1rw
* cell instance $7358 r0 *1 113.505,38.22
X$7358 388 29 389 644 645 cell_1rw
* cell instance $7359 r0 *1 114.21,38.22
X$7359 390 29 391 644 645 cell_1rw
* cell instance $7360 r0 *1 114.915,38.22
X$7360 392 29 393 644 645 cell_1rw
* cell instance $7361 r0 *1 115.62,38.22
X$7361 394 29 395 644 645 cell_1rw
* cell instance $7362 r0 *1 116.325,38.22
X$7362 396 29 397 644 645 cell_1rw
* cell instance $7363 r0 *1 117.03,38.22
X$7363 398 29 399 644 645 cell_1rw
* cell instance $7364 r0 *1 117.735,38.22
X$7364 400 29 401 644 645 cell_1rw
* cell instance $7365 r0 *1 118.44,38.22
X$7365 402 29 403 644 645 cell_1rw
* cell instance $7366 r0 *1 119.145,38.22
X$7366 404 29 405 644 645 cell_1rw
* cell instance $7367 r0 *1 119.85,38.22
X$7367 406 29 407 644 645 cell_1rw
* cell instance $7368 r0 *1 120.555,38.22
X$7368 408 29 409 644 645 cell_1rw
* cell instance $7369 r0 *1 121.26,38.22
X$7369 410 29 411 644 645 cell_1rw
* cell instance $7370 r0 *1 121.965,38.22
X$7370 412 29 413 644 645 cell_1rw
* cell instance $7371 r0 *1 122.67,38.22
X$7371 414 29 415 644 645 cell_1rw
* cell instance $7372 r0 *1 123.375,38.22
X$7372 416 29 417 644 645 cell_1rw
* cell instance $7373 r0 *1 124.08,38.22
X$7373 418 29 419 644 645 cell_1rw
* cell instance $7374 r0 *1 124.785,38.22
X$7374 420 29 421 644 645 cell_1rw
* cell instance $7375 r0 *1 125.49,38.22
X$7375 422 29 423 644 645 cell_1rw
* cell instance $7376 r0 *1 126.195,38.22
X$7376 424 29 425 644 645 cell_1rw
* cell instance $7377 r0 *1 126.9,38.22
X$7377 426 29 427 644 645 cell_1rw
* cell instance $7378 r0 *1 127.605,38.22
X$7378 428 29 429 644 645 cell_1rw
* cell instance $7379 r0 *1 128.31,38.22
X$7379 430 29 431 644 645 cell_1rw
* cell instance $7380 r0 *1 129.015,38.22
X$7380 432 29 433 644 645 cell_1rw
* cell instance $7381 r0 *1 129.72,38.22
X$7381 434 29 435 644 645 cell_1rw
* cell instance $7382 r0 *1 130.425,38.22
X$7382 436 29 437 644 645 cell_1rw
* cell instance $7383 r0 *1 131.13,38.22
X$7383 438 29 439 644 645 cell_1rw
* cell instance $7384 r0 *1 131.835,38.22
X$7384 440 29 441 644 645 cell_1rw
* cell instance $7385 r0 *1 132.54,38.22
X$7385 442 29 443 644 645 cell_1rw
* cell instance $7386 r0 *1 133.245,38.22
X$7386 444 29 445 644 645 cell_1rw
* cell instance $7387 r0 *1 133.95,38.22
X$7387 446 29 447 644 645 cell_1rw
* cell instance $7388 r0 *1 134.655,38.22
X$7388 448 29 449 644 645 cell_1rw
* cell instance $7389 r0 *1 135.36,38.22
X$7389 450 29 451 644 645 cell_1rw
* cell instance $7390 r0 *1 136.065,38.22
X$7390 452 29 453 644 645 cell_1rw
* cell instance $7391 r0 *1 136.77,38.22
X$7391 454 29 455 644 645 cell_1rw
* cell instance $7392 r0 *1 137.475,38.22
X$7392 456 29 457 644 645 cell_1rw
* cell instance $7393 r0 *1 138.18,38.22
X$7393 458 29 459 644 645 cell_1rw
* cell instance $7394 r0 *1 138.885,38.22
X$7394 460 29 461 644 645 cell_1rw
* cell instance $7395 r0 *1 139.59,38.22
X$7395 462 29 463 644 645 cell_1rw
* cell instance $7396 r0 *1 140.295,38.22
X$7396 464 29 465 644 645 cell_1rw
* cell instance $7397 r0 *1 141,38.22
X$7397 466 29 467 644 645 cell_1rw
* cell instance $7398 r0 *1 141.705,38.22
X$7398 468 29 469 644 645 cell_1rw
* cell instance $7399 r0 *1 142.41,38.22
X$7399 470 29 471 644 645 cell_1rw
* cell instance $7400 r0 *1 143.115,38.22
X$7400 472 29 473 644 645 cell_1rw
* cell instance $7401 r0 *1 143.82,38.22
X$7401 474 29 475 644 645 cell_1rw
* cell instance $7402 r0 *1 144.525,38.22
X$7402 476 29 477 644 645 cell_1rw
* cell instance $7403 r0 *1 145.23,38.22
X$7403 478 29 479 644 645 cell_1rw
* cell instance $7404 r0 *1 145.935,38.22
X$7404 480 29 481 644 645 cell_1rw
* cell instance $7405 r0 *1 146.64,38.22
X$7405 482 29 483 644 645 cell_1rw
* cell instance $7406 r0 *1 147.345,38.22
X$7406 484 29 485 644 645 cell_1rw
* cell instance $7407 r0 *1 148.05,38.22
X$7407 486 29 487 644 645 cell_1rw
* cell instance $7408 r0 *1 148.755,38.22
X$7408 488 29 489 644 645 cell_1rw
* cell instance $7409 r0 *1 149.46,38.22
X$7409 490 29 491 644 645 cell_1rw
* cell instance $7410 r0 *1 150.165,38.22
X$7410 492 29 493 644 645 cell_1rw
* cell instance $7411 r0 *1 150.87,38.22
X$7411 494 29 495 644 645 cell_1rw
* cell instance $7412 r0 *1 151.575,38.22
X$7412 496 29 497 644 645 cell_1rw
* cell instance $7413 r0 *1 152.28,38.22
X$7413 498 29 499 644 645 cell_1rw
* cell instance $7414 r0 *1 152.985,38.22
X$7414 500 29 501 644 645 cell_1rw
* cell instance $7415 r0 *1 153.69,38.22
X$7415 502 29 503 644 645 cell_1rw
* cell instance $7416 r0 *1 154.395,38.22
X$7416 504 29 505 644 645 cell_1rw
* cell instance $7417 r0 *1 155.1,38.22
X$7417 506 29 507 644 645 cell_1rw
* cell instance $7418 r0 *1 155.805,38.22
X$7418 508 29 509 644 645 cell_1rw
* cell instance $7419 r0 *1 156.51,38.22
X$7419 510 29 511 644 645 cell_1rw
* cell instance $7420 r0 *1 157.215,38.22
X$7420 512 29 513 644 645 cell_1rw
* cell instance $7421 r0 *1 157.92,38.22
X$7421 514 29 515 644 645 cell_1rw
* cell instance $7422 r0 *1 158.625,38.22
X$7422 516 29 517 644 645 cell_1rw
* cell instance $7423 r0 *1 159.33,38.22
X$7423 518 29 519 644 645 cell_1rw
* cell instance $7424 r0 *1 160.035,38.22
X$7424 520 29 521 644 645 cell_1rw
* cell instance $7425 r0 *1 160.74,38.22
X$7425 522 29 523 644 645 cell_1rw
* cell instance $7426 r0 *1 161.445,38.22
X$7426 524 29 525 644 645 cell_1rw
* cell instance $7427 r0 *1 162.15,38.22
X$7427 526 29 527 644 645 cell_1rw
* cell instance $7428 r0 *1 162.855,38.22
X$7428 528 29 529 644 645 cell_1rw
* cell instance $7429 r0 *1 163.56,38.22
X$7429 530 29 531 644 645 cell_1rw
* cell instance $7430 r0 *1 164.265,38.22
X$7430 532 29 533 644 645 cell_1rw
* cell instance $7431 r0 *1 164.97,38.22
X$7431 534 29 535 644 645 cell_1rw
* cell instance $7432 r0 *1 165.675,38.22
X$7432 536 29 537 644 645 cell_1rw
* cell instance $7433 r0 *1 166.38,38.22
X$7433 538 29 539 644 645 cell_1rw
* cell instance $7434 r0 *1 167.085,38.22
X$7434 540 29 541 644 645 cell_1rw
* cell instance $7435 r0 *1 167.79,38.22
X$7435 542 29 543 644 645 cell_1rw
* cell instance $7436 r0 *1 168.495,38.22
X$7436 544 29 545 644 645 cell_1rw
* cell instance $7437 r0 *1 169.2,38.22
X$7437 546 29 547 644 645 cell_1rw
* cell instance $7438 r0 *1 169.905,38.22
X$7438 548 29 549 644 645 cell_1rw
* cell instance $7439 r0 *1 170.61,38.22
X$7439 550 29 551 644 645 cell_1rw
* cell instance $7440 r0 *1 171.315,38.22
X$7440 552 29 553 644 645 cell_1rw
* cell instance $7441 r0 *1 172.02,38.22
X$7441 554 29 555 644 645 cell_1rw
* cell instance $7442 r0 *1 172.725,38.22
X$7442 556 29 557 644 645 cell_1rw
* cell instance $7443 r0 *1 173.43,38.22
X$7443 558 29 559 644 645 cell_1rw
* cell instance $7444 r0 *1 174.135,38.22
X$7444 560 29 561 644 645 cell_1rw
* cell instance $7445 r0 *1 174.84,38.22
X$7445 562 29 563 644 645 cell_1rw
* cell instance $7446 r0 *1 175.545,38.22
X$7446 564 29 565 644 645 cell_1rw
* cell instance $7447 r0 *1 176.25,38.22
X$7447 566 29 567 644 645 cell_1rw
* cell instance $7448 r0 *1 176.955,38.22
X$7448 568 29 569 644 645 cell_1rw
* cell instance $7449 r0 *1 177.66,38.22
X$7449 570 29 571 644 645 cell_1rw
* cell instance $7450 r0 *1 178.365,38.22
X$7450 572 29 573 644 645 cell_1rw
* cell instance $7451 r0 *1 179.07,38.22
X$7451 574 29 575 644 645 cell_1rw
* cell instance $7452 r0 *1 179.775,38.22
X$7452 576 29 577 644 645 cell_1rw
* cell instance $7453 r0 *1 180.48,38.22
X$7453 578 29 579 644 645 cell_1rw
* cell instance $7454 m0 *1 0.705,40.95
X$7454 67 30 68 644 645 cell_1rw
* cell instance $7455 m0 *1 0,40.95
X$7455 65 30 66 644 645 cell_1rw
* cell instance $7456 m0 *1 1.41,40.95
X$7456 69 30 70 644 645 cell_1rw
* cell instance $7457 m0 *1 2.115,40.95
X$7457 71 30 72 644 645 cell_1rw
* cell instance $7458 m0 *1 2.82,40.95
X$7458 73 30 74 644 645 cell_1rw
* cell instance $7459 m0 *1 3.525,40.95
X$7459 75 30 76 644 645 cell_1rw
* cell instance $7460 m0 *1 4.23,40.95
X$7460 77 30 78 644 645 cell_1rw
* cell instance $7461 m0 *1 4.935,40.95
X$7461 79 30 80 644 645 cell_1rw
* cell instance $7462 m0 *1 5.64,40.95
X$7462 81 30 82 644 645 cell_1rw
* cell instance $7463 m0 *1 6.345,40.95
X$7463 83 30 84 644 645 cell_1rw
* cell instance $7464 m0 *1 7.05,40.95
X$7464 85 30 86 644 645 cell_1rw
* cell instance $7465 m0 *1 7.755,40.95
X$7465 87 30 88 644 645 cell_1rw
* cell instance $7466 m0 *1 8.46,40.95
X$7466 89 30 90 644 645 cell_1rw
* cell instance $7467 m0 *1 9.165,40.95
X$7467 91 30 92 644 645 cell_1rw
* cell instance $7468 m0 *1 9.87,40.95
X$7468 93 30 94 644 645 cell_1rw
* cell instance $7469 m0 *1 10.575,40.95
X$7469 95 30 96 644 645 cell_1rw
* cell instance $7470 m0 *1 11.28,40.95
X$7470 97 30 98 644 645 cell_1rw
* cell instance $7471 m0 *1 11.985,40.95
X$7471 99 30 100 644 645 cell_1rw
* cell instance $7472 m0 *1 12.69,40.95
X$7472 101 30 102 644 645 cell_1rw
* cell instance $7473 m0 *1 13.395,40.95
X$7473 103 30 104 644 645 cell_1rw
* cell instance $7474 m0 *1 14.1,40.95
X$7474 105 30 106 644 645 cell_1rw
* cell instance $7475 m0 *1 14.805,40.95
X$7475 107 30 108 644 645 cell_1rw
* cell instance $7476 m0 *1 15.51,40.95
X$7476 109 30 110 644 645 cell_1rw
* cell instance $7477 m0 *1 16.215,40.95
X$7477 111 30 112 644 645 cell_1rw
* cell instance $7478 m0 *1 16.92,40.95
X$7478 113 30 114 644 645 cell_1rw
* cell instance $7479 m0 *1 17.625,40.95
X$7479 115 30 116 644 645 cell_1rw
* cell instance $7480 m0 *1 18.33,40.95
X$7480 117 30 118 644 645 cell_1rw
* cell instance $7481 m0 *1 19.035,40.95
X$7481 119 30 120 644 645 cell_1rw
* cell instance $7482 m0 *1 19.74,40.95
X$7482 121 30 122 644 645 cell_1rw
* cell instance $7483 m0 *1 20.445,40.95
X$7483 123 30 124 644 645 cell_1rw
* cell instance $7484 m0 *1 21.15,40.95
X$7484 125 30 126 644 645 cell_1rw
* cell instance $7485 m0 *1 21.855,40.95
X$7485 127 30 128 644 645 cell_1rw
* cell instance $7486 m0 *1 22.56,40.95
X$7486 129 30 130 644 645 cell_1rw
* cell instance $7487 m0 *1 23.265,40.95
X$7487 131 30 132 644 645 cell_1rw
* cell instance $7488 m0 *1 23.97,40.95
X$7488 133 30 134 644 645 cell_1rw
* cell instance $7489 m0 *1 24.675,40.95
X$7489 135 30 136 644 645 cell_1rw
* cell instance $7490 m0 *1 25.38,40.95
X$7490 137 30 138 644 645 cell_1rw
* cell instance $7491 m0 *1 26.085,40.95
X$7491 139 30 140 644 645 cell_1rw
* cell instance $7492 m0 *1 26.79,40.95
X$7492 141 30 142 644 645 cell_1rw
* cell instance $7493 m0 *1 27.495,40.95
X$7493 143 30 144 644 645 cell_1rw
* cell instance $7494 m0 *1 28.2,40.95
X$7494 145 30 146 644 645 cell_1rw
* cell instance $7495 m0 *1 28.905,40.95
X$7495 147 30 148 644 645 cell_1rw
* cell instance $7496 m0 *1 29.61,40.95
X$7496 149 30 150 644 645 cell_1rw
* cell instance $7497 m0 *1 30.315,40.95
X$7497 151 30 152 644 645 cell_1rw
* cell instance $7498 m0 *1 31.02,40.95
X$7498 153 30 154 644 645 cell_1rw
* cell instance $7499 m0 *1 31.725,40.95
X$7499 155 30 156 644 645 cell_1rw
* cell instance $7500 m0 *1 32.43,40.95
X$7500 157 30 158 644 645 cell_1rw
* cell instance $7501 m0 *1 33.135,40.95
X$7501 159 30 160 644 645 cell_1rw
* cell instance $7502 m0 *1 33.84,40.95
X$7502 161 30 162 644 645 cell_1rw
* cell instance $7503 m0 *1 34.545,40.95
X$7503 163 30 164 644 645 cell_1rw
* cell instance $7504 m0 *1 35.25,40.95
X$7504 165 30 166 644 645 cell_1rw
* cell instance $7505 m0 *1 35.955,40.95
X$7505 167 30 168 644 645 cell_1rw
* cell instance $7506 m0 *1 36.66,40.95
X$7506 169 30 170 644 645 cell_1rw
* cell instance $7507 m0 *1 37.365,40.95
X$7507 171 30 172 644 645 cell_1rw
* cell instance $7508 m0 *1 38.07,40.95
X$7508 173 30 174 644 645 cell_1rw
* cell instance $7509 m0 *1 38.775,40.95
X$7509 175 30 176 644 645 cell_1rw
* cell instance $7510 m0 *1 39.48,40.95
X$7510 177 30 178 644 645 cell_1rw
* cell instance $7511 m0 *1 40.185,40.95
X$7511 179 30 180 644 645 cell_1rw
* cell instance $7512 m0 *1 40.89,40.95
X$7512 181 30 182 644 645 cell_1rw
* cell instance $7513 m0 *1 41.595,40.95
X$7513 183 30 184 644 645 cell_1rw
* cell instance $7514 m0 *1 42.3,40.95
X$7514 185 30 186 644 645 cell_1rw
* cell instance $7515 m0 *1 43.005,40.95
X$7515 187 30 188 644 645 cell_1rw
* cell instance $7516 m0 *1 43.71,40.95
X$7516 189 30 190 644 645 cell_1rw
* cell instance $7517 m0 *1 44.415,40.95
X$7517 191 30 192 644 645 cell_1rw
* cell instance $7518 m0 *1 45.12,40.95
X$7518 193 30 194 644 645 cell_1rw
* cell instance $7519 m0 *1 45.825,40.95
X$7519 195 30 196 644 645 cell_1rw
* cell instance $7520 m0 *1 46.53,40.95
X$7520 197 30 198 644 645 cell_1rw
* cell instance $7521 m0 *1 47.235,40.95
X$7521 199 30 200 644 645 cell_1rw
* cell instance $7522 m0 *1 47.94,40.95
X$7522 201 30 202 644 645 cell_1rw
* cell instance $7523 m0 *1 48.645,40.95
X$7523 203 30 204 644 645 cell_1rw
* cell instance $7524 m0 *1 49.35,40.95
X$7524 205 30 206 644 645 cell_1rw
* cell instance $7525 m0 *1 50.055,40.95
X$7525 207 30 208 644 645 cell_1rw
* cell instance $7526 m0 *1 50.76,40.95
X$7526 209 30 210 644 645 cell_1rw
* cell instance $7527 m0 *1 51.465,40.95
X$7527 211 30 212 644 645 cell_1rw
* cell instance $7528 m0 *1 52.17,40.95
X$7528 213 30 214 644 645 cell_1rw
* cell instance $7529 m0 *1 52.875,40.95
X$7529 215 30 216 644 645 cell_1rw
* cell instance $7530 m0 *1 53.58,40.95
X$7530 217 30 218 644 645 cell_1rw
* cell instance $7531 m0 *1 54.285,40.95
X$7531 219 30 220 644 645 cell_1rw
* cell instance $7532 m0 *1 54.99,40.95
X$7532 221 30 222 644 645 cell_1rw
* cell instance $7533 m0 *1 55.695,40.95
X$7533 223 30 224 644 645 cell_1rw
* cell instance $7534 m0 *1 56.4,40.95
X$7534 225 30 226 644 645 cell_1rw
* cell instance $7535 m0 *1 57.105,40.95
X$7535 227 30 228 644 645 cell_1rw
* cell instance $7536 m0 *1 57.81,40.95
X$7536 229 30 230 644 645 cell_1rw
* cell instance $7537 m0 *1 58.515,40.95
X$7537 231 30 232 644 645 cell_1rw
* cell instance $7538 m0 *1 59.22,40.95
X$7538 233 30 234 644 645 cell_1rw
* cell instance $7539 m0 *1 59.925,40.95
X$7539 235 30 236 644 645 cell_1rw
* cell instance $7540 m0 *1 60.63,40.95
X$7540 237 30 238 644 645 cell_1rw
* cell instance $7541 m0 *1 61.335,40.95
X$7541 239 30 240 644 645 cell_1rw
* cell instance $7542 m0 *1 62.04,40.95
X$7542 241 30 242 644 645 cell_1rw
* cell instance $7543 m0 *1 62.745,40.95
X$7543 243 30 244 644 645 cell_1rw
* cell instance $7544 m0 *1 63.45,40.95
X$7544 245 30 246 644 645 cell_1rw
* cell instance $7545 m0 *1 64.155,40.95
X$7545 247 30 248 644 645 cell_1rw
* cell instance $7546 m0 *1 64.86,40.95
X$7546 249 30 250 644 645 cell_1rw
* cell instance $7547 m0 *1 65.565,40.95
X$7547 251 30 252 644 645 cell_1rw
* cell instance $7548 m0 *1 66.27,40.95
X$7548 253 30 254 644 645 cell_1rw
* cell instance $7549 m0 *1 66.975,40.95
X$7549 255 30 256 644 645 cell_1rw
* cell instance $7550 m0 *1 67.68,40.95
X$7550 257 30 258 644 645 cell_1rw
* cell instance $7551 m0 *1 68.385,40.95
X$7551 259 30 260 644 645 cell_1rw
* cell instance $7552 m0 *1 69.09,40.95
X$7552 261 30 262 644 645 cell_1rw
* cell instance $7553 m0 *1 69.795,40.95
X$7553 263 30 264 644 645 cell_1rw
* cell instance $7554 m0 *1 70.5,40.95
X$7554 265 30 266 644 645 cell_1rw
* cell instance $7555 m0 *1 71.205,40.95
X$7555 267 30 268 644 645 cell_1rw
* cell instance $7556 m0 *1 71.91,40.95
X$7556 269 30 270 644 645 cell_1rw
* cell instance $7557 m0 *1 72.615,40.95
X$7557 271 30 272 644 645 cell_1rw
* cell instance $7558 m0 *1 73.32,40.95
X$7558 273 30 274 644 645 cell_1rw
* cell instance $7559 m0 *1 74.025,40.95
X$7559 275 30 276 644 645 cell_1rw
* cell instance $7560 m0 *1 74.73,40.95
X$7560 277 30 278 644 645 cell_1rw
* cell instance $7561 m0 *1 75.435,40.95
X$7561 279 30 280 644 645 cell_1rw
* cell instance $7562 m0 *1 76.14,40.95
X$7562 281 30 282 644 645 cell_1rw
* cell instance $7563 m0 *1 76.845,40.95
X$7563 283 30 284 644 645 cell_1rw
* cell instance $7564 m0 *1 77.55,40.95
X$7564 285 30 286 644 645 cell_1rw
* cell instance $7565 m0 *1 78.255,40.95
X$7565 287 30 288 644 645 cell_1rw
* cell instance $7566 m0 *1 78.96,40.95
X$7566 289 30 290 644 645 cell_1rw
* cell instance $7567 m0 *1 79.665,40.95
X$7567 291 30 292 644 645 cell_1rw
* cell instance $7568 m0 *1 80.37,40.95
X$7568 293 30 294 644 645 cell_1rw
* cell instance $7569 m0 *1 81.075,40.95
X$7569 295 30 296 644 645 cell_1rw
* cell instance $7570 m0 *1 81.78,40.95
X$7570 297 30 298 644 645 cell_1rw
* cell instance $7571 m0 *1 82.485,40.95
X$7571 299 30 300 644 645 cell_1rw
* cell instance $7572 m0 *1 83.19,40.95
X$7572 301 30 302 644 645 cell_1rw
* cell instance $7573 m0 *1 83.895,40.95
X$7573 303 30 304 644 645 cell_1rw
* cell instance $7574 m0 *1 84.6,40.95
X$7574 305 30 306 644 645 cell_1rw
* cell instance $7575 m0 *1 85.305,40.95
X$7575 307 30 308 644 645 cell_1rw
* cell instance $7576 m0 *1 86.01,40.95
X$7576 309 30 310 644 645 cell_1rw
* cell instance $7577 m0 *1 86.715,40.95
X$7577 311 30 312 644 645 cell_1rw
* cell instance $7578 m0 *1 87.42,40.95
X$7578 313 30 314 644 645 cell_1rw
* cell instance $7579 m0 *1 88.125,40.95
X$7579 315 30 316 644 645 cell_1rw
* cell instance $7580 m0 *1 88.83,40.95
X$7580 317 30 318 644 645 cell_1rw
* cell instance $7581 m0 *1 89.535,40.95
X$7581 319 30 320 644 645 cell_1rw
* cell instance $7582 m0 *1 90.24,40.95
X$7582 321 30 323 644 645 cell_1rw
* cell instance $7583 m0 *1 90.945,40.95
X$7583 324 30 325 644 645 cell_1rw
* cell instance $7584 m0 *1 91.65,40.95
X$7584 326 30 327 644 645 cell_1rw
* cell instance $7585 m0 *1 92.355,40.95
X$7585 328 30 329 644 645 cell_1rw
* cell instance $7586 m0 *1 93.06,40.95
X$7586 330 30 331 644 645 cell_1rw
* cell instance $7587 m0 *1 93.765,40.95
X$7587 332 30 333 644 645 cell_1rw
* cell instance $7588 m0 *1 94.47,40.95
X$7588 334 30 335 644 645 cell_1rw
* cell instance $7589 m0 *1 95.175,40.95
X$7589 336 30 337 644 645 cell_1rw
* cell instance $7590 m0 *1 95.88,40.95
X$7590 338 30 339 644 645 cell_1rw
* cell instance $7591 m0 *1 96.585,40.95
X$7591 340 30 341 644 645 cell_1rw
* cell instance $7592 m0 *1 97.29,40.95
X$7592 342 30 343 644 645 cell_1rw
* cell instance $7593 m0 *1 97.995,40.95
X$7593 344 30 345 644 645 cell_1rw
* cell instance $7594 m0 *1 98.7,40.95
X$7594 346 30 347 644 645 cell_1rw
* cell instance $7595 m0 *1 99.405,40.95
X$7595 348 30 349 644 645 cell_1rw
* cell instance $7596 m0 *1 100.11,40.95
X$7596 350 30 351 644 645 cell_1rw
* cell instance $7597 m0 *1 100.815,40.95
X$7597 352 30 353 644 645 cell_1rw
* cell instance $7598 m0 *1 101.52,40.95
X$7598 354 30 355 644 645 cell_1rw
* cell instance $7599 m0 *1 102.225,40.95
X$7599 356 30 357 644 645 cell_1rw
* cell instance $7600 m0 *1 102.93,40.95
X$7600 358 30 359 644 645 cell_1rw
* cell instance $7601 m0 *1 103.635,40.95
X$7601 360 30 361 644 645 cell_1rw
* cell instance $7602 m0 *1 104.34,40.95
X$7602 362 30 363 644 645 cell_1rw
* cell instance $7603 m0 *1 105.045,40.95
X$7603 364 30 365 644 645 cell_1rw
* cell instance $7604 m0 *1 105.75,40.95
X$7604 366 30 367 644 645 cell_1rw
* cell instance $7605 m0 *1 106.455,40.95
X$7605 368 30 369 644 645 cell_1rw
* cell instance $7606 m0 *1 107.16,40.95
X$7606 370 30 371 644 645 cell_1rw
* cell instance $7607 m0 *1 107.865,40.95
X$7607 372 30 373 644 645 cell_1rw
* cell instance $7608 m0 *1 108.57,40.95
X$7608 374 30 375 644 645 cell_1rw
* cell instance $7609 m0 *1 109.275,40.95
X$7609 376 30 377 644 645 cell_1rw
* cell instance $7610 m0 *1 109.98,40.95
X$7610 378 30 379 644 645 cell_1rw
* cell instance $7611 m0 *1 110.685,40.95
X$7611 380 30 381 644 645 cell_1rw
* cell instance $7612 m0 *1 111.39,40.95
X$7612 382 30 383 644 645 cell_1rw
* cell instance $7613 m0 *1 112.095,40.95
X$7613 384 30 385 644 645 cell_1rw
* cell instance $7614 m0 *1 112.8,40.95
X$7614 386 30 387 644 645 cell_1rw
* cell instance $7615 m0 *1 113.505,40.95
X$7615 388 30 389 644 645 cell_1rw
* cell instance $7616 m0 *1 114.21,40.95
X$7616 390 30 391 644 645 cell_1rw
* cell instance $7617 m0 *1 114.915,40.95
X$7617 392 30 393 644 645 cell_1rw
* cell instance $7618 m0 *1 115.62,40.95
X$7618 394 30 395 644 645 cell_1rw
* cell instance $7619 m0 *1 116.325,40.95
X$7619 396 30 397 644 645 cell_1rw
* cell instance $7620 m0 *1 117.03,40.95
X$7620 398 30 399 644 645 cell_1rw
* cell instance $7621 m0 *1 117.735,40.95
X$7621 400 30 401 644 645 cell_1rw
* cell instance $7622 m0 *1 118.44,40.95
X$7622 402 30 403 644 645 cell_1rw
* cell instance $7623 m0 *1 119.145,40.95
X$7623 404 30 405 644 645 cell_1rw
* cell instance $7624 m0 *1 119.85,40.95
X$7624 406 30 407 644 645 cell_1rw
* cell instance $7625 m0 *1 120.555,40.95
X$7625 408 30 409 644 645 cell_1rw
* cell instance $7626 m0 *1 121.26,40.95
X$7626 410 30 411 644 645 cell_1rw
* cell instance $7627 m0 *1 121.965,40.95
X$7627 412 30 413 644 645 cell_1rw
* cell instance $7628 m0 *1 122.67,40.95
X$7628 414 30 415 644 645 cell_1rw
* cell instance $7629 m0 *1 123.375,40.95
X$7629 416 30 417 644 645 cell_1rw
* cell instance $7630 m0 *1 124.08,40.95
X$7630 418 30 419 644 645 cell_1rw
* cell instance $7631 m0 *1 124.785,40.95
X$7631 420 30 421 644 645 cell_1rw
* cell instance $7632 m0 *1 125.49,40.95
X$7632 422 30 423 644 645 cell_1rw
* cell instance $7633 m0 *1 126.195,40.95
X$7633 424 30 425 644 645 cell_1rw
* cell instance $7634 m0 *1 126.9,40.95
X$7634 426 30 427 644 645 cell_1rw
* cell instance $7635 m0 *1 127.605,40.95
X$7635 428 30 429 644 645 cell_1rw
* cell instance $7636 m0 *1 128.31,40.95
X$7636 430 30 431 644 645 cell_1rw
* cell instance $7637 m0 *1 129.015,40.95
X$7637 432 30 433 644 645 cell_1rw
* cell instance $7638 m0 *1 129.72,40.95
X$7638 434 30 435 644 645 cell_1rw
* cell instance $7639 m0 *1 130.425,40.95
X$7639 436 30 437 644 645 cell_1rw
* cell instance $7640 m0 *1 131.13,40.95
X$7640 438 30 439 644 645 cell_1rw
* cell instance $7641 m0 *1 131.835,40.95
X$7641 440 30 441 644 645 cell_1rw
* cell instance $7642 m0 *1 132.54,40.95
X$7642 442 30 443 644 645 cell_1rw
* cell instance $7643 m0 *1 133.245,40.95
X$7643 444 30 445 644 645 cell_1rw
* cell instance $7644 m0 *1 133.95,40.95
X$7644 446 30 447 644 645 cell_1rw
* cell instance $7645 m0 *1 134.655,40.95
X$7645 448 30 449 644 645 cell_1rw
* cell instance $7646 m0 *1 135.36,40.95
X$7646 450 30 451 644 645 cell_1rw
* cell instance $7647 m0 *1 136.065,40.95
X$7647 452 30 453 644 645 cell_1rw
* cell instance $7648 m0 *1 136.77,40.95
X$7648 454 30 455 644 645 cell_1rw
* cell instance $7649 m0 *1 137.475,40.95
X$7649 456 30 457 644 645 cell_1rw
* cell instance $7650 m0 *1 138.18,40.95
X$7650 458 30 459 644 645 cell_1rw
* cell instance $7651 m0 *1 138.885,40.95
X$7651 460 30 461 644 645 cell_1rw
* cell instance $7652 m0 *1 139.59,40.95
X$7652 462 30 463 644 645 cell_1rw
* cell instance $7653 m0 *1 140.295,40.95
X$7653 464 30 465 644 645 cell_1rw
* cell instance $7654 m0 *1 141,40.95
X$7654 466 30 467 644 645 cell_1rw
* cell instance $7655 m0 *1 141.705,40.95
X$7655 468 30 469 644 645 cell_1rw
* cell instance $7656 m0 *1 142.41,40.95
X$7656 470 30 471 644 645 cell_1rw
* cell instance $7657 m0 *1 143.115,40.95
X$7657 472 30 473 644 645 cell_1rw
* cell instance $7658 m0 *1 143.82,40.95
X$7658 474 30 475 644 645 cell_1rw
* cell instance $7659 m0 *1 144.525,40.95
X$7659 476 30 477 644 645 cell_1rw
* cell instance $7660 m0 *1 145.23,40.95
X$7660 478 30 479 644 645 cell_1rw
* cell instance $7661 m0 *1 145.935,40.95
X$7661 480 30 481 644 645 cell_1rw
* cell instance $7662 m0 *1 146.64,40.95
X$7662 482 30 483 644 645 cell_1rw
* cell instance $7663 m0 *1 147.345,40.95
X$7663 484 30 485 644 645 cell_1rw
* cell instance $7664 m0 *1 148.05,40.95
X$7664 486 30 487 644 645 cell_1rw
* cell instance $7665 m0 *1 148.755,40.95
X$7665 488 30 489 644 645 cell_1rw
* cell instance $7666 m0 *1 149.46,40.95
X$7666 490 30 491 644 645 cell_1rw
* cell instance $7667 m0 *1 150.165,40.95
X$7667 492 30 493 644 645 cell_1rw
* cell instance $7668 m0 *1 150.87,40.95
X$7668 494 30 495 644 645 cell_1rw
* cell instance $7669 m0 *1 151.575,40.95
X$7669 496 30 497 644 645 cell_1rw
* cell instance $7670 m0 *1 152.28,40.95
X$7670 498 30 499 644 645 cell_1rw
* cell instance $7671 m0 *1 152.985,40.95
X$7671 500 30 501 644 645 cell_1rw
* cell instance $7672 m0 *1 153.69,40.95
X$7672 502 30 503 644 645 cell_1rw
* cell instance $7673 m0 *1 154.395,40.95
X$7673 504 30 505 644 645 cell_1rw
* cell instance $7674 m0 *1 155.1,40.95
X$7674 506 30 507 644 645 cell_1rw
* cell instance $7675 m0 *1 155.805,40.95
X$7675 508 30 509 644 645 cell_1rw
* cell instance $7676 m0 *1 156.51,40.95
X$7676 510 30 511 644 645 cell_1rw
* cell instance $7677 m0 *1 157.215,40.95
X$7677 512 30 513 644 645 cell_1rw
* cell instance $7678 m0 *1 157.92,40.95
X$7678 514 30 515 644 645 cell_1rw
* cell instance $7679 m0 *1 158.625,40.95
X$7679 516 30 517 644 645 cell_1rw
* cell instance $7680 m0 *1 159.33,40.95
X$7680 518 30 519 644 645 cell_1rw
* cell instance $7681 m0 *1 160.035,40.95
X$7681 520 30 521 644 645 cell_1rw
* cell instance $7682 m0 *1 160.74,40.95
X$7682 522 30 523 644 645 cell_1rw
* cell instance $7683 m0 *1 161.445,40.95
X$7683 524 30 525 644 645 cell_1rw
* cell instance $7684 m0 *1 162.15,40.95
X$7684 526 30 527 644 645 cell_1rw
* cell instance $7685 m0 *1 162.855,40.95
X$7685 528 30 529 644 645 cell_1rw
* cell instance $7686 m0 *1 163.56,40.95
X$7686 530 30 531 644 645 cell_1rw
* cell instance $7687 m0 *1 164.265,40.95
X$7687 532 30 533 644 645 cell_1rw
* cell instance $7688 m0 *1 164.97,40.95
X$7688 534 30 535 644 645 cell_1rw
* cell instance $7689 m0 *1 165.675,40.95
X$7689 536 30 537 644 645 cell_1rw
* cell instance $7690 m0 *1 166.38,40.95
X$7690 538 30 539 644 645 cell_1rw
* cell instance $7691 m0 *1 167.085,40.95
X$7691 540 30 541 644 645 cell_1rw
* cell instance $7692 m0 *1 167.79,40.95
X$7692 542 30 543 644 645 cell_1rw
* cell instance $7693 m0 *1 168.495,40.95
X$7693 544 30 545 644 645 cell_1rw
* cell instance $7694 m0 *1 169.2,40.95
X$7694 546 30 547 644 645 cell_1rw
* cell instance $7695 m0 *1 169.905,40.95
X$7695 548 30 549 644 645 cell_1rw
* cell instance $7696 m0 *1 170.61,40.95
X$7696 550 30 551 644 645 cell_1rw
* cell instance $7697 m0 *1 171.315,40.95
X$7697 552 30 553 644 645 cell_1rw
* cell instance $7698 m0 *1 172.02,40.95
X$7698 554 30 555 644 645 cell_1rw
* cell instance $7699 m0 *1 172.725,40.95
X$7699 556 30 557 644 645 cell_1rw
* cell instance $7700 m0 *1 173.43,40.95
X$7700 558 30 559 644 645 cell_1rw
* cell instance $7701 m0 *1 174.135,40.95
X$7701 560 30 561 644 645 cell_1rw
* cell instance $7702 m0 *1 174.84,40.95
X$7702 562 30 563 644 645 cell_1rw
* cell instance $7703 m0 *1 175.545,40.95
X$7703 564 30 565 644 645 cell_1rw
* cell instance $7704 m0 *1 176.25,40.95
X$7704 566 30 567 644 645 cell_1rw
* cell instance $7705 m0 *1 176.955,40.95
X$7705 568 30 569 644 645 cell_1rw
* cell instance $7706 m0 *1 177.66,40.95
X$7706 570 30 571 644 645 cell_1rw
* cell instance $7707 m0 *1 178.365,40.95
X$7707 572 30 573 644 645 cell_1rw
* cell instance $7708 m0 *1 179.07,40.95
X$7708 574 30 575 644 645 cell_1rw
* cell instance $7709 m0 *1 179.775,40.95
X$7709 576 30 577 644 645 cell_1rw
* cell instance $7710 m0 *1 180.48,40.95
X$7710 578 30 579 644 645 cell_1rw
* cell instance $7711 r0 *1 0.705,40.95
X$7711 67 31 68 644 645 cell_1rw
* cell instance $7712 r0 *1 0,40.95
X$7712 65 31 66 644 645 cell_1rw
* cell instance $7713 r0 *1 1.41,40.95
X$7713 69 31 70 644 645 cell_1rw
* cell instance $7714 r0 *1 2.115,40.95
X$7714 71 31 72 644 645 cell_1rw
* cell instance $7715 r0 *1 2.82,40.95
X$7715 73 31 74 644 645 cell_1rw
* cell instance $7716 r0 *1 3.525,40.95
X$7716 75 31 76 644 645 cell_1rw
* cell instance $7717 r0 *1 4.23,40.95
X$7717 77 31 78 644 645 cell_1rw
* cell instance $7718 r0 *1 4.935,40.95
X$7718 79 31 80 644 645 cell_1rw
* cell instance $7719 r0 *1 5.64,40.95
X$7719 81 31 82 644 645 cell_1rw
* cell instance $7720 r0 *1 6.345,40.95
X$7720 83 31 84 644 645 cell_1rw
* cell instance $7721 r0 *1 7.05,40.95
X$7721 85 31 86 644 645 cell_1rw
* cell instance $7722 r0 *1 7.755,40.95
X$7722 87 31 88 644 645 cell_1rw
* cell instance $7723 r0 *1 8.46,40.95
X$7723 89 31 90 644 645 cell_1rw
* cell instance $7724 r0 *1 9.165,40.95
X$7724 91 31 92 644 645 cell_1rw
* cell instance $7725 r0 *1 9.87,40.95
X$7725 93 31 94 644 645 cell_1rw
* cell instance $7726 r0 *1 10.575,40.95
X$7726 95 31 96 644 645 cell_1rw
* cell instance $7727 r0 *1 11.28,40.95
X$7727 97 31 98 644 645 cell_1rw
* cell instance $7728 r0 *1 11.985,40.95
X$7728 99 31 100 644 645 cell_1rw
* cell instance $7729 r0 *1 12.69,40.95
X$7729 101 31 102 644 645 cell_1rw
* cell instance $7730 r0 *1 13.395,40.95
X$7730 103 31 104 644 645 cell_1rw
* cell instance $7731 r0 *1 14.1,40.95
X$7731 105 31 106 644 645 cell_1rw
* cell instance $7732 r0 *1 14.805,40.95
X$7732 107 31 108 644 645 cell_1rw
* cell instance $7733 r0 *1 15.51,40.95
X$7733 109 31 110 644 645 cell_1rw
* cell instance $7734 r0 *1 16.215,40.95
X$7734 111 31 112 644 645 cell_1rw
* cell instance $7735 r0 *1 16.92,40.95
X$7735 113 31 114 644 645 cell_1rw
* cell instance $7736 r0 *1 17.625,40.95
X$7736 115 31 116 644 645 cell_1rw
* cell instance $7737 r0 *1 18.33,40.95
X$7737 117 31 118 644 645 cell_1rw
* cell instance $7738 r0 *1 19.035,40.95
X$7738 119 31 120 644 645 cell_1rw
* cell instance $7739 r0 *1 19.74,40.95
X$7739 121 31 122 644 645 cell_1rw
* cell instance $7740 r0 *1 20.445,40.95
X$7740 123 31 124 644 645 cell_1rw
* cell instance $7741 r0 *1 21.15,40.95
X$7741 125 31 126 644 645 cell_1rw
* cell instance $7742 r0 *1 21.855,40.95
X$7742 127 31 128 644 645 cell_1rw
* cell instance $7743 r0 *1 22.56,40.95
X$7743 129 31 130 644 645 cell_1rw
* cell instance $7744 r0 *1 23.265,40.95
X$7744 131 31 132 644 645 cell_1rw
* cell instance $7745 r0 *1 23.97,40.95
X$7745 133 31 134 644 645 cell_1rw
* cell instance $7746 r0 *1 24.675,40.95
X$7746 135 31 136 644 645 cell_1rw
* cell instance $7747 r0 *1 25.38,40.95
X$7747 137 31 138 644 645 cell_1rw
* cell instance $7748 r0 *1 26.085,40.95
X$7748 139 31 140 644 645 cell_1rw
* cell instance $7749 r0 *1 26.79,40.95
X$7749 141 31 142 644 645 cell_1rw
* cell instance $7750 r0 *1 27.495,40.95
X$7750 143 31 144 644 645 cell_1rw
* cell instance $7751 r0 *1 28.2,40.95
X$7751 145 31 146 644 645 cell_1rw
* cell instance $7752 r0 *1 28.905,40.95
X$7752 147 31 148 644 645 cell_1rw
* cell instance $7753 r0 *1 29.61,40.95
X$7753 149 31 150 644 645 cell_1rw
* cell instance $7754 r0 *1 30.315,40.95
X$7754 151 31 152 644 645 cell_1rw
* cell instance $7755 r0 *1 31.02,40.95
X$7755 153 31 154 644 645 cell_1rw
* cell instance $7756 r0 *1 31.725,40.95
X$7756 155 31 156 644 645 cell_1rw
* cell instance $7757 r0 *1 32.43,40.95
X$7757 157 31 158 644 645 cell_1rw
* cell instance $7758 r0 *1 33.135,40.95
X$7758 159 31 160 644 645 cell_1rw
* cell instance $7759 r0 *1 33.84,40.95
X$7759 161 31 162 644 645 cell_1rw
* cell instance $7760 r0 *1 34.545,40.95
X$7760 163 31 164 644 645 cell_1rw
* cell instance $7761 r0 *1 35.25,40.95
X$7761 165 31 166 644 645 cell_1rw
* cell instance $7762 r0 *1 35.955,40.95
X$7762 167 31 168 644 645 cell_1rw
* cell instance $7763 r0 *1 36.66,40.95
X$7763 169 31 170 644 645 cell_1rw
* cell instance $7764 r0 *1 37.365,40.95
X$7764 171 31 172 644 645 cell_1rw
* cell instance $7765 r0 *1 38.07,40.95
X$7765 173 31 174 644 645 cell_1rw
* cell instance $7766 r0 *1 38.775,40.95
X$7766 175 31 176 644 645 cell_1rw
* cell instance $7767 r0 *1 39.48,40.95
X$7767 177 31 178 644 645 cell_1rw
* cell instance $7768 r0 *1 40.185,40.95
X$7768 179 31 180 644 645 cell_1rw
* cell instance $7769 r0 *1 40.89,40.95
X$7769 181 31 182 644 645 cell_1rw
* cell instance $7770 r0 *1 41.595,40.95
X$7770 183 31 184 644 645 cell_1rw
* cell instance $7771 r0 *1 42.3,40.95
X$7771 185 31 186 644 645 cell_1rw
* cell instance $7772 r0 *1 43.005,40.95
X$7772 187 31 188 644 645 cell_1rw
* cell instance $7773 r0 *1 43.71,40.95
X$7773 189 31 190 644 645 cell_1rw
* cell instance $7774 r0 *1 44.415,40.95
X$7774 191 31 192 644 645 cell_1rw
* cell instance $7775 r0 *1 45.12,40.95
X$7775 193 31 194 644 645 cell_1rw
* cell instance $7776 r0 *1 45.825,40.95
X$7776 195 31 196 644 645 cell_1rw
* cell instance $7777 r0 *1 46.53,40.95
X$7777 197 31 198 644 645 cell_1rw
* cell instance $7778 r0 *1 47.235,40.95
X$7778 199 31 200 644 645 cell_1rw
* cell instance $7779 r0 *1 47.94,40.95
X$7779 201 31 202 644 645 cell_1rw
* cell instance $7780 r0 *1 48.645,40.95
X$7780 203 31 204 644 645 cell_1rw
* cell instance $7781 r0 *1 49.35,40.95
X$7781 205 31 206 644 645 cell_1rw
* cell instance $7782 r0 *1 50.055,40.95
X$7782 207 31 208 644 645 cell_1rw
* cell instance $7783 r0 *1 50.76,40.95
X$7783 209 31 210 644 645 cell_1rw
* cell instance $7784 r0 *1 51.465,40.95
X$7784 211 31 212 644 645 cell_1rw
* cell instance $7785 r0 *1 52.17,40.95
X$7785 213 31 214 644 645 cell_1rw
* cell instance $7786 r0 *1 52.875,40.95
X$7786 215 31 216 644 645 cell_1rw
* cell instance $7787 r0 *1 53.58,40.95
X$7787 217 31 218 644 645 cell_1rw
* cell instance $7788 r0 *1 54.285,40.95
X$7788 219 31 220 644 645 cell_1rw
* cell instance $7789 r0 *1 54.99,40.95
X$7789 221 31 222 644 645 cell_1rw
* cell instance $7790 r0 *1 55.695,40.95
X$7790 223 31 224 644 645 cell_1rw
* cell instance $7791 r0 *1 56.4,40.95
X$7791 225 31 226 644 645 cell_1rw
* cell instance $7792 r0 *1 57.105,40.95
X$7792 227 31 228 644 645 cell_1rw
* cell instance $7793 r0 *1 57.81,40.95
X$7793 229 31 230 644 645 cell_1rw
* cell instance $7794 r0 *1 58.515,40.95
X$7794 231 31 232 644 645 cell_1rw
* cell instance $7795 r0 *1 59.22,40.95
X$7795 233 31 234 644 645 cell_1rw
* cell instance $7796 r0 *1 59.925,40.95
X$7796 235 31 236 644 645 cell_1rw
* cell instance $7797 r0 *1 60.63,40.95
X$7797 237 31 238 644 645 cell_1rw
* cell instance $7798 r0 *1 61.335,40.95
X$7798 239 31 240 644 645 cell_1rw
* cell instance $7799 r0 *1 62.04,40.95
X$7799 241 31 242 644 645 cell_1rw
* cell instance $7800 r0 *1 62.745,40.95
X$7800 243 31 244 644 645 cell_1rw
* cell instance $7801 r0 *1 63.45,40.95
X$7801 245 31 246 644 645 cell_1rw
* cell instance $7802 r0 *1 64.155,40.95
X$7802 247 31 248 644 645 cell_1rw
* cell instance $7803 r0 *1 64.86,40.95
X$7803 249 31 250 644 645 cell_1rw
* cell instance $7804 r0 *1 65.565,40.95
X$7804 251 31 252 644 645 cell_1rw
* cell instance $7805 r0 *1 66.27,40.95
X$7805 253 31 254 644 645 cell_1rw
* cell instance $7806 r0 *1 66.975,40.95
X$7806 255 31 256 644 645 cell_1rw
* cell instance $7807 r0 *1 67.68,40.95
X$7807 257 31 258 644 645 cell_1rw
* cell instance $7808 r0 *1 68.385,40.95
X$7808 259 31 260 644 645 cell_1rw
* cell instance $7809 r0 *1 69.09,40.95
X$7809 261 31 262 644 645 cell_1rw
* cell instance $7810 r0 *1 69.795,40.95
X$7810 263 31 264 644 645 cell_1rw
* cell instance $7811 r0 *1 70.5,40.95
X$7811 265 31 266 644 645 cell_1rw
* cell instance $7812 r0 *1 71.205,40.95
X$7812 267 31 268 644 645 cell_1rw
* cell instance $7813 r0 *1 71.91,40.95
X$7813 269 31 270 644 645 cell_1rw
* cell instance $7814 r0 *1 72.615,40.95
X$7814 271 31 272 644 645 cell_1rw
* cell instance $7815 r0 *1 73.32,40.95
X$7815 273 31 274 644 645 cell_1rw
* cell instance $7816 r0 *1 74.025,40.95
X$7816 275 31 276 644 645 cell_1rw
* cell instance $7817 r0 *1 74.73,40.95
X$7817 277 31 278 644 645 cell_1rw
* cell instance $7818 r0 *1 75.435,40.95
X$7818 279 31 280 644 645 cell_1rw
* cell instance $7819 r0 *1 76.14,40.95
X$7819 281 31 282 644 645 cell_1rw
* cell instance $7820 r0 *1 76.845,40.95
X$7820 283 31 284 644 645 cell_1rw
* cell instance $7821 r0 *1 77.55,40.95
X$7821 285 31 286 644 645 cell_1rw
* cell instance $7822 r0 *1 78.255,40.95
X$7822 287 31 288 644 645 cell_1rw
* cell instance $7823 r0 *1 78.96,40.95
X$7823 289 31 290 644 645 cell_1rw
* cell instance $7824 r0 *1 79.665,40.95
X$7824 291 31 292 644 645 cell_1rw
* cell instance $7825 r0 *1 80.37,40.95
X$7825 293 31 294 644 645 cell_1rw
* cell instance $7826 r0 *1 81.075,40.95
X$7826 295 31 296 644 645 cell_1rw
* cell instance $7827 r0 *1 81.78,40.95
X$7827 297 31 298 644 645 cell_1rw
* cell instance $7828 r0 *1 82.485,40.95
X$7828 299 31 300 644 645 cell_1rw
* cell instance $7829 r0 *1 83.19,40.95
X$7829 301 31 302 644 645 cell_1rw
* cell instance $7830 r0 *1 83.895,40.95
X$7830 303 31 304 644 645 cell_1rw
* cell instance $7831 r0 *1 84.6,40.95
X$7831 305 31 306 644 645 cell_1rw
* cell instance $7832 r0 *1 85.305,40.95
X$7832 307 31 308 644 645 cell_1rw
* cell instance $7833 r0 *1 86.01,40.95
X$7833 309 31 310 644 645 cell_1rw
* cell instance $7834 r0 *1 86.715,40.95
X$7834 311 31 312 644 645 cell_1rw
* cell instance $7835 r0 *1 87.42,40.95
X$7835 313 31 314 644 645 cell_1rw
* cell instance $7836 r0 *1 88.125,40.95
X$7836 315 31 316 644 645 cell_1rw
* cell instance $7837 r0 *1 88.83,40.95
X$7837 317 31 318 644 645 cell_1rw
* cell instance $7838 r0 *1 89.535,40.95
X$7838 319 31 320 644 645 cell_1rw
* cell instance $7839 r0 *1 90.24,40.95
X$7839 321 31 323 644 645 cell_1rw
* cell instance $7840 r0 *1 90.945,40.95
X$7840 324 31 325 644 645 cell_1rw
* cell instance $7841 r0 *1 91.65,40.95
X$7841 326 31 327 644 645 cell_1rw
* cell instance $7842 r0 *1 92.355,40.95
X$7842 328 31 329 644 645 cell_1rw
* cell instance $7843 r0 *1 93.06,40.95
X$7843 330 31 331 644 645 cell_1rw
* cell instance $7844 r0 *1 93.765,40.95
X$7844 332 31 333 644 645 cell_1rw
* cell instance $7845 r0 *1 94.47,40.95
X$7845 334 31 335 644 645 cell_1rw
* cell instance $7846 r0 *1 95.175,40.95
X$7846 336 31 337 644 645 cell_1rw
* cell instance $7847 r0 *1 95.88,40.95
X$7847 338 31 339 644 645 cell_1rw
* cell instance $7848 r0 *1 96.585,40.95
X$7848 340 31 341 644 645 cell_1rw
* cell instance $7849 r0 *1 97.29,40.95
X$7849 342 31 343 644 645 cell_1rw
* cell instance $7850 r0 *1 97.995,40.95
X$7850 344 31 345 644 645 cell_1rw
* cell instance $7851 r0 *1 98.7,40.95
X$7851 346 31 347 644 645 cell_1rw
* cell instance $7852 r0 *1 99.405,40.95
X$7852 348 31 349 644 645 cell_1rw
* cell instance $7853 r0 *1 100.11,40.95
X$7853 350 31 351 644 645 cell_1rw
* cell instance $7854 r0 *1 100.815,40.95
X$7854 352 31 353 644 645 cell_1rw
* cell instance $7855 r0 *1 101.52,40.95
X$7855 354 31 355 644 645 cell_1rw
* cell instance $7856 r0 *1 102.225,40.95
X$7856 356 31 357 644 645 cell_1rw
* cell instance $7857 r0 *1 102.93,40.95
X$7857 358 31 359 644 645 cell_1rw
* cell instance $7858 r0 *1 103.635,40.95
X$7858 360 31 361 644 645 cell_1rw
* cell instance $7859 r0 *1 104.34,40.95
X$7859 362 31 363 644 645 cell_1rw
* cell instance $7860 r0 *1 105.045,40.95
X$7860 364 31 365 644 645 cell_1rw
* cell instance $7861 r0 *1 105.75,40.95
X$7861 366 31 367 644 645 cell_1rw
* cell instance $7862 r0 *1 106.455,40.95
X$7862 368 31 369 644 645 cell_1rw
* cell instance $7863 r0 *1 107.16,40.95
X$7863 370 31 371 644 645 cell_1rw
* cell instance $7864 r0 *1 107.865,40.95
X$7864 372 31 373 644 645 cell_1rw
* cell instance $7865 r0 *1 108.57,40.95
X$7865 374 31 375 644 645 cell_1rw
* cell instance $7866 r0 *1 109.275,40.95
X$7866 376 31 377 644 645 cell_1rw
* cell instance $7867 r0 *1 109.98,40.95
X$7867 378 31 379 644 645 cell_1rw
* cell instance $7868 r0 *1 110.685,40.95
X$7868 380 31 381 644 645 cell_1rw
* cell instance $7869 r0 *1 111.39,40.95
X$7869 382 31 383 644 645 cell_1rw
* cell instance $7870 r0 *1 112.095,40.95
X$7870 384 31 385 644 645 cell_1rw
* cell instance $7871 r0 *1 112.8,40.95
X$7871 386 31 387 644 645 cell_1rw
* cell instance $7872 r0 *1 113.505,40.95
X$7872 388 31 389 644 645 cell_1rw
* cell instance $7873 r0 *1 114.21,40.95
X$7873 390 31 391 644 645 cell_1rw
* cell instance $7874 r0 *1 114.915,40.95
X$7874 392 31 393 644 645 cell_1rw
* cell instance $7875 r0 *1 115.62,40.95
X$7875 394 31 395 644 645 cell_1rw
* cell instance $7876 r0 *1 116.325,40.95
X$7876 396 31 397 644 645 cell_1rw
* cell instance $7877 r0 *1 117.03,40.95
X$7877 398 31 399 644 645 cell_1rw
* cell instance $7878 r0 *1 117.735,40.95
X$7878 400 31 401 644 645 cell_1rw
* cell instance $7879 r0 *1 118.44,40.95
X$7879 402 31 403 644 645 cell_1rw
* cell instance $7880 r0 *1 119.145,40.95
X$7880 404 31 405 644 645 cell_1rw
* cell instance $7881 r0 *1 119.85,40.95
X$7881 406 31 407 644 645 cell_1rw
* cell instance $7882 r0 *1 120.555,40.95
X$7882 408 31 409 644 645 cell_1rw
* cell instance $7883 r0 *1 121.26,40.95
X$7883 410 31 411 644 645 cell_1rw
* cell instance $7884 r0 *1 121.965,40.95
X$7884 412 31 413 644 645 cell_1rw
* cell instance $7885 r0 *1 122.67,40.95
X$7885 414 31 415 644 645 cell_1rw
* cell instance $7886 r0 *1 123.375,40.95
X$7886 416 31 417 644 645 cell_1rw
* cell instance $7887 r0 *1 124.08,40.95
X$7887 418 31 419 644 645 cell_1rw
* cell instance $7888 r0 *1 124.785,40.95
X$7888 420 31 421 644 645 cell_1rw
* cell instance $7889 r0 *1 125.49,40.95
X$7889 422 31 423 644 645 cell_1rw
* cell instance $7890 r0 *1 126.195,40.95
X$7890 424 31 425 644 645 cell_1rw
* cell instance $7891 r0 *1 126.9,40.95
X$7891 426 31 427 644 645 cell_1rw
* cell instance $7892 r0 *1 127.605,40.95
X$7892 428 31 429 644 645 cell_1rw
* cell instance $7893 r0 *1 128.31,40.95
X$7893 430 31 431 644 645 cell_1rw
* cell instance $7894 r0 *1 129.015,40.95
X$7894 432 31 433 644 645 cell_1rw
* cell instance $7895 r0 *1 129.72,40.95
X$7895 434 31 435 644 645 cell_1rw
* cell instance $7896 r0 *1 130.425,40.95
X$7896 436 31 437 644 645 cell_1rw
* cell instance $7897 r0 *1 131.13,40.95
X$7897 438 31 439 644 645 cell_1rw
* cell instance $7898 r0 *1 131.835,40.95
X$7898 440 31 441 644 645 cell_1rw
* cell instance $7899 r0 *1 132.54,40.95
X$7899 442 31 443 644 645 cell_1rw
* cell instance $7900 r0 *1 133.245,40.95
X$7900 444 31 445 644 645 cell_1rw
* cell instance $7901 r0 *1 133.95,40.95
X$7901 446 31 447 644 645 cell_1rw
* cell instance $7902 r0 *1 134.655,40.95
X$7902 448 31 449 644 645 cell_1rw
* cell instance $7903 r0 *1 135.36,40.95
X$7903 450 31 451 644 645 cell_1rw
* cell instance $7904 r0 *1 136.065,40.95
X$7904 452 31 453 644 645 cell_1rw
* cell instance $7905 r0 *1 136.77,40.95
X$7905 454 31 455 644 645 cell_1rw
* cell instance $7906 r0 *1 137.475,40.95
X$7906 456 31 457 644 645 cell_1rw
* cell instance $7907 r0 *1 138.18,40.95
X$7907 458 31 459 644 645 cell_1rw
* cell instance $7908 r0 *1 138.885,40.95
X$7908 460 31 461 644 645 cell_1rw
* cell instance $7909 r0 *1 139.59,40.95
X$7909 462 31 463 644 645 cell_1rw
* cell instance $7910 r0 *1 140.295,40.95
X$7910 464 31 465 644 645 cell_1rw
* cell instance $7911 r0 *1 141,40.95
X$7911 466 31 467 644 645 cell_1rw
* cell instance $7912 r0 *1 141.705,40.95
X$7912 468 31 469 644 645 cell_1rw
* cell instance $7913 r0 *1 142.41,40.95
X$7913 470 31 471 644 645 cell_1rw
* cell instance $7914 r0 *1 143.115,40.95
X$7914 472 31 473 644 645 cell_1rw
* cell instance $7915 r0 *1 143.82,40.95
X$7915 474 31 475 644 645 cell_1rw
* cell instance $7916 r0 *1 144.525,40.95
X$7916 476 31 477 644 645 cell_1rw
* cell instance $7917 r0 *1 145.23,40.95
X$7917 478 31 479 644 645 cell_1rw
* cell instance $7918 r0 *1 145.935,40.95
X$7918 480 31 481 644 645 cell_1rw
* cell instance $7919 r0 *1 146.64,40.95
X$7919 482 31 483 644 645 cell_1rw
* cell instance $7920 r0 *1 147.345,40.95
X$7920 484 31 485 644 645 cell_1rw
* cell instance $7921 r0 *1 148.05,40.95
X$7921 486 31 487 644 645 cell_1rw
* cell instance $7922 r0 *1 148.755,40.95
X$7922 488 31 489 644 645 cell_1rw
* cell instance $7923 r0 *1 149.46,40.95
X$7923 490 31 491 644 645 cell_1rw
* cell instance $7924 r0 *1 150.165,40.95
X$7924 492 31 493 644 645 cell_1rw
* cell instance $7925 r0 *1 150.87,40.95
X$7925 494 31 495 644 645 cell_1rw
* cell instance $7926 r0 *1 151.575,40.95
X$7926 496 31 497 644 645 cell_1rw
* cell instance $7927 r0 *1 152.28,40.95
X$7927 498 31 499 644 645 cell_1rw
* cell instance $7928 r0 *1 152.985,40.95
X$7928 500 31 501 644 645 cell_1rw
* cell instance $7929 r0 *1 153.69,40.95
X$7929 502 31 503 644 645 cell_1rw
* cell instance $7930 r0 *1 154.395,40.95
X$7930 504 31 505 644 645 cell_1rw
* cell instance $7931 r0 *1 155.1,40.95
X$7931 506 31 507 644 645 cell_1rw
* cell instance $7932 r0 *1 155.805,40.95
X$7932 508 31 509 644 645 cell_1rw
* cell instance $7933 r0 *1 156.51,40.95
X$7933 510 31 511 644 645 cell_1rw
* cell instance $7934 r0 *1 157.215,40.95
X$7934 512 31 513 644 645 cell_1rw
* cell instance $7935 r0 *1 157.92,40.95
X$7935 514 31 515 644 645 cell_1rw
* cell instance $7936 r0 *1 158.625,40.95
X$7936 516 31 517 644 645 cell_1rw
* cell instance $7937 r0 *1 159.33,40.95
X$7937 518 31 519 644 645 cell_1rw
* cell instance $7938 r0 *1 160.035,40.95
X$7938 520 31 521 644 645 cell_1rw
* cell instance $7939 r0 *1 160.74,40.95
X$7939 522 31 523 644 645 cell_1rw
* cell instance $7940 r0 *1 161.445,40.95
X$7940 524 31 525 644 645 cell_1rw
* cell instance $7941 r0 *1 162.15,40.95
X$7941 526 31 527 644 645 cell_1rw
* cell instance $7942 r0 *1 162.855,40.95
X$7942 528 31 529 644 645 cell_1rw
* cell instance $7943 r0 *1 163.56,40.95
X$7943 530 31 531 644 645 cell_1rw
* cell instance $7944 r0 *1 164.265,40.95
X$7944 532 31 533 644 645 cell_1rw
* cell instance $7945 r0 *1 164.97,40.95
X$7945 534 31 535 644 645 cell_1rw
* cell instance $7946 r0 *1 165.675,40.95
X$7946 536 31 537 644 645 cell_1rw
* cell instance $7947 r0 *1 166.38,40.95
X$7947 538 31 539 644 645 cell_1rw
* cell instance $7948 r0 *1 167.085,40.95
X$7948 540 31 541 644 645 cell_1rw
* cell instance $7949 r0 *1 167.79,40.95
X$7949 542 31 543 644 645 cell_1rw
* cell instance $7950 r0 *1 168.495,40.95
X$7950 544 31 545 644 645 cell_1rw
* cell instance $7951 r0 *1 169.2,40.95
X$7951 546 31 547 644 645 cell_1rw
* cell instance $7952 r0 *1 169.905,40.95
X$7952 548 31 549 644 645 cell_1rw
* cell instance $7953 r0 *1 170.61,40.95
X$7953 550 31 551 644 645 cell_1rw
* cell instance $7954 r0 *1 171.315,40.95
X$7954 552 31 553 644 645 cell_1rw
* cell instance $7955 r0 *1 172.02,40.95
X$7955 554 31 555 644 645 cell_1rw
* cell instance $7956 r0 *1 172.725,40.95
X$7956 556 31 557 644 645 cell_1rw
* cell instance $7957 r0 *1 173.43,40.95
X$7957 558 31 559 644 645 cell_1rw
* cell instance $7958 r0 *1 174.135,40.95
X$7958 560 31 561 644 645 cell_1rw
* cell instance $7959 r0 *1 174.84,40.95
X$7959 562 31 563 644 645 cell_1rw
* cell instance $7960 r0 *1 175.545,40.95
X$7960 564 31 565 644 645 cell_1rw
* cell instance $7961 r0 *1 176.25,40.95
X$7961 566 31 567 644 645 cell_1rw
* cell instance $7962 r0 *1 176.955,40.95
X$7962 568 31 569 644 645 cell_1rw
* cell instance $7963 r0 *1 177.66,40.95
X$7963 570 31 571 644 645 cell_1rw
* cell instance $7964 r0 *1 178.365,40.95
X$7964 572 31 573 644 645 cell_1rw
* cell instance $7965 r0 *1 179.07,40.95
X$7965 574 31 575 644 645 cell_1rw
* cell instance $7966 r0 *1 179.775,40.95
X$7966 576 31 577 644 645 cell_1rw
* cell instance $7967 r0 *1 180.48,40.95
X$7967 578 31 579 644 645 cell_1rw
* cell instance $7968 m0 *1 0.705,43.68
X$7968 67 32 68 644 645 cell_1rw
* cell instance $7969 m0 *1 0,43.68
X$7969 65 32 66 644 645 cell_1rw
* cell instance $7970 m0 *1 1.41,43.68
X$7970 69 32 70 644 645 cell_1rw
* cell instance $7971 m0 *1 2.115,43.68
X$7971 71 32 72 644 645 cell_1rw
* cell instance $7972 m0 *1 2.82,43.68
X$7972 73 32 74 644 645 cell_1rw
* cell instance $7973 m0 *1 3.525,43.68
X$7973 75 32 76 644 645 cell_1rw
* cell instance $7974 m0 *1 4.23,43.68
X$7974 77 32 78 644 645 cell_1rw
* cell instance $7975 m0 *1 4.935,43.68
X$7975 79 32 80 644 645 cell_1rw
* cell instance $7976 m0 *1 5.64,43.68
X$7976 81 32 82 644 645 cell_1rw
* cell instance $7977 m0 *1 6.345,43.68
X$7977 83 32 84 644 645 cell_1rw
* cell instance $7978 m0 *1 7.05,43.68
X$7978 85 32 86 644 645 cell_1rw
* cell instance $7979 m0 *1 7.755,43.68
X$7979 87 32 88 644 645 cell_1rw
* cell instance $7980 m0 *1 8.46,43.68
X$7980 89 32 90 644 645 cell_1rw
* cell instance $7981 m0 *1 9.165,43.68
X$7981 91 32 92 644 645 cell_1rw
* cell instance $7982 m0 *1 9.87,43.68
X$7982 93 32 94 644 645 cell_1rw
* cell instance $7983 m0 *1 10.575,43.68
X$7983 95 32 96 644 645 cell_1rw
* cell instance $7984 m0 *1 11.28,43.68
X$7984 97 32 98 644 645 cell_1rw
* cell instance $7985 m0 *1 11.985,43.68
X$7985 99 32 100 644 645 cell_1rw
* cell instance $7986 m0 *1 12.69,43.68
X$7986 101 32 102 644 645 cell_1rw
* cell instance $7987 m0 *1 13.395,43.68
X$7987 103 32 104 644 645 cell_1rw
* cell instance $7988 m0 *1 14.1,43.68
X$7988 105 32 106 644 645 cell_1rw
* cell instance $7989 m0 *1 14.805,43.68
X$7989 107 32 108 644 645 cell_1rw
* cell instance $7990 m0 *1 15.51,43.68
X$7990 109 32 110 644 645 cell_1rw
* cell instance $7991 m0 *1 16.215,43.68
X$7991 111 32 112 644 645 cell_1rw
* cell instance $7992 m0 *1 16.92,43.68
X$7992 113 32 114 644 645 cell_1rw
* cell instance $7993 m0 *1 17.625,43.68
X$7993 115 32 116 644 645 cell_1rw
* cell instance $7994 m0 *1 18.33,43.68
X$7994 117 32 118 644 645 cell_1rw
* cell instance $7995 m0 *1 19.035,43.68
X$7995 119 32 120 644 645 cell_1rw
* cell instance $7996 m0 *1 19.74,43.68
X$7996 121 32 122 644 645 cell_1rw
* cell instance $7997 m0 *1 20.445,43.68
X$7997 123 32 124 644 645 cell_1rw
* cell instance $7998 m0 *1 21.15,43.68
X$7998 125 32 126 644 645 cell_1rw
* cell instance $7999 m0 *1 21.855,43.68
X$7999 127 32 128 644 645 cell_1rw
* cell instance $8000 m0 *1 22.56,43.68
X$8000 129 32 130 644 645 cell_1rw
* cell instance $8001 m0 *1 23.265,43.68
X$8001 131 32 132 644 645 cell_1rw
* cell instance $8002 m0 *1 23.97,43.68
X$8002 133 32 134 644 645 cell_1rw
* cell instance $8003 m0 *1 24.675,43.68
X$8003 135 32 136 644 645 cell_1rw
* cell instance $8004 m0 *1 25.38,43.68
X$8004 137 32 138 644 645 cell_1rw
* cell instance $8005 m0 *1 26.085,43.68
X$8005 139 32 140 644 645 cell_1rw
* cell instance $8006 m0 *1 26.79,43.68
X$8006 141 32 142 644 645 cell_1rw
* cell instance $8007 m0 *1 27.495,43.68
X$8007 143 32 144 644 645 cell_1rw
* cell instance $8008 m0 *1 28.2,43.68
X$8008 145 32 146 644 645 cell_1rw
* cell instance $8009 m0 *1 28.905,43.68
X$8009 147 32 148 644 645 cell_1rw
* cell instance $8010 m0 *1 29.61,43.68
X$8010 149 32 150 644 645 cell_1rw
* cell instance $8011 m0 *1 30.315,43.68
X$8011 151 32 152 644 645 cell_1rw
* cell instance $8012 m0 *1 31.02,43.68
X$8012 153 32 154 644 645 cell_1rw
* cell instance $8013 m0 *1 31.725,43.68
X$8013 155 32 156 644 645 cell_1rw
* cell instance $8014 m0 *1 32.43,43.68
X$8014 157 32 158 644 645 cell_1rw
* cell instance $8015 m0 *1 33.135,43.68
X$8015 159 32 160 644 645 cell_1rw
* cell instance $8016 m0 *1 33.84,43.68
X$8016 161 32 162 644 645 cell_1rw
* cell instance $8017 m0 *1 34.545,43.68
X$8017 163 32 164 644 645 cell_1rw
* cell instance $8018 m0 *1 35.25,43.68
X$8018 165 32 166 644 645 cell_1rw
* cell instance $8019 m0 *1 35.955,43.68
X$8019 167 32 168 644 645 cell_1rw
* cell instance $8020 m0 *1 36.66,43.68
X$8020 169 32 170 644 645 cell_1rw
* cell instance $8021 m0 *1 37.365,43.68
X$8021 171 32 172 644 645 cell_1rw
* cell instance $8022 m0 *1 38.07,43.68
X$8022 173 32 174 644 645 cell_1rw
* cell instance $8023 m0 *1 38.775,43.68
X$8023 175 32 176 644 645 cell_1rw
* cell instance $8024 m0 *1 39.48,43.68
X$8024 177 32 178 644 645 cell_1rw
* cell instance $8025 m0 *1 40.185,43.68
X$8025 179 32 180 644 645 cell_1rw
* cell instance $8026 m0 *1 40.89,43.68
X$8026 181 32 182 644 645 cell_1rw
* cell instance $8027 m0 *1 41.595,43.68
X$8027 183 32 184 644 645 cell_1rw
* cell instance $8028 m0 *1 42.3,43.68
X$8028 185 32 186 644 645 cell_1rw
* cell instance $8029 m0 *1 43.005,43.68
X$8029 187 32 188 644 645 cell_1rw
* cell instance $8030 m0 *1 43.71,43.68
X$8030 189 32 190 644 645 cell_1rw
* cell instance $8031 m0 *1 44.415,43.68
X$8031 191 32 192 644 645 cell_1rw
* cell instance $8032 m0 *1 45.12,43.68
X$8032 193 32 194 644 645 cell_1rw
* cell instance $8033 m0 *1 45.825,43.68
X$8033 195 32 196 644 645 cell_1rw
* cell instance $8034 m0 *1 46.53,43.68
X$8034 197 32 198 644 645 cell_1rw
* cell instance $8035 m0 *1 47.235,43.68
X$8035 199 32 200 644 645 cell_1rw
* cell instance $8036 m0 *1 47.94,43.68
X$8036 201 32 202 644 645 cell_1rw
* cell instance $8037 m0 *1 48.645,43.68
X$8037 203 32 204 644 645 cell_1rw
* cell instance $8038 m0 *1 49.35,43.68
X$8038 205 32 206 644 645 cell_1rw
* cell instance $8039 m0 *1 50.055,43.68
X$8039 207 32 208 644 645 cell_1rw
* cell instance $8040 m0 *1 50.76,43.68
X$8040 209 32 210 644 645 cell_1rw
* cell instance $8041 m0 *1 51.465,43.68
X$8041 211 32 212 644 645 cell_1rw
* cell instance $8042 m0 *1 52.17,43.68
X$8042 213 32 214 644 645 cell_1rw
* cell instance $8043 m0 *1 52.875,43.68
X$8043 215 32 216 644 645 cell_1rw
* cell instance $8044 m0 *1 53.58,43.68
X$8044 217 32 218 644 645 cell_1rw
* cell instance $8045 m0 *1 54.285,43.68
X$8045 219 32 220 644 645 cell_1rw
* cell instance $8046 m0 *1 54.99,43.68
X$8046 221 32 222 644 645 cell_1rw
* cell instance $8047 m0 *1 55.695,43.68
X$8047 223 32 224 644 645 cell_1rw
* cell instance $8048 m0 *1 56.4,43.68
X$8048 225 32 226 644 645 cell_1rw
* cell instance $8049 m0 *1 57.105,43.68
X$8049 227 32 228 644 645 cell_1rw
* cell instance $8050 m0 *1 57.81,43.68
X$8050 229 32 230 644 645 cell_1rw
* cell instance $8051 m0 *1 58.515,43.68
X$8051 231 32 232 644 645 cell_1rw
* cell instance $8052 m0 *1 59.22,43.68
X$8052 233 32 234 644 645 cell_1rw
* cell instance $8053 m0 *1 59.925,43.68
X$8053 235 32 236 644 645 cell_1rw
* cell instance $8054 m0 *1 60.63,43.68
X$8054 237 32 238 644 645 cell_1rw
* cell instance $8055 m0 *1 61.335,43.68
X$8055 239 32 240 644 645 cell_1rw
* cell instance $8056 m0 *1 62.04,43.68
X$8056 241 32 242 644 645 cell_1rw
* cell instance $8057 m0 *1 62.745,43.68
X$8057 243 32 244 644 645 cell_1rw
* cell instance $8058 m0 *1 63.45,43.68
X$8058 245 32 246 644 645 cell_1rw
* cell instance $8059 m0 *1 64.155,43.68
X$8059 247 32 248 644 645 cell_1rw
* cell instance $8060 m0 *1 64.86,43.68
X$8060 249 32 250 644 645 cell_1rw
* cell instance $8061 m0 *1 65.565,43.68
X$8061 251 32 252 644 645 cell_1rw
* cell instance $8062 m0 *1 66.27,43.68
X$8062 253 32 254 644 645 cell_1rw
* cell instance $8063 m0 *1 66.975,43.68
X$8063 255 32 256 644 645 cell_1rw
* cell instance $8064 m0 *1 67.68,43.68
X$8064 257 32 258 644 645 cell_1rw
* cell instance $8065 m0 *1 68.385,43.68
X$8065 259 32 260 644 645 cell_1rw
* cell instance $8066 m0 *1 69.09,43.68
X$8066 261 32 262 644 645 cell_1rw
* cell instance $8067 m0 *1 69.795,43.68
X$8067 263 32 264 644 645 cell_1rw
* cell instance $8068 m0 *1 70.5,43.68
X$8068 265 32 266 644 645 cell_1rw
* cell instance $8069 m0 *1 71.205,43.68
X$8069 267 32 268 644 645 cell_1rw
* cell instance $8070 m0 *1 71.91,43.68
X$8070 269 32 270 644 645 cell_1rw
* cell instance $8071 m0 *1 72.615,43.68
X$8071 271 32 272 644 645 cell_1rw
* cell instance $8072 m0 *1 73.32,43.68
X$8072 273 32 274 644 645 cell_1rw
* cell instance $8073 m0 *1 74.025,43.68
X$8073 275 32 276 644 645 cell_1rw
* cell instance $8074 m0 *1 74.73,43.68
X$8074 277 32 278 644 645 cell_1rw
* cell instance $8075 m0 *1 75.435,43.68
X$8075 279 32 280 644 645 cell_1rw
* cell instance $8076 m0 *1 76.14,43.68
X$8076 281 32 282 644 645 cell_1rw
* cell instance $8077 m0 *1 76.845,43.68
X$8077 283 32 284 644 645 cell_1rw
* cell instance $8078 m0 *1 77.55,43.68
X$8078 285 32 286 644 645 cell_1rw
* cell instance $8079 m0 *1 78.255,43.68
X$8079 287 32 288 644 645 cell_1rw
* cell instance $8080 m0 *1 78.96,43.68
X$8080 289 32 290 644 645 cell_1rw
* cell instance $8081 m0 *1 79.665,43.68
X$8081 291 32 292 644 645 cell_1rw
* cell instance $8082 m0 *1 80.37,43.68
X$8082 293 32 294 644 645 cell_1rw
* cell instance $8083 m0 *1 81.075,43.68
X$8083 295 32 296 644 645 cell_1rw
* cell instance $8084 m0 *1 81.78,43.68
X$8084 297 32 298 644 645 cell_1rw
* cell instance $8085 m0 *1 82.485,43.68
X$8085 299 32 300 644 645 cell_1rw
* cell instance $8086 m0 *1 83.19,43.68
X$8086 301 32 302 644 645 cell_1rw
* cell instance $8087 m0 *1 83.895,43.68
X$8087 303 32 304 644 645 cell_1rw
* cell instance $8088 m0 *1 84.6,43.68
X$8088 305 32 306 644 645 cell_1rw
* cell instance $8089 m0 *1 85.305,43.68
X$8089 307 32 308 644 645 cell_1rw
* cell instance $8090 m0 *1 86.01,43.68
X$8090 309 32 310 644 645 cell_1rw
* cell instance $8091 m0 *1 86.715,43.68
X$8091 311 32 312 644 645 cell_1rw
* cell instance $8092 m0 *1 87.42,43.68
X$8092 313 32 314 644 645 cell_1rw
* cell instance $8093 m0 *1 88.125,43.68
X$8093 315 32 316 644 645 cell_1rw
* cell instance $8094 m0 *1 88.83,43.68
X$8094 317 32 318 644 645 cell_1rw
* cell instance $8095 m0 *1 89.535,43.68
X$8095 319 32 320 644 645 cell_1rw
* cell instance $8096 m0 *1 90.24,43.68
X$8096 321 32 323 644 645 cell_1rw
* cell instance $8097 m0 *1 90.945,43.68
X$8097 324 32 325 644 645 cell_1rw
* cell instance $8098 m0 *1 91.65,43.68
X$8098 326 32 327 644 645 cell_1rw
* cell instance $8099 m0 *1 92.355,43.68
X$8099 328 32 329 644 645 cell_1rw
* cell instance $8100 m0 *1 93.06,43.68
X$8100 330 32 331 644 645 cell_1rw
* cell instance $8101 m0 *1 93.765,43.68
X$8101 332 32 333 644 645 cell_1rw
* cell instance $8102 m0 *1 94.47,43.68
X$8102 334 32 335 644 645 cell_1rw
* cell instance $8103 m0 *1 95.175,43.68
X$8103 336 32 337 644 645 cell_1rw
* cell instance $8104 m0 *1 95.88,43.68
X$8104 338 32 339 644 645 cell_1rw
* cell instance $8105 m0 *1 96.585,43.68
X$8105 340 32 341 644 645 cell_1rw
* cell instance $8106 m0 *1 97.29,43.68
X$8106 342 32 343 644 645 cell_1rw
* cell instance $8107 m0 *1 97.995,43.68
X$8107 344 32 345 644 645 cell_1rw
* cell instance $8108 m0 *1 98.7,43.68
X$8108 346 32 347 644 645 cell_1rw
* cell instance $8109 m0 *1 99.405,43.68
X$8109 348 32 349 644 645 cell_1rw
* cell instance $8110 m0 *1 100.11,43.68
X$8110 350 32 351 644 645 cell_1rw
* cell instance $8111 m0 *1 100.815,43.68
X$8111 352 32 353 644 645 cell_1rw
* cell instance $8112 m0 *1 101.52,43.68
X$8112 354 32 355 644 645 cell_1rw
* cell instance $8113 m0 *1 102.225,43.68
X$8113 356 32 357 644 645 cell_1rw
* cell instance $8114 m0 *1 102.93,43.68
X$8114 358 32 359 644 645 cell_1rw
* cell instance $8115 m0 *1 103.635,43.68
X$8115 360 32 361 644 645 cell_1rw
* cell instance $8116 m0 *1 104.34,43.68
X$8116 362 32 363 644 645 cell_1rw
* cell instance $8117 m0 *1 105.045,43.68
X$8117 364 32 365 644 645 cell_1rw
* cell instance $8118 m0 *1 105.75,43.68
X$8118 366 32 367 644 645 cell_1rw
* cell instance $8119 m0 *1 106.455,43.68
X$8119 368 32 369 644 645 cell_1rw
* cell instance $8120 m0 *1 107.16,43.68
X$8120 370 32 371 644 645 cell_1rw
* cell instance $8121 m0 *1 107.865,43.68
X$8121 372 32 373 644 645 cell_1rw
* cell instance $8122 m0 *1 108.57,43.68
X$8122 374 32 375 644 645 cell_1rw
* cell instance $8123 m0 *1 109.275,43.68
X$8123 376 32 377 644 645 cell_1rw
* cell instance $8124 m0 *1 109.98,43.68
X$8124 378 32 379 644 645 cell_1rw
* cell instance $8125 m0 *1 110.685,43.68
X$8125 380 32 381 644 645 cell_1rw
* cell instance $8126 m0 *1 111.39,43.68
X$8126 382 32 383 644 645 cell_1rw
* cell instance $8127 m0 *1 112.095,43.68
X$8127 384 32 385 644 645 cell_1rw
* cell instance $8128 m0 *1 112.8,43.68
X$8128 386 32 387 644 645 cell_1rw
* cell instance $8129 m0 *1 113.505,43.68
X$8129 388 32 389 644 645 cell_1rw
* cell instance $8130 m0 *1 114.21,43.68
X$8130 390 32 391 644 645 cell_1rw
* cell instance $8131 m0 *1 114.915,43.68
X$8131 392 32 393 644 645 cell_1rw
* cell instance $8132 m0 *1 115.62,43.68
X$8132 394 32 395 644 645 cell_1rw
* cell instance $8133 m0 *1 116.325,43.68
X$8133 396 32 397 644 645 cell_1rw
* cell instance $8134 m0 *1 117.03,43.68
X$8134 398 32 399 644 645 cell_1rw
* cell instance $8135 m0 *1 117.735,43.68
X$8135 400 32 401 644 645 cell_1rw
* cell instance $8136 m0 *1 118.44,43.68
X$8136 402 32 403 644 645 cell_1rw
* cell instance $8137 m0 *1 119.145,43.68
X$8137 404 32 405 644 645 cell_1rw
* cell instance $8138 m0 *1 119.85,43.68
X$8138 406 32 407 644 645 cell_1rw
* cell instance $8139 m0 *1 120.555,43.68
X$8139 408 32 409 644 645 cell_1rw
* cell instance $8140 m0 *1 121.26,43.68
X$8140 410 32 411 644 645 cell_1rw
* cell instance $8141 m0 *1 121.965,43.68
X$8141 412 32 413 644 645 cell_1rw
* cell instance $8142 m0 *1 122.67,43.68
X$8142 414 32 415 644 645 cell_1rw
* cell instance $8143 m0 *1 123.375,43.68
X$8143 416 32 417 644 645 cell_1rw
* cell instance $8144 m0 *1 124.08,43.68
X$8144 418 32 419 644 645 cell_1rw
* cell instance $8145 m0 *1 124.785,43.68
X$8145 420 32 421 644 645 cell_1rw
* cell instance $8146 m0 *1 125.49,43.68
X$8146 422 32 423 644 645 cell_1rw
* cell instance $8147 m0 *1 126.195,43.68
X$8147 424 32 425 644 645 cell_1rw
* cell instance $8148 m0 *1 126.9,43.68
X$8148 426 32 427 644 645 cell_1rw
* cell instance $8149 m0 *1 127.605,43.68
X$8149 428 32 429 644 645 cell_1rw
* cell instance $8150 m0 *1 128.31,43.68
X$8150 430 32 431 644 645 cell_1rw
* cell instance $8151 m0 *1 129.015,43.68
X$8151 432 32 433 644 645 cell_1rw
* cell instance $8152 m0 *1 129.72,43.68
X$8152 434 32 435 644 645 cell_1rw
* cell instance $8153 m0 *1 130.425,43.68
X$8153 436 32 437 644 645 cell_1rw
* cell instance $8154 m0 *1 131.13,43.68
X$8154 438 32 439 644 645 cell_1rw
* cell instance $8155 m0 *1 131.835,43.68
X$8155 440 32 441 644 645 cell_1rw
* cell instance $8156 m0 *1 132.54,43.68
X$8156 442 32 443 644 645 cell_1rw
* cell instance $8157 m0 *1 133.245,43.68
X$8157 444 32 445 644 645 cell_1rw
* cell instance $8158 m0 *1 133.95,43.68
X$8158 446 32 447 644 645 cell_1rw
* cell instance $8159 m0 *1 134.655,43.68
X$8159 448 32 449 644 645 cell_1rw
* cell instance $8160 m0 *1 135.36,43.68
X$8160 450 32 451 644 645 cell_1rw
* cell instance $8161 m0 *1 136.065,43.68
X$8161 452 32 453 644 645 cell_1rw
* cell instance $8162 m0 *1 136.77,43.68
X$8162 454 32 455 644 645 cell_1rw
* cell instance $8163 m0 *1 137.475,43.68
X$8163 456 32 457 644 645 cell_1rw
* cell instance $8164 m0 *1 138.18,43.68
X$8164 458 32 459 644 645 cell_1rw
* cell instance $8165 m0 *1 138.885,43.68
X$8165 460 32 461 644 645 cell_1rw
* cell instance $8166 m0 *1 139.59,43.68
X$8166 462 32 463 644 645 cell_1rw
* cell instance $8167 m0 *1 140.295,43.68
X$8167 464 32 465 644 645 cell_1rw
* cell instance $8168 m0 *1 141,43.68
X$8168 466 32 467 644 645 cell_1rw
* cell instance $8169 m0 *1 141.705,43.68
X$8169 468 32 469 644 645 cell_1rw
* cell instance $8170 m0 *1 142.41,43.68
X$8170 470 32 471 644 645 cell_1rw
* cell instance $8171 m0 *1 143.115,43.68
X$8171 472 32 473 644 645 cell_1rw
* cell instance $8172 m0 *1 143.82,43.68
X$8172 474 32 475 644 645 cell_1rw
* cell instance $8173 m0 *1 144.525,43.68
X$8173 476 32 477 644 645 cell_1rw
* cell instance $8174 m0 *1 145.23,43.68
X$8174 478 32 479 644 645 cell_1rw
* cell instance $8175 m0 *1 145.935,43.68
X$8175 480 32 481 644 645 cell_1rw
* cell instance $8176 m0 *1 146.64,43.68
X$8176 482 32 483 644 645 cell_1rw
* cell instance $8177 m0 *1 147.345,43.68
X$8177 484 32 485 644 645 cell_1rw
* cell instance $8178 m0 *1 148.05,43.68
X$8178 486 32 487 644 645 cell_1rw
* cell instance $8179 m0 *1 148.755,43.68
X$8179 488 32 489 644 645 cell_1rw
* cell instance $8180 m0 *1 149.46,43.68
X$8180 490 32 491 644 645 cell_1rw
* cell instance $8181 m0 *1 150.165,43.68
X$8181 492 32 493 644 645 cell_1rw
* cell instance $8182 m0 *1 150.87,43.68
X$8182 494 32 495 644 645 cell_1rw
* cell instance $8183 m0 *1 151.575,43.68
X$8183 496 32 497 644 645 cell_1rw
* cell instance $8184 m0 *1 152.28,43.68
X$8184 498 32 499 644 645 cell_1rw
* cell instance $8185 m0 *1 152.985,43.68
X$8185 500 32 501 644 645 cell_1rw
* cell instance $8186 m0 *1 153.69,43.68
X$8186 502 32 503 644 645 cell_1rw
* cell instance $8187 m0 *1 154.395,43.68
X$8187 504 32 505 644 645 cell_1rw
* cell instance $8188 m0 *1 155.1,43.68
X$8188 506 32 507 644 645 cell_1rw
* cell instance $8189 m0 *1 155.805,43.68
X$8189 508 32 509 644 645 cell_1rw
* cell instance $8190 m0 *1 156.51,43.68
X$8190 510 32 511 644 645 cell_1rw
* cell instance $8191 m0 *1 157.215,43.68
X$8191 512 32 513 644 645 cell_1rw
* cell instance $8192 m0 *1 157.92,43.68
X$8192 514 32 515 644 645 cell_1rw
* cell instance $8193 m0 *1 158.625,43.68
X$8193 516 32 517 644 645 cell_1rw
* cell instance $8194 m0 *1 159.33,43.68
X$8194 518 32 519 644 645 cell_1rw
* cell instance $8195 m0 *1 160.035,43.68
X$8195 520 32 521 644 645 cell_1rw
* cell instance $8196 m0 *1 160.74,43.68
X$8196 522 32 523 644 645 cell_1rw
* cell instance $8197 m0 *1 161.445,43.68
X$8197 524 32 525 644 645 cell_1rw
* cell instance $8198 m0 *1 162.15,43.68
X$8198 526 32 527 644 645 cell_1rw
* cell instance $8199 m0 *1 162.855,43.68
X$8199 528 32 529 644 645 cell_1rw
* cell instance $8200 m0 *1 163.56,43.68
X$8200 530 32 531 644 645 cell_1rw
* cell instance $8201 m0 *1 164.265,43.68
X$8201 532 32 533 644 645 cell_1rw
* cell instance $8202 m0 *1 164.97,43.68
X$8202 534 32 535 644 645 cell_1rw
* cell instance $8203 m0 *1 165.675,43.68
X$8203 536 32 537 644 645 cell_1rw
* cell instance $8204 m0 *1 166.38,43.68
X$8204 538 32 539 644 645 cell_1rw
* cell instance $8205 m0 *1 167.085,43.68
X$8205 540 32 541 644 645 cell_1rw
* cell instance $8206 m0 *1 167.79,43.68
X$8206 542 32 543 644 645 cell_1rw
* cell instance $8207 m0 *1 168.495,43.68
X$8207 544 32 545 644 645 cell_1rw
* cell instance $8208 m0 *1 169.2,43.68
X$8208 546 32 547 644 645 cell_1rw
* cell instance $8209 m0 *1 169.905,43.68
X$8209 548 32 549 644 645 cell_1rw
* cell instance $8210 m0 *1 170.61,43.68
X$8210 550 32 551 644 645 cell_1rw
* cell instance $8211 m0 *1 171.315,43.68
X$8211 552 32 553 644 645 cell_1rw
* cell instance $8212 m0 *1 172.02,43.68
X$8212 554 32 555 644 645 cell_1rw
* cell instance $8213 m0 *1 172.725,43.68
X$8213 556 32 557 644 645 cell_1rw
* cell instance $8214 m0 *1 173.43,43.68
X$8214 558 32 559 644 645 cell_1rw
* cell instance $8215 m0 *1 174.135,43.68
X$8215 560 32 561 644 645 cell_1rw
* cell instance $8216 m0 *1 174.84,43.68
X$8216 562 32 563 644 645 cell_1rw
* cell instance $8217 m0 *1 175.545,43.68
X$8217 564 32 565 644 645 cell_1rw
* cell instance $8218 m0 *1 176.25,43.68
X$8218 566 32 567 644 645 cell_1rw
* cell instance $8219 m0 *1 176.955,43.68
X$8219 568 32 569 644 645 cell_1rw
* cell instance $8220 m0 *1 177.66,43.68
X$8220 570 32 571 644 645 cell_1rw
* cell instance $8221 m0 *1 178.365,43.68
X$8221 572 32 573 644 645 cell_1rw
* cell instance $8222 m0 *1 179.07,43.68
X$8222 574 32 575 644 645 cell_1rw
* cell instance $8223 m0 *1 179.775,43.68
X$8223 576 32 577 644 645 cell_1rw
* cell instance $8224 m0 *1 180.48,43.68
X$8224 578 32 579 644 645 cell_1rw
* cell instance $8225 r0 *1 0.705,43.68
X$8225 67 33 68 644 645 cell_1rw
* cell instance $8226 r0 *1 0,43.68
X$8226 65 33 66 644 645 cell_1rw
* cell instance $8227 r0 *1 1.41,43.68
X$8227 69 33 70 644 645 cell_1rw
* cell instance $8228 r0 *1 2.115,43.68
X$8228 71 33 72 644 645 cell_1rw
* cell instance $8229 r0 *1 2.82,43.68
X$8229 73 33 74 644 645 cell_1rw
* cell instance $8230 r0 *1 3.525,43.68
X$8230 75 33 76 644 645 cell_1rw
* cell instance $8231 r0 *1 4.23,43.68
X$8231 77 33 78 644 645 cell_1rw
* cell instance $8232 r0 *1 4.935,43.68
X$8232 79 33 80 644 645 cell_1rw
* cell instance $8233 r0 *1 5.64,43.68
X$8233 81 33 82 644 645 cell_1rw
* cell instance $8234 r0 *1 6.345,43.68
X$8234 83 33 84 644 645 cell_1rw
* cell instance $8235 r0 *1 7.05,43.68
X$8235 85 33 86 644 645 cell_1rw
* cell instance $8236 r0 *1 7.755,43.68
X$8236 87 33 88 644 645 cell_1rw
* cell instance $8237 r0 *1 8.46,43.68
X$8237 89 33 90 644 645 cell_1rw
* cell instance $8238 r0 *1 9.165,43.68
X$8238 91 33 92 644 645 cell_1rw
* cell instance $8239 r0 *1 9.87,43.68
X$8239 93 33 94 644 645 cell_1rw
* cell instance $8240 r0 *1 10.575,43.68
X$8240 95 33 96 644 645 cell_1rw
* cell instance $8241 r0 *1 11.28,43.68
X$8241 97 33 98 644 645 cell_1rw
* cell instance $8242 r0 *1 11.985,43.68
X$8242 99 33 100 644 645 cell_1rw
* cell instance $8243 r0 *1 12.69,43.68
X$8243 101 33 102 644 645 cell_1rw
* cell instance $8244 r0 *1 13.395,43.68
X$8244 103 33 104 644 645 cell_1rw
* cell instance $8245 r0 *1 14.1,43.68
X$8245 105 33 106 644 645 cell_1rw
* cell instance $8246 r0 *1 14.805,43.68
X$8246 107 33 108 644 645 cell_1rw
* cell instance $8247 r0 *1 15.51,43.68
X$8247 109 33 110 644 645 cell_1rw
* cell instance $8248 r0 *1 16.215,43.68
X$8248 111 33 112 644 645 cell_1rw
* cell instance $8249 r0 *1 16.92,43.68
X$8249 113 33 114 644 645 cell_1rw
* cell instance $8250 r0 *1 17.625,43.68
X$8250 115 33 116 644 645 cell_1rw
* cell instance $8251 r0 *1 18.33,43.68
X$8251 117 33 118 644 645 cell_1rw
* cell instance $8252 r0 *1 19.035,43.68
X$8252 119 33 120 644 645 cell_1rw
* cell instance $8253 r0 *1 19.74,43.68
X$8253 121 33 122 644 645 cell_1rw
* cell instance $8254 r0 *1 20.445,43.68
X$8254 123 33 124 644 645 cell_1rw
* cell instance $8255 r0 *1 21.15,43.68
X$8255 125 33 126 644 645 cell_1rw
* cell instance $8256 r0 *1 21.855,43.68
X$8256 127 33 128 644 645 cell_1rw
* cell instance $8257 r0 *1 22.56,43.68
X$8257 129 33 130 644 645 cell_1rw
* cell instance $8258 r0 *1 23.265,43.68
X$8258 131 33 132 644 645 cell_1rw
* cell instance $8259 r0 *1 23.97,43.68
X$8259 133 33 134 644 645 cell_1rw
* cell instance $8260 r0 *1 24.675,43.68
X$8260 135 33 136 644 645 cell_1rw
* cell instance $8261 r0 *1 25.38,43.68
X$8261 137 33 138 644 645 cell_1rw
* cell instance $8262 r0 *1 26.085,43.68
X$8262 139 33 140 644 645 cell_1rw
* cell instance $8263 r0 *1 26.79,43.68
X$8263 141 33 142 644 645 cell_1rw
* cell instance $8264 r0 *1 27.495,43.68
X$8264 143 33 144 644 645 cell_1rw
* cell instance $8265 r0 *1 28.2,43.68
X$8265 145 33 146 644 645 cell_1rw
* cell instance $8266 r0 *1 28.905,43.68
X$8266 147 33 148 644 645 cell_1rw
* cell instance $8267 r0 *1 29.61,43.68
X$8267 149 33 150 644 645 cell_1rw
* cell instance $8268 r0 *1 30.315,43.68
X$8268 151 33 152 644 645 cell_1rw
* cell instance $8269 r0 *1 31.02,43.68
X$8269 153 33 154 644 645 cell_1rw
* cell instance $8270 r0 *1 31.725,43.68
X$8270 155 33 156 644 645 cell_1rw
* cell instance $8271 r0 *1 32.43,43.68
X$8271 157 33 158 644 645 cell_1rw
* cell instance $8272 r0 *1 33.135,43.68
X$8272 159 33 160 644 645 cell_1rw
* cell instance $8273 r0 *1 33.84,43.68
X$8273 161 33 162 644 645 cell_1rw
* cell instance $8274 r0 *1 34.545,43.68
X$8274 163 33 164 644 645 cell_1rw
* cell instance $8275 r0 *1 35.25,43.68
X$8275 165 33 166 644 645 cell_1rw
* cell instance $8276 r0 *1 35.955,43.68
X$8276 167 33 168 644 645 cell_1rw
* cell instance $8277 r0 *1 36.66,43.68
X$8277 169 33 170 644 645 cell_1rw
* cell instance $8278 r0 *1 37.365,43.68
X$8278 171 33 172 644 645 cell_1rw
* cell instance $8279 r0 *1 38.07,43.68
X$8279 173 33 174 644 645 cell_1rw
* cell instance $8280 r0 *1 38.775,43.68
X$8280 175 33 176 644 645 cell_1rw
* cell instance $8281 r0 *1 39.48,43.68
X$8281 177 33 178 644 645 cell_1rw
* cell instance $8282 r0 *1 40.185,43.68
X$8282 179 33 180 644 645 cell_1rw
* cell instance $8283 r0 *1 40.89,43.68
X$8283 181 33 182 644 645 cell_1rw
* cell instance $8284 r0 *1 41.595,43.68
X$8284 183 33 184 644 645 cell_1rw
* cell instance $8285 r0 *1 42.3,43.68
X$8285 185 33 186 644 645 cell_1rw
* cell instance $8286 r0 *1 43.005,43.68
X$8286 187 33 188 644 645 cell_1rw
* cell instance $8287 r0 *1 43.71,43.68
X$8287 189 33 190 644 645 cell_1rw
* cell instance $8288 r0 *1 44.415,43.68
X$8288 191 33 192 644 645 cell_1rw
* cell instance $8289 r0 *1 45.12,43.68
X$8289 193 33 194 644 645 cell_1rw
* cell instance $8290 r0 *1 45.825,43.68
X$8290 195 33 196 644 645 cell_1rw
* cell instance $8291 r0 *1 46.53,43.68
X$8291 197 33 198 644 645 cell_1rw
* cell instance $8292 r0 *1 47.235,43.68
X$8292 199 33 200 644 645 cell_1rw
* cell instance $8293 r0 *1 47.94,43.68
X$8293 201 33 202 644 645 cell_1rw
* cell instance $8294 r0 *1 48.645,43.68
X$8294 203 33 204 644 645 cell_1rw
* cell instance $8295 r0 *1 49.35,43.68
X$8295 205 33 206 644 645 cell_1rw
* cell instance $8296 r0 *1 50.055,43.68
X$8296 207 33 208 644 645 cell_1rw
* cell instance $8297 r0 *1 50.76,43.68
X$8297 209 33 210 644 645 cell_1rw
* cell instance $8298 r0 *1 51.465,43.68
X$8298 211 33 212 644 645 cell_1rw
* cell instance $8299 r0 *1 52.17,43.68
X$8299 213 33 214 644 645 cell_1rw
* cell instance $8300 r0 *1 52.875,43.68
X$8300 215 33 216 644 645 cell_1rw
* cell instance $8301 r0 *1 53.58,43.68
X$8301 217 33 218 644 645 cell_1rw
* cell instance $8302 r0 *1 54.285,43.68
X$8302 219 33 220 644 645 cell_1rw
* cell instance $8303 r0 *1 54.99,43.68
X$8303 221 33 222 644 645 cell_1rw
* cell instance $8304 r0 *1 55.695,43.68
X$8304 223 33 224 644 645 cell_1rw
* cell instance $8305 r0 *1 56.4,43.68
X$8305 225 33 226 644 645 cell_1rw
* cell instance $8306 r0 *1 57.105,43.68
X$8306 227 33 228 644 645 cell_1rw
* cell instance $8307 r0 *1 57.81,43.68
X$8307 229 33 230 644 645 cell_1rw
* cell instance $8308 r0 *1 58.515,43.68
X$8308 231 33 232 644 645 cell_1rw
* cell instance $8309 r0 *1 59.22,43.68
X$8309 233 33 234 644 645 cell_1rw
* cell instance $8310 r0 *1 59.925,43.68
X$8310 235 33 236 644 645 cell_1rw
* cell instance $8311 r0 *1 60.63,43.68
X$8311 237 33 238 644 645 cell_1rw
* cell instance $8312 r0 *1 61.335,43.68
X$8312 239 33 240 644 645 cell_1rw
* cell instance $8313 r0 *1 62.04,43.68
X$8313 241 33 242 644 645 cell_1rw
* cell instance $8314 r0 *1 62.745,43.68
X$8314 243 33 244 644 645 cell_1rw
* cell instance $8315 r0 *1 63.45,43.68
X$8315 245 33 246 644 645 cell_1rw
* cell instance $8316 r0 *1 64.155,43.68
X$8316 247 33 248 644 645 cell_1rw
* cell instance $8317 r0 *1 64.86,43.68
X$8317 249 33 250 644 645 cell_1rw
* cell instance $8318 r0 *1 65.565,43.68
X$8318 251 33 252 644 645 cell_1rw
* cell instance $8319 r0 *1 66.27,43.68
X$8319 253 33 254 644 645 cell_1rw
* cell instance $8320 r0 *1 66.975,43.68
X$8320 255 33 256 644 645 cell_1rw
* cell instance $8321 r0 *1 67.68,43.68
X$8321 257 33 258 644 645 cell_1rw
* cell instance $8322 r0 *1 68.385,43.68
X$8322 259 33 260 644 645 cell_1rw
* cell instance $8323 r0 *1 69.09,43.68
X$8323 261 33 262 644 645 cell_1rw
* cell instance $8324 r0 *1 69.795,43.68
X$8324 263 33 264 644 645 cell_1rw
* cell instance $8325 r0 *1 70.5,43.68
X$8325 265 33 266 644 645 cell_1rw
* cell instance $8326 r0 *1 71.205,43.68
X$8326 267 33 268 644 645 cell_1rw
* cell instance $8327 r0 *1 71.91,43.68
X$8327 269 33 270 644 645 cell_1rw
* cell instance $8328 r0 *1 72.615,43.68
X$8328 271 33 272 644 645 cell_1rw
* cell instance $8329 r0 *1 73.32,43.68
X$8329 273 33 274 644 645 cell_1rw
* cell instance $8330 r0 *1 74.025,43.68
X$8330 275 33 276 644 645 cell_1rw
* cell instance $8331 r0 *1 74.73,43.68
X$8331 277 33 278 644 645 cell_1rw
* cell instance $8332 r0 *1 75.435,43.68
X$8332 279 33 280 644 645 cell_1rw
* cell instance $8333 r0 *1 76.14,43.68
X$8333 281 33 282 644 645 cell_1rw
* cell instance $8334 r0 *1 76.845,43.68
X$8334 283 33 284 644 645 cell_1rw
* cell instance $8335 r0 *1 77.55,43.68
X$8335 285 33 286 644 645 cell_1rw
* cell instance $8336 r0 *1 78.255,43.68
X$8336 287 33 288 644 645 cell_1rw
* cell instance $8337 r0 *1 78.96,43.68
X$8337 289 33 290 644 645 cell_1rw
* cell instance $8338 r0 *1 79.665,43.68
X$8338 291 33 292 644 645 cell_1rw
* cell instance $8339 r0 *1 80.37,43.68
X$8339 293 33 294 644 645 cell_1rw
* cell instance $8340 r0 *1 81.075,43.68
X$8340 295 33 296 644 645 cell_1rw
* cell instance $8341 r0 *1 81.78,43.68
X$8341 297 33 298 644 645 cell_1rw
* cell instance $8342 r0 *1 82.485,43.68
X$8342 299 33 300 644 645 cell_1rw
* cell instance $8343 r0 *1 83.19,43.68
X$8343 301 33 302 644 645 cell_1rw
* cell instance $8344 r0 *1 83.895,43.68
X$8344 303 33 304 644 645 cell_1rw
* cell instance $8345 r0 *1 84.6,43.68
X$8345 305 33 306 644 645 cell_1rw
* cell instance $8346 r0 *1 85.305,43.68
X$8346 307 33 308 644 645 cell_1rw
* cell instance $8347 r0 *1 86.01,43.68
X$8347 309 33 310 644 645 cell_1rw
* cell instance $8348 r0 *1 86.715,43.68
X$8348 311 33 312 644 645 cell_1rw
* cell instance $8349 r0 *1 87.42,43.68
X$8349 313 33 314 644 645 cell_1rw
* cell instance $8350 r0 *1 88.125,43.68
X$8350 315 33 316 644 645 cell_1rw
* cell instance $8351 r0 *1 88.83,43.68
X$8351 317 33 318 644 645 cell_1rw
* cell instance $8352 r0 *1 89.535,43.68
X$8352 319 33 320 644 645 cell_1rw
* cell instance $8353 r0 *1 90.24,43.68
X$8353 321 33 323 644 645 cell_1rw
* cell instance $8354 r0 *1 90.945,43.68
X$8354 324 33 325 644 645 cell_1rw
* cell instance $8355 r0 *1 91.65,43.68
X$8355 326 33 327 644 645 cell_1rw
* cell instance $8356 r0 *1 92.355,43.68
X$8356 328 33 329 644 645 cell_1rw
* cell instance $8357 r0 *1 93.06,43.68
X$8357 330 33 331 644 645 cell_1rw
* cell instance $8358 r0 *1 93.765,43.68
X$8358 332 33 333 644 645 cell_1rw
* cell instance $8359 r0 *1 94.47,43.68
X$8359 334 33 335 644 645 cell_1rw
* cell instance $8360 r0 *1 95.175,43.68
X$8360 336 33 337 644 645 cell_1rw
* cell instance $8361 r0 *1 95.88,43.68
X$8361 338 33 339 644 645 cell_1rw
* cell instance $8362 r0 *1 96.585,43.68
X$8362 340 33 341 644 645 cell_1rw
* cell instance $8363 r0 *1 97.29,43.68
X$8363 342 33 343 644 645 cell_1rw
* cell instance $8364 r0 *1 97.995,43.68
X$8364 344 33 345 644 645 cell_1rw
* cell instance $8365 r0 *1 98.7,43.68
X$8365 346 33 347 644 645 cell_1rw
* cell instance $8366 r0 *1 99.405,43.68
X$8366 348 33 349 644 645 cell_1rw
* cell instance $8367 r0 *1 100.11,43.68
X$8367 350 33 351 644 645 cell_1rw
* cell instance $8368 r0 *1 100.815,43.68
X$8368 352 33 353 644 645 cell_1rw
* cell instance $8369 r0 *1 101.52,43.68
X$8369 354 33 355 644 645 cell_1rw
* cell instance $8370 r0 *1 102.225,43.68
X$8370 356 33 357 644 645 cell_1rw
* cell instance $8371 r0 *1 102.93,43.68
X$8371 358 33 359 644 645 cell_1rw
* cell instance $8372 r0 *1 103.635,43.68
X$8372 360 33 361 644 645 cell_1rw
* cell instance $8373 r0 *1 104.34,43.68
X$8373 362 33 363 644 645 cell_1rw
* cell instance $8374 r0 *1 105.045,43.68
X$8374 364 33 365 644 645 cell_1rw
* cell instance $8375 r0 *1 105.75,43.68
X$8375 366 33 367 644 645 cell_1rw
* cell instance $8376 r0 *1 106.455,43.68
X$8376 368 33 369 644 645 cell_1rw
* cell instance $8377 r0 *1 107.16,43.68
X$8377 370 33 371 644 645 cell_1rw
* cell instance $8378 r0 *1 107.865,43.68
X$8378 372 33 373 644 645 cell_1rw
* cell instance $8379 r0 *1 108.57,43.68
X$8379 374 33 375 644 645 cell_1rw
* cell instance $8380 r0 *1 109.275,43.68
X$8380 376 33 377 644 645 cell_1rw
* cell instance $8381 r0 *1 109.98,43.68
X$8381 378 33 379 644 645 cell_1rw
* cell instance $8382 r0 *1 110.685,43.68
X$8382 380 33 381 644 645 cell_1rw
* cell instance $8383 r0 *1 111.39,43.68
X$8383 382 33 383 644 645 cell_1rw
* cell instance $8384 r0 *1 112.095,43.68
X$8384 384 33 385 644 645 cell_1rw
* cell instance $8385 r0 *1 112.8,43.68
X$8385 386 33 387 644 645 cell_1rw
* cell instance $8386 r0 *1 113.505,43.68
X$8386 388 33 389 644 645 cell_1rw
* cell instance $8387 r0 *1 114.21,43.68
X$8387 390 33 391 644 645 cell_1rw
* cell instance $8388 r0 *1 114.915,43.68
X$8388 392 33 393 644 645 cell_1rw
* cell instance $8389 r0 *1 115.62,43.68
X$8389 394 33 395 644 645 cell_1rw
* cell instance $8390 r0 *1 116.325,43.68
X$8390 396 33 397 644 645 cell_1rw
* cell instance $8391 r0 *1 117.03,43.68
X$8391 398 33 399 644 645 cell_1rw
* cell instance $8392 r0 *1 117.735,43.68
X$8392 400 33 401 644 645 cell_1rw
* cell instance $8393 r0 *1 118.44,43.68
X$8393 402 33 403 644 645 cell_1rw
* cell instance $8394 r0 *1 119.145,43.68
X$8394 404 33 405 644 645 cell_1rw
* cell instance $8395 r0 *1 119.85,43.68
X$8395 406 33 407 644 645 cell_1rw
* cell instance $8396 r0 *1 120.555,43.68
X$8396 408 33 409 644 645 cell_1rw
* cell instance $8397 r0 *1 121.26,43.68
X$8397 410 33 411 644 645 cell_1rw
* cell instance $8398 r0 *1 121.965,43.68
X$8398 412 33 413 644 645 cell_1rw
* cell instance $8399 r0 *1 122.67,43.68
X$8399 414 33 415 644 645 cell_1rw
* cell instance $8400 r0 *1 123.375,43.68
X$8400 416 33 417 644 645 cell_1rw
* cell instance $8401 r0 *1 124.08,43.68
X$8401 418 33 419 644 645 cell_1rw
* cell instance $8402 r0 *1 124.785,43.68
X$8402 420 33 421 644 645 cell_1rw
* cell instance $8403 r0 *1 125.49,43.68
X$8403 422 33 423 644 645 cell_1rw
* cell instance $8404 r0 *1 126.195,43.68
X$8404 424 33 425 644 645 cell_1rw
* cell instance $8405 r0 *1 126.9,43.68
X$8405 426 33 427 644 645 cell_1rw
* cell instance $8406 r0 *1 127.605,43.68
X$8406 428 33 429 644 645 cell_1rw
* cell instance $8407 r0 *1 128.31,43.68
X$8407 430 33 431 644 645 cell_1rw
* cell instance $8408 r0 *1 129.015,43.68
X$8408 432 33 433 644 645 cell_1rw
* cell instance $8409 r0 *1 129.72,43.68
X$8409 434 33 435 644 645 cell_1rw
* cell instance $8410 r0 *1 130.425,43.68
X$8410 436 33 437 644 645 cell_1rw
* cell instance $8411 r0 *1 131.13,43.68
X$8411 438 33 439 644 645 cell_1rw
* cell instance $8412 r0 *1 131.835,43.68
X$8412 440 33 441 644 645 cell_1rw
* cell instance $8413 r0 *1 132.54,43.68
X$8413 442 33 443 644 645 cell_1rw
* cell instance $8414 r0 *1 133.245,43.68
X$8414 444 33 445 644 645 cell_1rw
* cell instance $8415 r0 *1 133.95,43.68
X$8415 446 33 447 644 645 cell_1rw
* cell instance $8416 r0 *1 134.655,43.68
X$8416 448 33 449 644 645 cell_1rw
* cell instance $8417 r0 *1 135.36,43.68
X$8417 450 33 451 644 645 cell_1rw
* cell instance $8418 r0 *1 136.065,43.68
X$8418 452 33 453 644 645 cell_1rw
* cell instance $8419 r0 *1 136.77,43.68
X$8419 454 33 455 644 645 cell_1rw
* cell instance $8420 r0 *1 137.475,43.68
X$8420 456 33 457 644 645 cell_1rw
* cell instance $8421 r0 *1 138.18,43.68
X$8421 458 33 459 644 645 cell_1rw
* cell instance $8422 r0 *1 138.885,43.68
X$8422 460 33 461 644 645 cell_1rw
* cell instance $8423 r0 *1 139.59,43.68
X$8423 462 33 463 644 645 cell_1rw
* cell instance $8424 r0 *1 140.295,43.68
X$8424 464 33 465 644 645 cell_1rw
* cell instance $8425 r0 *1 141,43.68
X$8425 466 33 467 644 645 cell_1rw
* cell instance $8426 r0 *1 141.705,43.68
X$8426 468 33 469 644 645 cell_1rw
* cell instance $8427 r0 *1 142.41,43.68
X$8427 470 33 471 644 645 cell_1rw
* cell instance $8428 r0 *1 143.115,43.68
X$8428 472 33 473 644 645 cell_1rw
* cell instance $8429 r0 *1 143.82,43.68
X$8429 474 33 475 644 645 cell_1rw
* cell instance $8430 r0 *1 144.525,43.68
X$8430 476 33 477 644 645 cell_1rw
* cell instance $8431 r0 *1 145.23,43.68
X$8431 478 33 479 644 645 cell_1rw
* cell instance $8432 r0 *1 145.935,43.68
X$8432 480 33 481 644 645 cell_1rw
* cell instance $8433 r0 *1 146.64,43.68
X$8433 482 33 483 644 645 cell_1rw
* cell instance $8434 r0 *1 147.345,43.68
X$8434 484 33 485 644 645 cell_1rw
* cell instance $8435 r0 *1 148.05,43.68
X$8435 486 33 487 644 645 cell_1rw
* cell instance $8436 r0 *1 148.755,43.68
X$8436 488 33 489 644 645 cell_1rw
* cell instance $8437 r0 *1 149.46,43.68
X$8437 490 33 491 644 645 cell_1rw
* cell instance $8438 r0 *1 150.165,43.68
X$8438 492 33 493 644 645 cell_1rw
* cell instance $8439 r0 *1 150.87,43.68
X$8439 494 33 495 644 645 cell_1rw
* cell instance $8440 r0 *1 151.575,43.68
X$8440 496 33 497 644 645 cell_1rw
* cell instance $8441 r0 *1 152.28,43.68
X$8441 498 33 499 644 645 cell_1rw
* cell instance $8442 r0 *1 152.985,43.68
X$8442 500 33 501 644 645 cell_1rw
* cell instance $8443 r0 *1 153.69,43.68
X$8443 502 33 503 644 645 cell_1rw
* cell instance $8444 r0 *1 154.395,43.68
X$8444 504 33 505 644 645 cell_1rw
* cell instance $8445 r0 *1 155.1,43.68
X$8445 506 33 507 644 645 cell_1rw
* cell instance $8446 r0 *1 155.805,43.68
X$8446 508 33 509 644 645 cell_1rw
* cell instance $8447 r0 *1 156.51,43.68
X$8447 510 33 511 644 645 cell_1rw
* cell instance $8448 r0 *1 157.215,43.68
X$8448 512 33 513 644 645 cell_1rw
* cell instance $8449 r0 *1 157.92,43.68
X$8449 514 33 515 644 645 cell_1rw
* cell instance $8450 r0 *1 158.625,43.68
X$8450 516 33 517 644 645 cell_1rw
* cell instance $8451 r0 *1 159.33,43.68
X$8451 518 33 519 644 645 cell_1rw
* cell instance $8452 r0 *1 160.035,43.68
X$8452 520 33 521 644 645 cell_1rw
* cell instance $8453 r0 *1 160.74,43.68
X$8453 522 33 523 644 645 cell_1rw
* cell instance $8454 r0 *1 161.445,43.68
X$8454 524 33 525 644 645 cell_1rw
* cell instance $8455 r0 *1 162.15,43.68
X$8455 526 33 527 644 645 cell_1rw
* cell instance $8456 r0 *1 162.855,43.68
X$8456 528 33 529 644 645 cell_1rw
* cell instance $8457 r0 *1 163.56,43.68
X$8457 530 33 531 644 645 cell_1rw
* cell instance $8458 r0 *1 164.265,43.68
X$8458 532 33 533 644 645 cell_1rw
* cell instance $8459 r0 *1 164.97,43.68
X$8459 534 33 535 644 645 cell_1rw
* cell instance $8460 r0 *1 165.675,43.68
X$8460 536 33 537 644 645 cell_1rw
* cell instance $8461 r0 *1 166.38,43.68
X$8461 538 33 539 644 645 cell_1rw
* cell instance $8462 r0 *1 167.085,43.68
X$8462 540 33 541 644 645 cell_1rw
* cell instance $8463 r0 *1 167.79,43.68
X$8463 542 33 543 644 645 cell_1rw
* cell instance $8464 r0 *1 168.495,43.68
X$8464 544 33 545 644 645 cell_1rw
* cell instance $8465 r0 *1 169.2,43.68
X$8465 546 33 547 644 645 cell_1rw
* cell instance $8466 r0 *1 169.905,43.68
X$8466 548 33 549 644 645 cell_1rw
* cell instance $8467 r0 *1 170.61,43.68
X$8467 550 33 551 644 645 cell_1rw
* cell instance $8468 r0 *1 171.315,43.68
X$8468 552 33 553 644 645 cell_1rw
* cell instance $8469 r0 *1 172.02,43.68
X$8469 554 33 555 644 645 cell_1rw
* cell instance $8470 r0 *1 172.725,43.68
X$8470 556 33 557 644 645 cell_1rw
* cell instance $8471 r0 *1 173.43,43.68
X$8471 558 33 559 644 645 cell_1rw
* cell instance $8472 r0 *1 174.135,43.68
X$8472 560 33 561 644 645 cell_1rw
* cell instance $8473 r0 *1 174.84,43.68
X$8473 562 33 563 644 645 cell_1rw
* cell instance $8474 r0 *1 175.545,43.68
X$8474 564 33 565 644 645 cell_1rw
* cell instance $8475 r0 *1 176.25,43.68
X$8475 566 33 567 644 645 cell_1rw
* cell instance $8476 r0 *1 176.955,43.68
X$8476 568 33 569 644 645 cell_1rw
* cell instance $8477 r0 *1 177.66,43.68
X$8477 570 33 571 644 645 cell_1rw
* cell instance $8478 r0 *1 178.365,43.68
X$8478 572 33 573 644 645 cell_1rw
* cell instance $8479 r0 *1 179.07,43.68
X$8479 574 33 575 644 645 cell_1rw
* cell instance $8480 r0 *1 179.775,43.68
X$8480 576 33 577 644 645 cell_1rw
* cell instance $8481 r0 *1 180.48,43.68
X$8481 578 33 579 644 645 cell_1rw
* cell instance $8482 m0 *1 0.705,46.41
X$8482 67 34 68 644 645 cell_1rw
* cell instance $8483 m0 *1 0,46.41
X$8483 65 34 66 644 645 cell_1rw
* cell instance $8484 m0 *1 1.41,46.41
X$8484 69 34 70 644 645 cell_1rw
* cell instance $8485 m0 *1 2.115,46.41
X$8485 71 34 72 644 645 cell_1rw
* cell instance $8486 m0 *1 2.82,46.41
X$8486 73 34 74 644 645 cell_1rw
* cell instance $8487 m0 *1 3.525,46.41
X$8487 75 34 76 644 645 cell_1rw
* cell instance $8488 m0 *1 4.23,46.41
X$8488 77 34 78 644 645 cell_1rw
* cell instance $8489 m0 *1 4.935,46.41
X$8489 79 34 80 644 645 cell_1rw
* cell instance $8490 m0 *1 5.64,46.41
X$8490 81 34 82 644 645 cell_1rw
* cell instance $8491 m0 *1 6.345,46.41
X$8491 83 34 84 644 645 cell_1rw
* cell instance $8492 m0 *1 7.05,46.41
X$8492 85 34 86 644 645 cell_1rw
* cell instance $8493 m0 *1 7.755,46.41
X$8493 87 34 88 644 645 cell_1rw
* cell instance $8494 m0 *1 8.46,46.41
X$8494 89 34 90 644 645 cell_1rw
* cell instance $8495 m0 *1 9.165,46.41
X$8495 91 34 92 644 645 cell_1rw
* cell instance $8496 m0 *1 9.87,46.41
X$8496 93 34 94 644 645 cell_1rw
* cell instance $8497 m0 *1 10.575,46.41
X$8497 95 34 96 644 645 cell_1rw
* cell instance $8498 m0 *1 11.28,46.41
X$8498 97 34 98 644 645 cell_1rw
* cell instance $8499 m0 *1 11.985,46.41
X$8499 99 34 100 644 645 cell_1rw
* cell instance $8500 m0 *1 12.69,46.41
X$8500 101 34 102 644 645 cell_1rw
* cell instance $8501 m0 *1 13.395,46.41
X$8501 103 34 104 644 645 cell_1rw
* cell instance $8502 m0 *1 14.1,46.41
X$8502 105 34 106 644 645 cell_1rw
* cell instance $8503 m0 *1 14.805,46.41
X$8503 107 34 108 644 645 cell_1rw
* cell instance $8504 m0 *1 15.51,46.41
X$8504 109 34 110 644 645 cell_1rw
* cell instance $8505 m0 *1 16.215,46.41
X$8505 111 34 112 644 645 cell_1rw
* cell instance $8506 m0 *1 16.92,46.41
X$8506 113 34 114 644 645 cell_1rw
* cell instance $8507 m0 *1 17.625,46.41
X$8507 115 34 116 644 645 cell_1rw
* cell instance $8508 m0 *1 18.33,46.41
X$8508 117 34 118 644 645 cell_1rw
* cell instance $8509 m0 *1 19.035,46.41
X$8509 119 34 120 644 645 cell_1rw
* cell instance $8510 m0 *1 19.74,46.41
X$8510 121 34 122 644 645 cell_1rw
* cell instance $8511 m0 *1 20.445,46.41
X$8511 123 34 124 644 645 cell_1rw
* cell instance $8512 m0 *1 21.15,46.41
X$8512 125 34 126 644 645 cell_1rw
* cell instance $8513 m0 *1 21.855,46.41
X$8513 127 34 128 644 645 cell_1rw
* cell instance $8514 m0 *1 22.56,46.41
X$8514 129 34 130 644 645 cell_1rw
* cell instance $8515 m0 *1 23.265,46.41
X$8515 131 34 132 644 645 cell_1rw
* cell instance $8516 m0 *1 23.97,46.41
X$8516 133 34 134 644 645 cell_1rw
* cell instance $8517 m0 *1 24.675,46.41
X$8517 135 34 136 644 645 cell_1rw
* cell instance $8518 m0 *1 25.38,46.41
X$8518 137 34 138 644 645 cell_1rw
* cell instance $8519 m0 *1 26.085,46.41
X$8519 139 34 140 644 645 cell_1rw
* cell instance $8520 m0 *1 26.79,46.41
X$8520 141 34 142 644 645 cell_1rw
* cell instance $8521 m0 *1 27.495,46.41
X$8521 143 34 144 644 645 cell_1rw
* cell instance $8522 m0 *1 28.2,46.41
X$8522 145 34 146 644 645 cell_1rw
* cell instance $8523 m0 *1 28.905,46.41
X$8523 147 34 148 644 645 cell_1rw
* cell instance $8524 m0 *1 29.61,46.41
X$8524 149 34 150 644 645 cell_1rw
* cell instance $8525 m0 *1 30.315,46.41
X$8525 151 34 152 644 645 cell_1rw
* cell instance $8526 m0 *1 31.02,46.41
X$8526 153 34 154 644 645 cell_1rw
* cell instance $8527 m0 *1 31.725,46.41
X$8527 155 34 156 644 645 cell_1rw
* cell instance $8528 m0 *1 32.43,46.41
X$8528 157 34 158 644 645 cell_1rw
* cell instance $8529 m0 *1 33.135,46.41
X$8529 159 34 160 644 645 cell_1rw
* cell instance $8530 m0 *1 33.84,46.41
X$8530 161 34 162 644 645 cell_1rw
* cell instance $8531 m0 *1 34.545,46.41
X$8531 163 34 164 644 645 cell_1rw
* cell instance $8532 m0 *1 35.25,46.41
X$8532 165 34 166 644 645 cell_1rw
* cell instance $8533 m0 *1 35.955,46.41
X$8533 167 34 168 644 645 cell_1rw
* cell instance $8534 m0 *1 36.66,46.41
X$8534 169 34 170 644 645 cell_1rw
* cell instance $8535 m0 *1 37.365,46.41
X$8535 171 34 172 644 645 cell_1rw
* cell instance $8536 m0 *1 38.07,46.41
X$8536 173 34 174 644 645 cell_1rw
* cell instance $8537 m0 *1 38.775,46.41
X$8537 175 34 176 644 645 cell_1rw
* cell instance $8538 m0 *1 39.48,46.41
X$8538 177 34 178 644 645 cell_1rw
* cell instance $8539 m0 *1 40.185,46.41
X$8539 179 34 180 644 645 cell_1rw
* cell instance $8540 m0 *1 40.89,46.41
X$8540 181 34 182 644 645 cell_1rw
* cell instance $8541 m0 *1 41.595,46.41
X$8541 183 34 184 644 645 cell_1rw
* cell instance $8542 m0 *1 42.3,46.41
X$8542 185 34 186 644 645 cell_1rw
* cell instance $8543 m0 *1 43.005,46.41
X$8543 187 34 188 644 645 cell_1rw
* cell instance $8544 m0 *1 43.71,46.41
X$8544 189 34 190 644 645 cell_1rw
* cell instance $8545 m0 *1 44.415,46.41
X$8545 191 34 192 644 645 cell_1rw
* cell instance $8546 m0 *1 45.12,46.41
X$8546 193 34 194 644 645 cell_1rw
* cell instance $8547 m0 *1 45.825,46.41
X$8547 195 34 196 644 645 cell_1rw
* cell instance $8548 m0 *1 46.53,46.41
X$8548 197 34 198 644 645 cell_1rw
* cell instance $8549 m0 *1 47.235,46.41
X$8549 199 34 200 644 645 cell_1rw
* cell instance $8550 m0 *1 47.94,46.41
X$8550 201 34 202 644 645 cell_1rw
* cell instance $8551 m0 *1 48.645,46.41
X$8551 203 34 204 644 645 cell_1rw
* cell instance $8552 m0 *1 49.35,46.41
X$8552 205 34 206 644 645 cell_1rw
* cell instance $8553 m0 *1 50.055,46.41
X$8553 207 34 208 644 645 cell_1rw
* cell instance $8554 m0 *1 50.76,46.41
X$8554 209 34 210 644 645 cell_1rw
* cell instance $8555 m0 *1 51.465,46.41
X$8555 211 34 212 644 645 cell_1rw
* cell instance $8556 m0 *1 52.17,46.41
X$8556 213 34 214 644 645 cell_1rw
* cell instance $8557 m0 *1 52.875,46.41
X$8557 215 34 216 644 645 cell_1rw
* cell instance $8558 m0 *1 53.58,46.41
X$8558 217 34 218 644 645 cell_1rw
* cell instance $8559 m0 *1 54.285,46.41
X$8559 219 34 220 644 645 cell_1rw
* cell instance $8560 m0 *1 54.99,46.41
X$8560 221 34 222 644 645 cell_1rw
* cell instance $8561 m0 *1 55.695,46.41
X$8561 223 34 224 644 645 cell_1rw
* cell instance $8562 m0 *1 56.4,46.41
X$8562 225 34 226 644 645 cell_1rw
* cell instance $8563 m0 *1 57.105,46.41
X$8563 227 34 228 644 645 cell_1rw
* cell instance $8564 m0 *1 57.81,46.41
X$8564 229 34 230 644 645 cell_1rw
* cell instance $8565 m0 *1 58.515,46.41
X$8565 231 34 232 644 645 cell_1rw
* cell instance $8566 m0 *1 59.22,46.41
X$8566 233 34 234 644 645 cell_1rw
* cell instance $8567 m0 *1 59.925,46.41
X$8567 235 34 236 644 645 cell_1rw
* cell instance $8568 m0 *1 60.63,46.41
X$8568 237 34 238 644 645 cell_1rw
* cell instance $8569 m0 *1 61.335,46.41
X$8569 239 34 240 644 645 cell_1rw
* cell instance $8570 m0 *1 62.04,46.41
X$8570 241 34 242 644 645 cell_1rw
* cell instance $8571 m0 *1 62.745,46.41
X$8571 243 34 244 644 645 cell_1rw
* cell instance $8572 m0 *1 63.45,46.41
X$8572 245 34 246 644 645 cell_1rw
* cell instance $8573 m0 *1 64.155,46.41
X$8573 247 34 248 644 645 cell_1rw
* cell instance $8574 m0 *1 64.86,46.41
X$8574 249 34 250 644 645 cell_1rw
* cell instance $8575 m0 *1 65.565,46.41
X$8575 251 34 252 644 645 cell_1rw
* cell instance $8576 m0 *1 66.27,46.41
X$8576 253 34 254 644 645 cell_1rw
* cell instance $8577 m0 *1 66.975,46.41
X$8577 255 34 256 644 645 cell_1rw
* cell instance $8578 m0 *1 67.68,46.41
X$8578 257 34 258 644 645 cell_1rw
* cell instance $8579 m0 *1 68.385,46.41
X$8579 259 34 260 644 645 cell_1rw
* cell instance $8580 m0 *1 69.09,46.41
X$8580 261 34 262 644 645 cell_1rw
* cell instance $8581 m0 *1 69.795,46.41
X$8581 263 34 264 644 645 cell_1rw
* cell instance $8582 m0 *1 70.5,46.41
X$8582 265 34 266 644 645 cell_1rw
* cell instance $8583 m0 *1 71.205,46.41
X$8583 267 34 268 644 645 cell_1rw
* cell instance $8584 m0 *1 71.91,46.41
X$8584 269 34 270 644 645 cell_1rw
* cell instance $8585 m0 *1 72.615,46.41
X$8585 271 34 272 644 645 cell_1rw
* cell instance $8586 m0 *1 73.32,46.41
X$8586 273 34 274 644 645 cell_1rw
* cell instance $8587 m0 *1 74.025,46.41
X$8587 275 34 276 644 645 cell_1rw
* cell instance $8588 m0 *1 74.73,46.41
X$8588 277 34 278 644 645 cell_1rw
* cell instance $8589 m0 *1 75.435,46.41
X$8589 279 34 280 644 645 cell_1rw
* cell instance $8590 m0 *1 76.14,46.41
X$8590 281 34 282 644 645 cell_1rw
* cell instance $8591 m0 *1 76.845,46.41
X$8591 283 34 284 644 645 cell_1rw
* cell instance $8592 m0 *1 77.55,46.41
X$8592 285 34 286 644 645 cell_1rw
* cell instance $8593 m0 *1 78.255,46.41
X$8593 287 34 288 644 645 cell_1rw
* cell instance $8594 m0 *1 78.96,46.41
X$8594 289 34 290 644 645 cell_1rw
* cell instance $8595 m0 *1 79.665,46.41
X$8595 291 34 292 644 645 cell_1rw
* cell instance $8596 m0 *1 80.37,46.41
X$8596 293 34 294 644 645 cell_1rw
* cell instance $8597 m0 *1 81.075,46.41
X$8597 295 34 296 644 645 cell_1rw
* cell instance $8598 m0 *1 81.78,46.41
X$8598 297 34 298 644 645 cell_1rw
* cell instance $8599 m0 *1 82.485,46.41
X$8599 299 34 300 644 645 cell_1rw
* cell instance $8600 m0 *1 83.19,46.41
X$8600 301 34 302 644 645 cell_1rw
* cell instance $8601 m0 *1 83.895,46.41
X$8601 303 34 304 644 645 cell_1rw
* cell instance $8602 m0 *1 84.6,46.41
X$8602 305 34 306 644 645 cell_1rw
* cell instance $8603 m0 *1 85.305,46.41
X$8603 307 34 308 644 645 cell_1rw
* cell instance $8604 m0 *1 86.01,46.41
X$8604 309 34 310 644 645 cell_1rw
* cell instance $8605 m0 *1 86.715,46.41
X$8605 311 34 312 644 645 cell_1rw
* cell instance $8606 m0 *1 87.42,46.41
X$8606 313 34 314 644 645 cell_1rw
* cell instance $8607 m0 *1 88.125,46.41
X$8607 315 34 316 644 645 cell_1rw
* cell instance $8608 m0 *1 88.83,46.41
X$8608 317 34 318 644 645 cell_1rw
* cell instance $8609 m0 *1 89.535,46.41
X$8609 319 34 320 644 645 cell_1rw
* cell instance $8610 m0 *1 90.24,46.41
X$8610 321 34 323 644 645 cell_1rw
* cell instance $8611 m0 *1 90.945,46.41
X$8611 324 34 325 644 645 cell_1rw
* cell instance $8612 m0 *1 91.65,46.41
X$8612 326 34 327 644 645 cell_1rw
* cell instance $8613 m0 *1 92.355,46.41
X$8613 328 34 329 644 645 cell_1rw
* cell instance $8614 m0 *1 93.06,46.41
X$8614 330 34 331 644 645 cell_1rw
* cell instance $8615 m0 *1 93.765,46.41
X$8615 332 34 333 644 645 cell_1rw
* cell instance $8616 m0 *1 94.47,46.41
X$8616 334 34 335 644 645 cell_1rw
* cell instance $8617 m0 *1 95.175,46.41
X$8617 336 34 337 644 645 cell_1rw
* cell instance $8618 m0 *1 95.88,46.41
X$8618 338 34 339 644 645 cell_1rw
* cell instance $8619 m0 *1 96.585,46.41
X$8619 340 34 341 644 645 cell_1rw
* cell instance $8620 m0 *1 97.29,46.41
X$8620 342 34 343 644 645 cell_1rw
* cell instance $8621 m0 *1 97.995,46.41
X$8621 344 34 345 644 645 cell_1rw
* cell instance $8622 m0 *1 98.7,46.41
X$8622 346 34 347 644 645 cell_1rw
* cell instance $8623 m0 *1 99.405,46.41
X$8623 348 34 349 644 645 cell_1rw
* cell instance $8624 m0 *1 100.11,46.41
X$8624 350 34 351 644 645 cell_1rw
* cell instance $8625 m0 *1 100.815,46.41
X$8625 352 34 353 644 645 cell_1rw
* cell instance $8626 m0 *1 101.52,46.41
X$8626 354 34 355 644 645 cell_1rw
* cell instance $8627 m0 *1 102.225,46.41
X$8627 356 34 357 644 645 cell_1rw
* cell instance $8628 m0 *1 102.93,46.41
X$8628 358 34 359 644 645 cell_1rw
* cell instance $8629 m0 *1 103.635,46.41
X$8629 360 34 361 644 645 cell_1rw
* cell instance $8630 m0 *1 104.34,46.41
X$8630 362 34 363 644 645 cell_1rw
* cell instance $8631 m0 *1 105.045,46.41
X$8631 364 34 365 644 645 cell_1rw
* cell instance $8632 m0 *1 105.75,46.41
X$8632 366 34 367 644 645 cell_1rw
* cell instance $8633 m0 *1 106.455,46.41
X$8633 368 34 369 644 645 cell_1rw
* cell instance $8634 m0 *1 107.16,46.41
X$8634 370 34 371 644 645 cell_1rw
* cell instance $8635 m0 *1 107.865,46.41
X$8635 372 34 373 644 645 cell_1rw
* cell instance $8636 m0 *1 108.57,46.41
X$8636 374 34 375 644 645 cell_1rw
* cell instance $8637 m0 *1 109.275,46.41
X$8637 376 34 377 644 645 cell_1rw
* cell instance $8638 m0 *1 109.98,46.41
X$8638 378 34 379 644 645 cell_1rw
* cell instance $8639 m0 *1 110.685,46.41
X$8639 380 34 381 644 645 cell_1rw
* cell instance $8640 m0 *1 111.39,46.41
X$8640 382 34 383 644 645 cell_1rw
* cell instance $8641 m0 *1 112.095,46.41
X$8641 384 34 385 644 645 cell_1rw
* cell instance $8642 m0 *1 112.8,46.41
X$8642 386 34 387 644 645 cell_1rw
* cell instance $8643 m0 *1 113.505,46.41
X$8643 388 34 389 644 645 cell_1rw
* cell instance $8644 m0 *1 114.21,46.41
X$8644 390 34 391 644 645 cell_1rw
* cell instance $8645 m0 *1 114.915,46.41
X$8645 392 34 393 644 645 cell_1rw
* cell instance $8646 m0 *1 115.62,46.41
X$8646 394 34 395 644 645 cell_1rw
* cell instance $8647 m0 *1 116.325,46.41
X$8647 396 34 397 644 645 cell_1rw
* cell instance $8648 m0 *1 117.03,46.41
X$8648 398 34 399 644 645 cell_1rw
* cell instance $8649 m0 *1 117.735,46.41
X$8649 400 34 401 644 645 cell_1rw
* cell instance $8650 m0 *1 118.44,46.41
X$8650 402 34 403 644 645 cell_1rw
* cell instance $8651 m0 *1 119.145,46.41
X$8651 404 34 405 644 645 cell_1rw
* cell instance $8652 m0 *1 119.85,46.41
X$8652 406 34 407 644 645 cell_1rw
* cell instance $8653 m0 *1 120.555,46.41
X$8653 408 34 409 644 645 cell_1rw
* cell instance $8654 m0 *1 121.26,46.41
X$8654 410 34 411 644 645 cell_1rw
* cell instance $8655 m0 *1 121.965,46.41
X$8655 412 34 413 644 645 cell_1rw
* cell instance $8656 m0 *1 122.67,46.41
X$8656 414 34 415 644 645 cell_1rw
* cell instance $8657 m0 *1 123.375,46.41
X$8657 416 34 417 644 645 cell_1rw
* cell instance $8658 m0 *1 124.08,46.41
X$8658 418 34 419 644 645 cell_1rw
* cell instance $8659 m0 *1 124.785,46.41
X$8659 420 34 421 644 645 cell_1rw
* cell instance $8660 m0 *1 125.49,46.41
X$8660 422 34 423 644 645 cell_1rw
* cell instance $8661 m0 *1 126.195,46.41
X$8661 424 34 425 644 645 cell_1rw
* cell instance $8662 m0 *1 126.9,46.41
X$8662 426 34 427 644 645 cell_1rw
* cell instance $8663 m0 *1 127.605,46.41
X$8663 428 34 429 644 645 cell_1rw
* cell instance $8664 m0 *1 128.31,46.41
X$8664 430 34 431 644 645 cell_1rw
* cell instance $8665 m0 *1 129.015,46.41
X$8665 432 34 433 644 645 cell_1rw
* cell instance $8666 m0 *1 129.72,46.41
X$8666 434 34 435 644 645 cell_1rw
* cell instance $8667 m0 *1 130.425,46.41
X$8667 436 34 437 644 645 cell_1rw
* cell instance $8668 m0 *1 131.13,46.41
X$8668 438 34 439 644 645 cell_1rw
* cell instance $8669 m0 *1 131.835,46.41
X$8669 440 34 441 644 645 cell_1rw
* cell instance $8670 m0 *1 132.54,46.41
X$8670 442 34 443 644 645 cell_1rw
* cell instance $8671 m0 *1 133.245,46.41
X$8671 444 34 445 644 645 cell_1rw
* cell instance $8672 m0 *1 133.95,46.41
X$8672 446 34 447 644 645 cell_1rw
* cell instance $8673 m0 *1 134.655,46.41
X$8673 448 34 449 644 645 cell_1rw
* cell instance $8674 m0 *1 135.36,46.41
X$8674 450 34 451 644 645 cell_1rw
* cell instance $8675 m0 *1 136.065,46.41
X$8675 452 34 453 644 645 cell_1rw
* cell instance $8676 m0 *1 136.77,46.41
X$8676 454 34 455 644 645 cell_1rw
* cell instance $8677 m0 *1 137.475,46.41
X$8677 456 34 457 644 645 cell_1rw
* cell instance $8678 m0 *1 138.18,46.41
X$8678 458 34 459 644 645 cell_1rw
* cell instance $8679 m0 *1 138.885,46.41
X$8679 460 34 461 644 645 cell_1rw
* cell instance $8680 m0 *1 139.59,46.41
X$8680 462 34 463 644 645 cell_1rw
* cell instance $8681 m0 *1 140.295,46.41
X$8681 464 34 465 644 645 cell_1rw
* cell instance $8682 m0 *1 141,46.41
X$8682 466 34 467 644 645 cell_1rw
* cell instance $8683 m0 *1 141.705,46.41
X$8683 468 34 469 644 645 cell_1rw
* cell instance $8684 m0 *1 142.41,46.41
X$8684 470 34 471 644 645 cell_1rw
* cell instance $8685 m0 *1 143.115,46.41
X$8685 472 34 473 644 645 cell_1rw
* cell instance $8686 m0 *1 143.82,46.41
X$8686 474 34 475 644 645 cell_1rw
* cell instance $8687 m0 *1 144.525,46.41
X$8687 476 34 477 644 645 cell_1rw
* cell instance $8688 m0 *1 145.23,46.41
X$8688 478 34 479 644 645 cell_1rw
* cell instance $8689 m0 *1 145.935,46.41
X$8689 480 34 481 644 645 cell_1rw
* cell instance $8690 m0 *1 146.64,46.41
X$8690 482 34 483 644 645 cell_1rw
* cell instance $8691 m0 *1 147.345,46.41
X$8691 484 34 485 644 645 cell_1rw
* cell instance $8692 m0 *1 148.05,46.41
X$8692 486 34 487 644 645 cell_1rw
* cell instance $8693 m0 *1 148.755,46.41
X$8693 488 34 489 644 645 cell_1rw
* cell instance $8694 m0 *1 149.46,46.41
X$8694 490 34 491 644 645 cell_1rw
* cell instance $8695 m0 *1 150.165,46.41
X$8695 492 34 493 644 645 cell_1rw
* cell instance $8696 m0 *1 150.87,46.41
X$8696 494 34 495 644 645 cell_1rw
* cell instance $8697 m0 *1 151.575,46.41
X$8697 496 34 497 644 645 cell_1rw
* cell instance $8698 m0 *1 152.28,46.41
X$8698 498 34 499 644 645 cell_1rw
* cell instance $8699 m0 *1 152.985,46.41
X$8699 500 34 501 644 645 cell_1rw
* cell instance $8700 m0 *1 153.69,46.41
X$8700 502 34 503 644 645 cell_1rw
* cell instance $8701 m0 *1 154.395,46.41
X$8701 504 34 505 644 645 cell_1rw
* cell instance $8702 m0 *1 155.1,46.41
X$8702 506 34 507 644 645 cell_1rw
* cell instance $8703 m0 *1 155.805,46.41
X$8703 508 34 509 644 645 cell_1rw
* cell instance $8704 m0 *1 156.51,46.41
X$8704 510 34 511 644 645 cell_1rw
* cell instance $8705 m0 *1 157.215,46.41
X$8705 512 34 513 644 645 cell_1rw
* cell instance $8706 m0 *1 157.92,46.41
X$8706 514 34 515 644 645 cell_1rw
* cell instance $8707 m0 *1 158.625,46.41
X$8707 516 34 517 644 645 cell_1rw
* cell instance $8708 m0 *1 159.33,46.41
X$8708 518 34 519 644 645 cell_1rw
* cell instance $8709 m0 *1 160.035,46.41
X$8709 520 34 521 644 645 cell_1rw
* cell instance $8710 m0 *1 160.74,46.41
X$8710 522 34 523 644 645 cell_1rw
* cell instance $8711 m0 *1 161.445,46.41
X$8711 524 34 525 644 645 cell_1rw
* cell instance $8712 m0 *1 162.15,46.41
X$8712 526 34 527 644 645 cell_1rw
* cell instance $8713 m0 *1 162.855,46.41
X$8713 528 34 529 644 645 cell_1rw
* cell instance $8714 m0 *1 163.56,46.41
X$8714 530 34 531 644 645 cell_1rw
* cell instance $8715 m0 *1 164.265,46.41
X$8715 532 34 533 644 645 cell_1rw
* cell instance $8716 m0 *1 164.97,46.41
X$8716 534 34 535 644 645 cell_1rw
* cell instance $8717 m0 *1 165.675,46.41
X$8717 536 34 537 644 645 cell_1rw
* cell instance $8718 m0 *1 166.38,46.41
X$8718 538 34 539 644 645 cell_1rw
* cell instance $8719 m0 *1 167.085,46.41
X$8719 540 34 541 644 645 cell_1rw
* cell instance $8720 m0 *1 167.79,46.41
X$8720 542 34 543 644 645 cell_1rw
* cell instance $8721 m0 *1 168.495,46.41
X$8721 544 34 545 644 645 cell_1rw
* cell instance $8722 m0 *1 169.2,46.41
X$8722 546 34 547 644 645 cell_1rw
* cell instance $8723 m0 *1 169.905,46.41
X$8723 548 34 549 644 645 cell_1rw
* cell instance $8724 m0 *1 170.61,46.41
X$8724 550 34 551 644 645 cell_1rw
* cell instance $8725 m0 *1 171.315,46.41
X$8725 552 34 553 644 645 cell_1rw
* cell instance $8726 m0 *1 172.02,46.41
X$8726 554 34 555 644 645 cell_1rw
* cell instance $8727 m0 *1 172.725,46.41
X$8727 556 34 557 644 645 cell_1rw
* cell instance $8728 m0 *1 173.43,46.41
X$8728 558 34 559 644 645 cell_1rw
* cell instance $8729 m0 *1 174.135,46.41
X$8729 560 34 561 644 645 cell_1rw
* cell instance $8730 m0 *1 174.84,46.41
X$8730 562 34 563 644 645 cell_1rw
* cell instance $8731 m0 *1 175.545,46.41
X$8731 564 34 565 644 645 cell_1rw
* cell instance $8732 m0 *1 176.25,46.41
X$8732 566 34 567 644 645 cell_1rw
* cell instance $8733 m0 *1 176.955,46.41
X$8733 568 34 569 644 645 cell_1rw
* cell instance $8734 m0 *1 177.66,46.41
X$8734 570 34 571 644 645 cell_1rw
* cell instance $8735 m0 *1 178.365,46.41
X$8735 572 34 573 644 645 cell_1rw
* cell instance $8736 m0 *1 179.07,46.41
X$8736 574 34 575 644 645 cell_1rw
* cell instance $8737 m0 *1 179.775,46.41
X$8737 576 34 577 644 645 cell_1rw
* cell instance $8738 m0 *1 180.48,46.41
X$8738 578 34 579 644 645 cell_1rw
* cell instance $8739 r0 *1 0.705,46.41
X$8739 67 35 68 644 645 cell_1rw
* cell instance $8740 r0 *1 0,46.41
X$8740 65 35 66 644 645 cell_1rw
* cell instance $8741 r0 *1 1.41,46.41
X$8741 69 35 70 644 645 cell_1rw
* cell instance $8742 r0 *1 2.115,46.41
X$8742 71 35 72 644 645 cell_1rw
* cell instance $8743 r0 *1 2.82,46.41
X$8743 73 35 74 644 645 cell_1rw
* cell instance $8744 r0 *1 3.525,46.41
X$8744 75 35 76 644 645 cell_1rw
* cell instance $8745 r0 *1 4.23,46.41
X$8745 77 35 78 644 645 cell_1rw
* cell instance $8746 r0 *1 4.935,46.41
X$8746 79 35 80 644 645 cell_1rw
* cell instance $8747 r0 *1 5.64,46.41
X$8747 81 35 82 644 645 cell_1rw
* cell instance $8748 r0 *1 6.345,46.41
X$8748 83 35 84 644 645 cell_1rw
* cell instance $8749 r0 *1 7.05,46.41
X$8749 85 35 86 644 645 cell_1rw
* cell instance $8750 r0 *1 7.755,46.41
X$8750 87 35 88 644 645 cell_1rw
* cell instance $8751 r0 *1 8.46,46.41
X$8751 89 35 90 644 645 cell_1rw
* cell instance $8752 r0 *1 9.165,46.41
X$8752 91 35 92 644 645 cell_1rw
* cell instance $8753 r0 *1 9.87,46.41
X$8753 93 35 94 644 645 cell_1rw
* cell instance $8754 r0 *1 10.575,46.41
X$8754 95 35 96 644 645 cell_1rw
* cell instance $8755 r0 *1 11.28,46.41
X$8755 97 35 98 644 645 cell_1rw
* cell instance $8756 r0 *1 11.985,46.41
X$8756 99 35 100 644 645 cell_1rw
* cell instance $8757 r0 *1 12.69,46.41
X$8757 101 35 102 644 645 cell_1rw
* cell instance $8758 r0 *1 13.395,46.41
X$8758 103 35 104 644 645 cell_1rw
* cell instance $8759 r0 *1 14.1,46.41
X$8759 105 35 106 644 645 cell_1rw
* cell instance $8760 r0 *1 14.805,46.41
X$8760 107 35 108 644 645 cell_1rw
* cell instance $8761 r0 *1 15.51,46.41
X$8761 109 35 110 644 645 cell_1rw
* cell instance $8762 r0 *1 16.215,46.41
X$8762 111 35 112 644 645 cell_1rw
* cell instance $8763 r0 *1 16.92,46.41
X$8763 113 35 114 644 645 cell_1rw
* cell instance $8764 r0 *1 17.625,46.41
X$8764 115 35 116 644 645 cell_1rw
* cell instance $8765 r0 *1 18.33,46.41
X$8765 117 35 118 644 645 cell_1rw
* cell instance $8766 r0 *1 19.035,46.41
X$8766 119 35 120 644 645 cell_1rw
* cell instance $8767 r0 *1 19.74,46.41
X$8767 121 35 122 644 645 cell_1rw
* cell instance $8768 r0 *1 20.445,46.41
X$8768 123 35 124 644 645 cell_1rw
* cell instance $8769 r0 *1 21.15,46.41
X$8769 125 35 126 644 645 cell_1rw
* cell instance $8770 r0 *1 21.855,46.41
X$8770 127 35 128 644 645 cell_1rw
* cell instance $8771 r0 *1 22.56,46.41
X$8771 129 35 130 644 645 cell_1rw
* cell instance $8772 r0 *1 23.265,46.41
X$8772 131 35 132 644 645 cell_1rw
* cell instance $8773 r0 *1 23.97,46.41
X$8773 133 35 134 644 645 cell_1rw
* cell instance $8774 r0 *1 24.675,46.41
X$8774 135 35 136 644 645 cell_1rw
* cell instance $8775 r0 *1 25.38,46.41
X$8775 137 35 138 644 645 cell_1rw
* cell instance $8776 r0 *1 26.085,46.41
X$8776 139 35 140 644 645 cell_1rw
* cell instance $8777 r0 *1 26.79,46.41
X$8777 141 35 142 644 645 cell_1rw
* cell instance $8778 r0 *1 27.495,46.41
X$8778 143 35 144 644 645 cell_1rw
* cell instance $8779 r0 *1 28.2,46.41
X$8779 145 35 146 644 645 cell_1rw
* cell instance $8780 r0 *1 28.905,46.41
X$8780 147 35 148 644 645 cell_1rw
* cell instance $8781 r0 *1 29.61,46.41
X$8781 149 35 150 644 645 cell_1rw
* cell instance $8782 r0 *1 30.315,46.41
X$8782 151 35 152 644 645 cell_1rw
* cell instance $8783 r0 *1 31.02,46.41
X$8783 153 35 154 644 645 cell_1rw
* cell instance $8784 r0 *1 31.725,46.41
X$8784 155 35 156 644 645 cell_1rw
* cell instance $8785 r0 *1 32.43,46.41
X$8785 157 35 158 644 645 cell_1rw
* cell instance $8786 r0 *1 33.135,46.41
X$8786 159 35 160 644 645 cell_1rw
* cell instance $8787 r0 *1 33.84,46.41
X$8787 161 35 162 644 645 cell_1rw
* cell instance $8788 r0 *1 34.545,46.41
X$8788 163 35 164 644 645 cell_1rw
* cell instance $8789 r0 *1 35.25,46.41
X$8789 165 35 166 644 645 cell_1rw
* cell instance $8790 r0 *1 35.955,46.41
X$8790 167 35 168 644 645 cell_1rw
* cell instance $8791 r0 *1 36.66,46.41
X$8791 169 35 170 644 645 cell_1rw
* cell instance $8792 r0 *1 37.365,46.41
X$8792 171 35 172 644 645 cell_1rw
* cell instance $8793 r0 *1 38.07,46.41
X$8793 173 35 174 644 645 cell_1rw
* cell instance $8794 r0 *1 38.775,46.41
X$8794 175 35 176 644 645 cell_1rw
* cell instance $8795 r0 *1 39.48,46.41
X$8795 177 35 178 644 645 cell_1rw
* cell instance $8796 r0 *1 40.185,46.41
X$8796 179 35 180 644 645 cell_1rw
* cell instance $8797 r0 *1 40.89,46.41
X$8797 181 35 182 644 645 cell_1rw
* cell instance $8798 r0 *1 41.595,46.41
X$8798 183 35 184 644 645 cell_1rw
* cell instance $8799 r0 *1 42.3,46.41
X$8799 185 35 186 644 645 cell_1rw
* cell instance $8800 r0 *1 43.005,46.41
X$8800 187 35 188 644 645 cell_1rw
* cell instance $8801 r0 *1 43.71,46.41
X$8801 189 35 190 644 645 cell_1rw
* cell instance $8802 r0 *1 44.415,46.41
X$8802 191 35 192 644 645 cell_1rw
* cell instance $8803 r0 *1 45.12,46.41
X$8803 193 35 194 644 645 cell_1rw
* cell instance $8804 r0 *1 45.825,46.41
X$8804 195 35 196 644 645 cell_1rw
* cell instance $8805 r0 *1 46.53,46.41
X$8805 197 35 198 644 645 cell_1rw
* cell instance $8806 r0 *1 47.235,46.41
X$8806 199 35 200 644 645 cell_1rw
* cell instance $8807 r0 *1 47.94,46.41
X$8807 201 35 202 644 645 cell_1rw
* cell instance $8808 r0 *1 48.645,46.41
X$8808 203 35 204 644 645 cell_1rw
* cell instance $8809 r0 *1 49.35,46.41
X$8809 205 35 206 644 645 cell_1rw
* cell instance $8810 r0 *1 50.055,46.41
X$8810 207 35 208 644 645 cell_1rw
* cell instance $8811 r0 *1 50.76,46.41
X$8811 209 35 210 644 645 cell_1rw
* cell instance $8812 r0 *1 51.465,46.41
X$8812 211 35 212 644 645 cell_1rw
* cell instance $8813 r0 *1 52.17,46.41
X$8813 213 35 214 644 645 cell_1rw
* cell instance $8814 r0 *1 52.875,46.41
X$8814 215 35 216 644 645 cell_1rw
* cell instance $8815 r0 *1 53.58,46.41
X$8815 217 35 218 644 645 cell_1rw
* cell instance $8816 r0 *1 54.285,46.41
X$8816 219 35 220 644 645 cell_1rw
* cell instance $8817 r0 *1 54.99,46.41
X$8817 221 35 222 644 645 cell_1rw
* cell instance $8818 r0 *1 55.695,46.41
X$8818 223 35 224 644 645 cell_1rw
* cell instance $8819 r0 *1 56.4,46.41
X$8819 225 35 226 644 645 cell_1rw
* cell instance $8820 r0 *1 57.105,46.41
X$8820 227 35 228 644 645 cell_1rw
* cell instance $8821 r0 *1 57.81,46.41
X$8821 229 35 230 644 645 cell_1rw
* cell instance $8822 r0 *1 58.515,46.41
X$8822 231 35 232 644 645 cell_1rw
* cell instance $8823 r0 *1 59.22,46.41
X$8823 233 35 234 644 645 cell_1rw
* cell instance $8824 r0 *1 59.925,46.41
X$8824 235 35 236 644 645 cell_1rw
* cell instance $8825 r0 *1 60.63,46.41
X$8825 237 35 238 644 645 cell_1rw
* cell instance $8826 r0 *1 61.335,46.41
X$8826 239 35 240 644 645 cell_1rw
* cell instance $8827 r0 *1 62.04,46.41
X$8827 241 35 242 644 645 cell_1rw
* cell instance $8828 r0 *1 62.745,46.41
X$8828 243 35 244 644 645 cell_1rw
* cell instance $8829 r0 *1 63.45,46.41
X$8829 245 35 246 644 645 cell_1rw
* cell instance $8830 r0 *1 64.155,46.41
X$8830 247 35 248 644 645 cell_1rw
* cell instance $8831 r0 *1 64.86,46.41
X$8831 249 35 250 644 645 cell_1rw
* cell instance $8832 r0 *1 65.565,46.41
X$8832 251 35 252 644 645 cell_1rw
* cell instance $8833 r0 *1 66.27,46.41
X$8833 253 35 254 644 645 cell_1rw
* cell instance $8834 r0 *1 66.975,46.41
X$8834 255 35 256 644 645 cell_1rw
* cell instance $8835 r0 *1 67.68,46.41
X$8835 257 35 258 644 645 cell_1rw
* cell instance $8836 r0 *1 68.385,46.41
X$8836 259 35 260 644 645 cell_1rw
* cell instance $8837 r0 *1 69.09,46.41
X$8837 261 35 262 644 645 cell_1rw
* cell instance $8838 r0 *1 69.795,46.41
X$8838 263 35 264 644 645 cell_1rw
* cell instance $8839 r0 *1 70.5,46.41
X$8839 265 35 266 644 645 cell_1rw
* cell instance $8840 r0 *1 71.205,46.41
X$8840 267 35 268 644 645 cell_1rw
* cell instance $8841 r0 *1 71.91,46.41
X$8841 269 35 270 644 645 cell_1rw
* cell instance $8842 r0 *1 72.615,46.41
X$8842 271 35 272 644 645 cell_1rw
* cell instance $8843 r0 *1 73.32,46.41
X$8843 273 35 274 644 645 cell_1rw
* cell instance $8844 r0 *1 74.025,46.41
X$8844 275 35 276 644 645 cell_1rw
* cell instance $8845 r0 *1 74.73,46.41
X$8845 277 35 278 644 645 cell_1rw
* cell instance $8846 r0 *1 75.435,46.41
X$8846 279 35 280 644 645 cell_1rw
* cell instance $8847 r0 *1 76.14,46.41
X$8847 281 35 282 644 645 cell_1rw
* cell instance $8848 r0 *1 76.845,46.41
X$8848 283 35 284 644 645 cell_1rw
* cell instance $8849 r0 *1 77.55,46.41
X$8849 285 35 286 644 645 cell_1rw
* cell instance $8850 r0 *1 78.255,46.41
X$8850 287 35 288 644 645 cell_1rw
* cell instance $8851 r0 *1 78.96,46.41
X$8851 289 35 290 644 645 cell_1rw
* cell instance $8852 r0 *1 79.665,46.41
X$8852 291 35 292 644 645 cell_1rw
* cell instance $8853 r0 *1 80.37,46.41
X$8853 293 35 294 644 645 cell_1rw
* cell instance $8854 r0 *1 81.075,46.41
X$8854 295 35 296 644 645 cell_1rw
* cell instance $8855 r0 *1 81.78,46.41
X$8855 297 35 298 644 645 cell_1rw
* cell instance $8856 r0 *1 82.485,46.41
X$8856 299 35 300 644 645 cell_1rw
* cell instance $8857 r0 *1 83.19,46.41
X$8857 301 35 302 644 645 cell_1rw
* cell instance $8858 r0 *1 83.895,46.41
X$8858 303 35 304 644 645 cell_1rw
* cell instance $8859 r0 *1 84.6,46.41
X$8859 305 35 306 644 645 cell_1rw
* cell instance $8860 r0 *1 85.305,46.41
X$8860 307 35 308 644 645 cell_1rw
* cell instance $8861 r0 *1 86.01,46.41
X$8861 309 35 310 644 645 cell_1rw
* cell instance $8862 r0 *1 86.715,46.41
X$8862 311 35 312 644 645 cell_1rw
* cell instance $8863 r0 *1 87.42,46.41
X$8863 313 35 314 644 645 cell_1rw
* cell instance $8864 r0 *1 88.125,46.41
X$8864 315 35 316 644 645 cell_1rw
* cell instance $8865 r0 *1 88.83,46.41
X$8865 317 35 318 644 645 cell_1rw
* cell instance $8866 r0 *1 89.535,46.41
X$8866 319 35 320 644 645 cell_1rw
* cell instance $8867 r0 *1 90.24,46.41
X$8867 321 35 323 644 645 cell_1rw
* cell instance $8868 r0 *1 90.945,46.41
X$8868 324 35 325 644 645 cell_1rw
* cell instance $8869 r0 *1 91.65,46.41
X$8869 326 35 327 644 645 cell_1rw
* cell instance $8870 r0 *1 92.355,46.41
X$8870 328 35 329 644 645 cell_1rw
* cell instance $8871 r0 *1 93.06,46.41
X$8871 330 35 331 644 645 cell_1rw
* cell instance $8872 r0 *1 93.765,46.41
X$8872 332 35 333 644 645 cell_1rw
* cell instance $8873 r0 *1 94.47,46.41
X$8873 334 35 335 644 645 cell_1rw
* cell instance $8874 r0 *1 95.175,46.41
X$8874 336 35 337 644 645 cell_1rw
* cell instance $8875 r0 *1 95.88,46.41
X$8875 338 35 339 644 645 cell_1rw
* cell instance $8876 r0 *1 96.585,46.41
X$8876 340 35 341 644 645 cell_1rw
* cell instance $8877 r0 *1 97.29,46.41
X$8877 342 35 343 644 645 cell_1rw
* cell instance $8878 r0 *1 97.995,46.41
X$8878 344 35 345 644 645 cell_1rw
* cell instance $8879 r0 *1 98.7,46.41
X$8879 346 35 347 644 645 cell_1rw
* cell instance $8880 r0 *1 99.405,46.41
X$8880 348 35 349 644 645 cell_1rw
* cell instance $8881 r0 *1 100.11,46.41
X$8881 350 35 351 644 645 cell_1rw
* cell instance $8882 r0 *1 100.815,46.41
X$8882 352 35 353 644 645 cell_1rw
* cell instance $8883 r0 *1 101.52,46.41
X$8883 354 35 355 644 645 cell_1rw
* cell instance $8884 r0 *1 102.225,46.41
X$8884 356 35 357 644 645 cell_1rw
* cell instance $8885 r0 *1 102.93,46.41
X$8885 358 35 359 644 645 cell_1rw
* cell instance $8886 r0 *1 103.635,46.41
X$8886 360 35 361 644 645 cell_1rw
* cell instance $8887 r0 *1 104.34,46.41
X$8887 362 35 363 644 645 cell_1rw
* cell instance $8888 r0 *1 105.045,46.41
X$8888 364 35 365 644 645 cell_1rw
* cell instance $8889 r0 *1 105.75,46.41
X$8889 366 35 367 644 645 cell_1rw
* cell instance $8890 r0 *1 106.455,46.41
X$8890 368 35 369 644 645 cell_1rw
* cell instance $8891 r0 *1 107.16,46.41
X$8891 370 35 371 644 645 cell_1rw
* cell instance $8892 r0 *1 107.865,46.41
X$8892 372 35 373 644 645 cell_1rw
* cell instance $8893 r0 *1 108.57,46.41
X$8893 374 35 375 644 645 cell_1rw
* cell instance $8894 r0 *1 109.275,46.41
X$8894 376 35 377 644 645 cell_1rw
* cell instance $8895 r0 *1 109.98,46.41
X$8895 378 35 379 644 645 cell_1rw
* cell instance $8896 r0 *1 110.685,46.41
X$8896 380 35 381 644 645 cell_1rw
* cell instance $8897 r0 *1 111.39,46.41
X$8897 382 35 383 644 645 cell_1rw
* cell instance $8898 r0 *1 112.095,46.41
X$8898 384 35 385 644 645 cell_1rw
* cell instance $8899 r0 *1 112.8,46.41
X$8899 386 35 387 644 645 cell_1rw
* cell instance $8900 r0 *1 113.505,46.41
X$8900 388 35 389 644 645 cell_1rw
* cell instance $8901 r0 *1 114.21,46.41
X$8901 390 35 391 644 645 cell_1rw
* cell instance $8902 r0 *1 114.915,46.41
X$8902 392 35 393 644 645 cell_1rw
* cell instance $8903 r0 *1 115.62,46.41
X$8903 394 35 395 644 645 cell_1rw
* cell instance $8904 r0 *1 116.325,46.41
X$8904 396 35 397 644 645 cell_1rw
* cell instance $8905 r0 *1 117.03,46.41
X$8905 398 35 399 644 645 cell_1rw
* cell instance $8906 r0 *1 117.735,46.41
X$8906 400 35 401 644 645 cell_1rw
* cell instance $8907 r0 *1 118.44,46.41
X$8907 402 35 403 644 645 cell_1rw
* cell instance $8908 r0 *1 119.145,46.41
X$8908 404 35 405 644 645 cell_1rw
* cell instance $8909 r0 *1 119.85,46.41
X$8909 406 35 407 644 645 cell_1rw
* cell instance $8910 r0 *1 120.555,46.41
X$8910 408 35 409 644 645 cell_1rw
* cell instance $8911 r0 *1 121.26,46.41
X$8911 410 35 411 644 645 cell_1rw
* cell instance $8912 r0 *1 121.965,46.41
X$8912 412 35 413 644 645 cell_1rw
* cell instance $8913 r0 *1 122.67,46.41
X$8913 414 35 415 644 645 cell_1rw
* cell instance $8914 r0 *1 123.375,46.41
X$8914 416 35 417 644 645 cell_1rw
* cell instance $8915 r0 *1 124.08,46.41
X$8915 418 35 419 644 645 cell_1rw
* cell instance $8916 r0 *1 124.785,46.41
X$8916 420 35 421 644 645 cell_1rw
* cell instance $8917 r0 *1 125.49,46.41
X$8917 422 35 423 644 645 cell_1rw
* cell instance $8918 r0 *1 126.195,46.41
X$8918 424 35 425 644 645 cell_1rw
* cell instance $8919 r0 *1 126.9,46.41
X$8919 426 35 427 644 645 cell_1rw
* cell instance $8920 r0 *1 127.605,46.41
X$8920 428 35 429 644 645 cell_1rw
* cell instance $8921 r0 *1 128.31,46.41
X$8921 430 35 431 644 645 cell_1rw
* cell instance $8922 r0 *1 129.015,46.41
X$8922 432 35 433 644 645 cell_1rw
* cell instance $8923 r0 *1 129.72,46.41
X$8923 434 35 435 644 645 cell_1rw
* cell instance $8924 r0 *1 130.425,46.41
X$8924 436 35 437 644 645 cell_1rw
* cell instance $8925 r0 *1 131.13,46.41
X$8925 438 35 439 644 645 cell_1rw
* cell instance $8926 r0 *1 131.835,46.41
X$8926 440 35 441 644 645 cell_1rw
* cell instance $8927 r0 *1 132.54,46.41
X$8927 442 35 443 644 645 cell_1rw
* cell instance $8928 r0 *1 133.245,46.41
X$8928 444 35 445 644 645 cell_1rw
* cell instance $8929 r0 *1 133.95,46.41
X$8929 446 35 447 644 645 cell_1rw
* cell instance $8930 r0 *1 134.655,46.41
X$8930 448 35 449 644 645 cell_1rw
* cell instance $8931 r0 *1 135.36,46.41
X$8931 450 35 451 644 645 cell_1rw
* cell instance $8932 r0 *1 136.065,46.41
X$8932 452 35 453 644 645 cell_1rw
* cell instance $8933 r0 *1 136.77,46.41
X$8933 454 35 455 644 645 cell_1rw
* cell instance $8934 r0 *1 137.475,46.41
X$8934 456 35 457 644 645 cell_1rw
* cell instance $8935 r0 *1 138.18,46.41
X$8935 458 35 459 644 645 cell_1rw
* cell instance $8936 r0 *1 138.885,46.41
X$8936 460 35 461 644 645 cell_1rw
* cell instance $8937 r0 *1 139.59,46.41
X$8937 462 35 463 644 645 cell_1rw
* cell instance $8938 r0 *1 140.295,46.41
X$8938 464 35 465 644 645 cell_1rw
* cell instance $8939 r0 *1 141,46.41
X$8939 466 35 467 644 645 cell_1rw
* cell instance $8940 r0 *1 141.705,46.41
X$8940 468 35 469 644 645 cell_1rw
* cell instance $8941 r0 *1 142.41,46.41
X$8941 470 35 471 644 645 cell_1rw
* cell instance $8942 r0 *1 143.115,46.41
X$8942 472 35 473 644 645 cell_1rw
* cell instance $8943 r0 *1 143.82,46.41
X$8943 474 35 475 644 645 cell_1rw
* cell instance $8944 r0 *1 144.525,46.41
X$8944 476 35 477 644 645 cell_1rw
* cell instance $8945 r0 *1 145.23,46.41
X$8945 478 35 479 644 645 cell_1rw
* cell instance $8946 r0 *1 145.935,46.41
X$8946 480 35 481 644 645 cell_1rw
* cell instance $8947 r0 *1 146.64,46.41
X$8947 482 35 483 644 645 cell_1rw
* cell instance $8948 r0 *1 147.345,46.41
X$8948 484 35 485 644 645 cell_1rw
* cell instance $8949 r0 *1 148.05,46.41
X$8949 486 35 487 644 645 cell_1rw
* cell instance $8950 r0 *1 148.755,46.41
X$8950 488 35 489 644 645 cell_1rw
* cell instance $8951 r0 *1 149.46,46.41
X$8951 490 35 491 644 645 cell_1rw
* cell instance $8952 r0 *1 150.165,46.41
X$8952 492 35 493 644 645 cell_1rw
* cell instance $8953 r0 *1 150.87,46.41
X$8953 494 35 495 644 645 cell_1rw
* cell instance $8954 r0 *1 151.575,46.41
X$8954 496 35 497 644 645 cell_1rw
* cell instance $8955 r0 *1 152.28,46.41
X$8955 498 35 499 644 645 cell_1rw
* cell instance $8956 r0 *1 152.985,46.41
X$8956 500 35 501 644 645 cell_1rw
* cell instance $8957 r0 *1 153.69,46.41
X$8957 502 35 503 644 645 cell_1rw
* cell instance $8958 r0 *1 154.395,46.41
X$8958 504 35 505 644 645 cell_1rw
* cell instance $8959 r0 *1 155.1,46.41
X$8959 506 35 507 644 645 cell_1rw
* cell instance $8960 r0 *1 155.805,46.41
X$8960 508 35 509 644 645 cell_1rw
* cell instance $8961 r0 *1 156.51,46.41
X$8961 510 35 511 644 645 cell_1rw
* cell instance $8962 r0 *1 157.215,46.41
X$8962 512 35 513 644 645 cell_1rw
* cell instance $8963 r0 *1 157.92,46.41
X$8963 514 35 515 644 645 cell_1rw
* cell instance $8964 r0 *1 158.625,46.41
X$8964 516 35 517 644 645 cell_1rw
* cell instance $8965 r0 *1 159.33,46.41
X$8965 518 35 519 644 645 cell_1rw
* cell instance $8966 r0 *1 160.035,46.41
X$8966 520 35 521 644 645 cell_1rw
* cell instance $8967 r0 *1 160.74,46.41
X$8967 522 35 523 644 645 cell_1rw
* cell instance $8968 r0 *1 161.445,46.41
X$8968 524 35 525 644 645 cell_1rw
* cell instance $8969 r0 *1 162.15,46.41
X$8969 526 35 527 644 645 cell_1rw
* cell instance $8970 r0 *1 162.855,46.41
X$8970 528 35 529 644 645 cell_1rw
* cell instance $8971 r0 *1 163.56,46.41
X$8971 530 35 531 644 645 cell_1rw
* cell instance $8972 r0 *1 164.265,46.41
X$8972 532 35 533 644 645 cell_1rw
* cell instance $8973 r0 *1 164.97,46.41
X$8973 534 35 535 644 645 cell_1rw
* cell instance $8974 r0 *1 165.675,46.41
X$8974 536 35 537 644 645 cell_1rw
* cell instance $8975 r0 *1 166.38,46.41
X$8975 538 35 539 644 645 cell_1rw
* cell instance $8976 r0 *1 167.085,46.41
X$8976 540 35 541 644 645 cell_1rw
* cell instance $8977 r0 *1 167.79,46.41
X$8977 542 35 543 644 645 cell_1rw
* cell instance $8978 r0 *1 168.495,46.41
X$8978 544 35 545 644 645 cell_1rw
* cell instance $8979 r0 *1 169.2,46.41
X$8979 546 35 547 644 645 cell_1rw
* cell instance $8980 r0 *1 169.905,46.41
X$8980 548 35 549 644 645 cell_1rw
* cell instance $8981 r0 *1 170.61,46.41
X$8981 550 35 551 644 645 cell_1rw
* cell instance $8982 r0 *1 171.315,46.41
X$8982 552 35 553 644 645 cell_1rw
* cell instance $8983 r0 *1 172.02,46.41
X$8983 554 35 555 644 645 cell_1rw
* cell instance $8984 r0 *1 172.725,46.41
X$8984 556 35 557 644 645 cell_1rw
* cell instance $8985 r0 *1 173.43,46.41
X$8985 558 35 559 644 645 cell_1rw
* cell instance $8986 r0 *1 174.135,46.41
X$8986 560 35 561 644 645 cell_1rw
* cell instance $8987 r0 *1 174.84,46.41
X$8987 562 35 563 644 645 cell_1rw
* cell instance $8988 r0 *1 175.545,46.41
X$8988 564 35 565 644 645 cell_1rw
* cell instance $8989 r0 *1 176.25,46.41
X$8989 566 35 567 644 645 cell_1rw
* cell instance $8990 r0 *1 176.955,46.41
X$8990 568 35 569 644 645 cell_1rw
* cell instance $8991 r0 *1 177.66,46.41
X$8991 570 35 571 644 645 cell_1rw
* cell instance $8992 r0 *1 178.365,46.41
X$8992 572 35 573 644 645 cell_1rw
* cell instance $8993 r0 *1 179.07,46.41
X$8993 574 35 575 644 645 cell_1rw
* cell instance $8994 r0 *1 179.775,46.41
X$8994 576 35 577 644 645 cell_1rw
* cell instance $8995 r0 *1 180.48,46.41
X$8995 578 35 579 644 645 cell_1rw
* cell instance $8996 m0 *1 0.705,49.14
X$8996 67 36 68 644 645 cell_1rw
* cell instance $8997 m0 *1 0,49.14
X$8997 65 36 66 644 645 cell_1rw
* cell instance $8998 m0 *1 1.41,49.14
X$8998 69 36 70 644 645 cell_1rw
* cell instance $8999 m0 *1 2.115,49.14
X$8999 71 36 72 644 645 cell_1rw
* cell instance $9000 m0 *1 2.82,49.14
X$9000 73 36 74 644 645 cell_1rw
* cell instance $9001 m0 *1 3.525,49.14
X$9001 75 36 76 644 645 cell_1rw
* cell instance $9002 m0 *1 4.23,49.14
X$9002 77 36 78 644 645 cell_1rw
* cell instance $9003 m0 *1 4.935,49.14
X$9003 79 36 80 644 645 cell_1rw
* cell instance $9004 m0 *1 5.64,49.14
X$9004 81 36 82 644 645 cell_1rw
* cell instance $9005 m0 *1 6.345,49.14
X$9005 83 36 84 644 645 cell_1rw
* cell instance $9006 m0 *1 7.05,49.14
X$9006 85 36 86 644 645 cell_1rw
* cell instance $9007 m0 *1 7.755,49.14
X$9007 87 36 88 644 645 cell_1rw
* cell instance $9008 m0 *1 8.46,49.14
X$9008 89 36 90 644 645 cell_1rw
* cell instance $9009 m0 *1 9.165,49.14
X$9009 91 36 92 644 645 cell_1rw
* cell instance $9010 m0 *1 9.87,49.14
X$9010 93 36 94 644 645 cell_1rw
* cell instance $9011 m0 *1 10.575,49.14
X$9011 95 36 96 644 645 cell_1rw
* cell instance $9012 m0 *1 11.28,49.14
X$9012 97 36 98 644 645 cell_1rw
* cell instance $9013 m0 *1 11.985,49.14
X$9013 99 36 100 644 645 cell_1rw
* cell instance $9014 m0 *1 12.69,49.14
X$9014 101 36 102 644 645 cell_1rw
* cell instance $9015 m0 *1 13.395,49.14
X$9015 103 36 104 644 645 cell_1rw
* cell instance $9016 m0 *1 14.1,49.14
X$9016 105 36 106 644 645 cell_1rw
* cell instance $9017 m0 *1 14.805,49.14
X$9017 107 36 108 644 645 cell_1rw
* cell instance $9018 m0 *1 15.51,49.14
X$9018 109 36 110 644 645 cell_1rw
* cell instance $9019 m0 *1 16.215,49.14
X$9019 111 36 112 644 645 cell_1rw
* cell instance $9020 m0 *1 16.92,49.14
X$9020 113 36 114 644 645 cell_1rw
* cell instance $9021 m0 *1 17.625,49.14
X$9021 115 36 116 644 645 cell_1rw
* cell instance $9022 m0 *1 18.33,49.14
X$9022 117 36 118 644 645 cell_1rw
* cell instance $9023 m0 *1 19.035,49.14
X$9023 119 36 120 644 645 cell_1rw
* cell instance $9024 m0 *1 19.74,49.14
X$9024 121 36 122 644 645 cell_1rw
* cell instance $9025 m0 *1 20.445,49.14
X$9025 123 36 124 644 645 cell_1rw
* cell instance $9026 m0 *1 21.15,49.14
X$9026 125 36 126 644 645 cell_1rw
* cell instance $9027 m0 *1 21.855,49.14
X$9027 127 36 128 644 645 cell_1rw
* cell instance $9028 m0 *1 22.56,49.14
X$9028 129 36 130 644 645 cell_1rw
* cell instance $9029 m0 *1 23.265,49.14
X$9029 131 36 132 644 645 cell_1rw
* cell instance $9030 m0 *1 23.97,49.14
X$9030 133 36 134 644 645 cell_1rw
* cell instance $9031 m0 *1 24.675,49.14
X$9031 135 36 136 644 645 cell_1rw
* cell instance $9032 m0 *1 25.38,49.14
X$9032 137 36 138 644 645 cell_1rw
* cell instance $9033 m0 *1 26.085,49.14
X$9033 139 36 140 644 645 cell_1rw
* cell instance $9034 m0 *1 26.79,49.14
X$9034 141 36 142 644 645 cell_1rw
* cell instance $9035 m0 *1 27.495,49.14
X$9035 143 36 144 644 645 cell_1rw
* cell instance $9036 m0 *1 28.2,49.14
X$9036 145 36 146 644 645 cell_1rw
* cell instance $9037 m0 *1 28.905,49.14
X$9037 147 36 148 644 645 cell_1rw
* cell instance $9038 m0 *1 29.61,49.14
X$9038 149 36 150 644 645 cell_1rw
* cell instance $9039 m0 *1 30.315,49.14
X$9039 151 36 152 644 645 cell_1rw
* cell instance $9040 m0 *1 31.02,49.14
X$9040 153 36 154 644 645 cell_1rw
* cell instance $9041 m0 *1 31.725,49.14
X$9041 155 36 156 644 645 cell_1rw
* cell instance $9042 m0 *1 32.43,49.14
X$9042 157 36 158 644 645 cell_1rw
* cell instance $9043 m0 *1 33.135,49.14
X$9043 159 36 160 644 645 cell_1rw
* cell instance $9044 m0 *1 33.84,49.14
X$9044 161 36 162 644 645 cell_1rw
* cell instance $9045 m0 *1 34.545,49.14
X$9045 163 36 164 644 645 cell_1rw
* cell instance $9046 m0 *1 35.25,49.14
X$9046 165 36 166 644 645 cell_1rw
* cell instance $9047 m0 *1 35.955,49.14
X$9047 167 36 168 644 645 cell_1rw
* cell instance $9048 m0 *1 36.66,49.14
X$9048 169 36 170 644 645 cell_1rw
* cell instance $9049 m0 *1 37.365,49.14
X$9049 171 36 172 644 645 cell_1rw
* cell instance $9050 m0 *1 38.07,49.14
X$9050 173 36 174 644 645 cell_1rw
* cell instance $9051 m0 *1 38.775,49.14
X$9051 175 36 176 644 645 cell_1rw
* cell instance $9052 m0 *1 39.48,49.14
X$9052 177 36 178 644 645 cell_1rw
* cell instance $9053 m0 *1 40.185,49.14
X$9053 179 36 180 644 645 cell_1rw
* cell instance $9054 m0 *1 40.89,49.14
X$9054 181 36 182 644 645 cell_1rw
* cell instance $9055 m0 *1 41.595,49.14
X$9055 183 36 184 644 645 cell_1rw
* cell instance $9056 m0 *1 42.3,49.14
X$9056 185 36 186 644 645 cell_1rw
* cell instance $9057 m0 *1 43.005,49.14
X$9057 187 36 188 644 645 cell_1rw
* cell instance $9058 m0 *1 43.71,49.14
X$9058 189 36 190 644 645 cell_1rw
* cell instance $9059 m0 *1 44.415,49.14
X$9059 191 36 192 644 645 cell_1rw
* cell instance $9060 m0 *1 45.12,49.14
X$9060 193 36 194 644 645 cell_1rw
* cell instance $9061 m0 *1 45.825,49.14
X$9061 195 36 196 644 645 cell_1rw
* cell instance $9062 m0 *1 46.53,49.14
X$9062 197 36 198 644 645 cell_1rw
* cell instance $9063 m0 *1 47.235,49.14
X$9063 199 36 200 644 645 cell_1rw
* cell instance $9064 m0 *1 47.94,49.14
X$9064 201 36 202 644 645 cell_1rw
* cell instance $9065 m0 *1 48.645,49.14
X$9065 203 36 204 644 645 cell_1rw
* cell instance $9066 m0 *1 49.35,49.14
X$9066 205 36 206 644 645 cell_1rw
* cell instance $9067 m0 *1 50.055,49.14
X$9067 207 36 208 644 645 cell_1rw
* cell instance $9068 m0 *1 50.76,49.14
X$9068 209 36 210 644 645 cell_1rw
* cell instance $9069 m0 *1 51.465,49.14
X$9069 211 36 212 644 645 cell_1rw
* cell instance $9070 m0 *1 52.17,49.14
X$9070 213 36 214 644 645 cell_1rw
* cell instance $9071 m0 *1 52.875,49.14
X$9071 215 36 216 644 645 cell_1rw
* cell instance $9072 m0 *1 53.58,49.14
X$9072 217 36 218 644 645 cell_1rw
* cell instance $9073 m0 *1 54.285,49.14
X$9073 219 36 220 644 645 cell_1rw
* cell instance $9074 m0 *1 54.99,49.14
X$9074 221 36 222 644 645 cell_1rw
* cell instance $9075 m0 *1 55.695,49.14
X$9075 223 36 224 644 645 cell_1rw
* cell instance $9076 m0 *1 56.4,49.14
X$9076 225 36 226 644 645 cell_1rw
* cell instance $9077 m0 *1 57.105,49.14
X$9077 227 36 228 644 645 cell_1rw
* cell instance $9078 m0 *1 57.81,49.14
X$9078 229 36 230 644 645 cell_1rw
* cell instance $9079 m0 *1 58.515,49.14
X$9079 231 36 232 644 645 cell_1rw
* cell instance $9080 m0 *1 59.22,49.14
X$9080 233 36 234 644 645 cell_1rw
* cell instance $9081 m0 *1 59.925,49.14
X$9081 235 36 236 644 645 cell_1rw
* cell instance $9082 m0 *1 60.63,49.14
X$9082 237 36 238 644 645 cell_1rw
* cell instance $9083 m0 *1 61.335,49.14
X$9083 239 36 240 644 645 cell_1rw
* cell instance $9084 m0 *1 62.04,49.14
X$9084 241 36 242 644 645 cell_1rw
* cell instance $9085 m0 *1 62.745,49.14
X$9085 243 36 244 644 645 cell_1rw
* cell instance $9086 m0 *1 63.45,49.14
X$9086 245 36 246 644 645 cell_1rw
* cell instance $9087 m0 *1 64.155,49.14
X$9087 247 36 248 644 645 cell_1rw
* cell instance $9088 m0 *1 64.86,49.14
X$9088 249 36 250 644 645 cell_1rw
* cell instance $9089 m0 *1 65.565,49.14
X$9089 251 36 252 644 645 cell_1rw
* cell instance $9090 m0 *1 66.27,49.14
X$9090 253 36 254 644 645 cell_1rw
* cell instance $9091 m0 *1 66.975,49.14
X$9091 255 36 256 644 645 cell_1rw
* cell instance $9092 m0 *1 67.68,49.14
X$9092 257 36 258 644 645 cell_1rw
* cell instance $9093 m0 *1 68.385,49.14
X$9093 259 36 260 644 645 cell_1rw
* cell instance $9094 m0 *1 69.09,49.14
X$9094 261 36 262 644 645 cell_1rw
* cell instance $9095 m0 *1 69.795,49.14
X$9095 263 36 264 644 645 cell_1rw
* cell instance $9096 m0 *1 70.5,49.14
X$9096 265 36 266 644 645 cell_1rw
* cell instance $9097 m0 *1 71.205,49.14
X$9097 267 36 268 644 645 cell_1rw
* cell instance $9098 m0 *1 71.91,49.14
X$9098 269 36 270 644 645 cell_1rw
* cell instance $9099 m0 *1 72.615,49.14
X$9099 271 36 272 644 645 cell_1rw
* cell instance $9100 m0 *1 73.32,49.14
X$9100 273 36 274 644 645 cell_1rw
* cell instance $9101 m0 *1 74.025,49.14
X$9101 275 36 276 644 645 cell_1rw
* cell instance $9102 m0 *1 74.73,49.14
X$9102 277 36 278 644 645 cell_1rw
* cell instance $9103 m0 *1 75.435,49.14
X$9103 279 36 280 644 645 cell_1rw
* cell instance $9104 m0 *1 76.14,49.14
X$9104 281 36 282 644 645 cell_1rw
* cell instance $9105 m0 *1 76.845,49.14
X$9105 283 36 284 644 645 cell_1rw
* cell instance $9106 m0 *1 77.55,49.14
X$9106 285 36 286 644 645 cell_1rw
* cell instance $9107 m0 *1 78.255,49.14
X$9107 287 36 288 644 645 cell_1rw
* cell instance $9108 m0 *1 78.96,49.14
X$9108 289 36 290 644 645 cell_1rw
* cell instance $9109 m0 *1 79.665,49.14
X$9109 291 36 292 644 645 cell_1rw
* cell instance $9110 m0 *1 80.37,49.14
X$9110 293 36 294 644 645 cell_1rw
* cell instance $9111 m0 *1 81.075,49.14
X$9111 295 36 296 644 645 cell_1rw
* cell instance $9112 m0 *1 81.78,49.14
X$9112 297 36 298 644 645 cell_1rw
* cell instance $9113 m0 *1 82.485,49.14
X$9113 299 36 300 644 645 cell_1rw
* cell instance $9114 m0 *1 83.19,49.14
X$9114 301 36 302 644 645 cell_1rw
* cell instance $9115 m0 *1 83.895,49.14
X$9115 303 36 304 644 645 cell_1rw
* cell instance $9116 m0 *1 84.6,49.14
X$9116 305 36 306 644 645 cell_1rw
* cell instance $9117 m0 *1 85.305,49.14
X$9117 307 36 308 644 645 cell_1rw
* cell instance $9118 m0 *1 86.01,49.14
X$9118 309 36 310 644 645 cell_1rw
* cell instance $9119 m0 *1 86.715,49.14
X$9119 311 36 312 644 645 cell_1rw
* cell instance $9120 m0 *1 87.42,49.14
X$9120 313 36 314 644 645 cell_1rw
* cell instance $9121 m0 *1 88.125,49.14
X$9121 315 36 316 644 645 cell_1rw
* cell instance $9122 m0 *1 88.83,49.14
X$9122 317 36 318 644 645 cell_1rw
* cell instance $9123 m0 *1 89.535,49.14
X$9123 319 36 320 644 645 cell_1rw
* cell instance $9124 m0 *1 90.24,49.14
X$9124 321 36 323 644 645 cell_1rw
* cell instance $9125 m0 *1 90.945,49.14
X$9125 324 36 325 644 645 cell_1rw
* cell instance $9126 m0 *1 91.65,49.14
X$9126 326 36 327 644 645 cell_1rw
* cell instance $9127 m0 *1 92.355,49.14
X$9127 328 36 329 644 645 cell_1rw
* cell instance $9128 m0 *1 93.06,49.14
X$9128 330 36 331 644 645 cell_1rw
* cell instance $9129 m0 *1 93.765,49.14
X$9129 332 36 333 644 645 cell_1rw
* cell instance $9130 m0 *1 94.47,49.14
X$9130 334 36 335 644 645 cell_1rw
* cell instance $9131 m0 *1 95.175,49.14
X$9131 336 36 337 644 645 cell_1rw
* cell instance $9132 m0 *1 95.88,49.14
X$9132 338 36 339 644 645 cell_1rw
* cell instance $9133 m0 *1 96.585,49.14
X$9133 340 36 341 644 645 cell_1rw
* cell instance $9134 m0 *1 97.29,49.14
X$9134 342 36 343 644 645 cell_1rw
* cell instance $9135 m0 *1 97.995,49.14
X$9135 344 36 345 644 645 cell_1rw
* cell instance $9136 m0 *1 98.7,49.14
X$9136 346 36 347 644 645 cell_1rw
* cell instance $9137 m0 *1 99.405,49.14
X$9137 348 36 349 644 645 cell_1rw
* cell instance $9138 m0 *1 100.11,49.14
X$9138 350 36 351 644 645 cell_1rw
* cell instance $9139 m0 *1 100.815,49.14
X$9139 352 36 353 644 645 cell_1rw
* cell instance $9140 m0 *1 101.52,49.14
X$9140 354 36 355 644 645 cell_1rw
* cell instance $9141 m0 *1 102.225,49.14
X$9141 356 36 357 644 645 cell_1rw
* cell instance $9142 m0 *1 102.93,49.14
X$9142 358 36 359 644 645 cell_1rw
* cell instance $9143 m0 *1 103.635,49.14
X$9143 360 36 361 644 645 cell_1rw
* cell instance $9144 m0 *1 104.34,49.14
X$9144 362 36 363 644 645 cell_1rw
* cell instance $9145 m0 *1 105.045,49.14
X$9145 364 36 365 644 645 cell_1rw
* cell instance $9146 m0 *1 105.75,49.14
X$9146 366 36 367 644 645 cell_1rw
* cell instance $9147 m0 *1 106.455,49.14
X$9147 368 36 369 644 645 cell_1rw
* cell instance $9148 m0 *1 107.16,49.14
X$9148 370 36 371 644 645 cell_1rw
* cell instance $9149 m0 *1 107.865,49.14
X$9149 372 36 373 644 645 cell_1rw
* cell instance $9150 m0 *1 108.57,49.14
X$9150 374 36 375 644 645 cell_1rw
* cell instance $9151 m0 *1 109.275,49.14
X$9151 376 36 377 644 645 cell_1rw
* cell instance $9152 m0 *1 109.98,49.14
X$9152 378 36 379 644 645 cell_1rw
* cell instance $9153 m0 *1 110.685,49.14
X$9153 380 36 381 644 645 cell_1rw
* cell instance $9154 m0 *1 111.39,49.14
X$9154 382 36 383 644 645 cell_1rw
* cell instance $9155 m0 *1 112.095,49.14
X$9155 384 36 385 644 645 cell_1rw
* cell instance $9156 m0 *1 112.8,49.14
X$9156 386 36 387 644 645 cell_1rw
* cell instance $9157 m0 *1 113.505,49.14
X$9157 388 36 389 644 645 cell_1rw
* cell instance $9158 m0 *1 114.21,49.14
X$9158 390 36 391 644 645 cell_1rw
* cell instance $9159 m0 *1 114.915,49.14
X$9159 392 36 393 644 645 cell_1rw
* cell instance $9160 m0 *1 115.62,49.14
X$9160 394 36 395 644 645 cell_1rw
* cell instance $9161 m0 *1 116.325,49.14
X$9161 396 36 397 644 645 cell_1rw
* cell instance $9162 m0 *1 117.03,49.14
X$9162 398 36 399 644 645 cell_1rw
* cell instance $9163 m0 *1 117.735,49.14
X$9163 400 36 401 644 645 cell_1rw
* cell instance $9164 m0 *1 118.44,49.14
X$9164 402 36 403 644 645 cell_1rw
* cell instance $9165 m0 *1 119.145,49.14
X$9165 404 36 405 644 645 cell_1rw
* cell instance $9166 m0 *1 119.85,49.14
X$9166 406 36 407 644 645 cell_1rw
* cell instance $9167 m0 *1 120.555,49.14
X$9167 408 36 409 644 645 cell_1rw
* cell instance $9168 m0 *1 121.26,49.14
X$9168 410 36 411 644 645 cell_1rw
* cell instance $9169 m0 *1 121.965,49.14
X$9169 412 36 413 644 645 cell_1rw
* cell instance $9170 m0 *1 122.67,49.14
X$9170 414 36 415 644 645 cell_1rw
* cell instance $9171 m0 *1 123.375,49.14
X$9171 416 36 417 644 645 cell_1rw
* cell instance $9172 m0 *1 124.08,49.14
X$9172 418 36 419 644 645 cell_1rw
* cell instance $9173 m0 *1 124.785,49.14
X$9173 420 36 421 644 645 cell_1rw
* cell instance $9174 m0 *1 125.49,49.14
X$9174 422 36 423 644 645 cell_1rw
* cell instance $9175 m0 *1 126.195,49.14
X$9175 424 36 425 644 645 cell_1rw
* cell instance $9176 m0 *1 126.9,49.14
X$9176 426 36 427 644 645 cell_1rw
* cell instance $9177 m0 *1 127.605,49.14
X$9177 428 36 429 644 645 cell_1rw
* cell instance $9178 m0 *1 128.31,49.14
X$9178 430 36 431 644 645 cell_1rw
* cell instance $9179 m0 *1 129.015,49.14
X$9179 432 36 433 644 645 cell_1rw
* cell instance $9180 m0 *1 129.72,49.14
X$9180 434 36 435 644 645 cell_1rw
* cell instance $9181 m0 *1 130.425,49.14
X$9181 436 36 437 644 645 cell_1rw
* cell instance $9182 m0 *1 131.13,49.14
X$9182 438 36 439 644 645 cell_1rw
* cell instance $9183 m0 *1 131.835,49.14
X$9183 440 36 441 644 645 cell_1rw
* cell instance $9184 m0 *1 132.54,49.14
X$9184 442 36 443 644 645 cell_1rw
* cell instance $9185 m0 *1 133.245,49.14
X$9185 444 36 445 644 645 cell_1rw
* cell instance $9186 m0 *1 133.95,49.14
X$9186 446 36 447 644 645 cell_1rw
* cell instance $9187 m0 *1 134.655,49.14
X$9187 448 36 449 644 645 cell_1rw
* cell instance $9188 m0 *1 135.36,49.14
X$9188 450 36 451 644 645 cell_1rw
* cell instance $9189 m0 *1 136.065,49.14
X$9189 452 36 453 644 645 cell_1rw
* cell instance $9190 m0 *1 136.77,49.14
X$9190 454 36 455 644 645 cell_1rw
* cell instance $9191 m0 *1 137.475,49.14
X$9191 456 36 457 644 645 cell_1rw
* cell instance $9192 m0 *1 138.18,49.14
X$9192 458 36 459 644 645 cell_1rw
* cell instance $9193 m0 *1 138.885,49.14
X$9193 460 36 461 644 645 cell_1rw
* cell instance $9194 m0 *1 139.59,49.14
X$9194 462 36 463 644 645 cell_1rw
* cell instance $9195 m0 *1 140.295,49.14
X$9195 464 36 465 644 645 cell_1rw
* cell instance $9196 m0 *1 141,49.14
X$9196 466 36 467 644 645 cell_1rw
* cell instance $9197 m0 *1 141.705,49.14
X$9197 468 36 469 644 645 cell_1rw
* cell instance $9198 m0 *1 142.41,49.14
X$9198 470 36 471 644 645 cell_1rw
* cell instance $9199 m0 *1 143.115,49.14
X$9199 472 36 473 644 645 cell_1rw
* cell instance $9200 m0 *1 143.82,49.14
X$9200 474 36 475 644 645 cell_1rw
* cell instance $9201 m0 *1 144.525,49.14
X$9201 476 36 477 644 645 cell_1rw
* cell instance $9202 m0 *1 145.23,49.14
X$9202 478 36 479 644 645 cell_1rw
* cell instance $9203 m0 *1 145.935,49.14
X$9203 480 36 481 644 645 cell_1rw
* cell instance $9204 m0 *1 146.64,49.14
X$9204 482 36 483 644 645 cell_1rw
* cell instance $9205 m0 *1 147.345,49.14
X$9205 484 36 485 644 645 cell_1rw
* cell instance $9206 m0 *1 148.05,49.14
X$9206 486 36 487 644 645 cell_1rw
* cell instance $9207 m0 *1 148.755,49.14
X$9207 488 36 489 644 645 cell_1rw
* cell instance $9208 m0 *1 149.46,49.14
X$9208 490 36 491 644 645 cell_1rw
* cell instance $9209 m0 *1 150.165,49.14
X$9209 492 36 493 644 645 cell_1rw
* cell instance $9210 m0 *1 150.87,49.14
X$9210 494 36 495 644 645 cell_1rw
* cell instance $9211 m0 *1 151.575,49.14
X$9211 496 36 497 644 645 cell_1rw
* cell instance $9212 m0 *1 152.28,49.14
X$9212 498 36 499 644 645 cell_1rw
* cell instance $9213 m0 *1 152.985,49.14
X$9213 500 36 501 644 645 cell_1rw
* cell instance $9214 m0 *1 153.69,49.14
X$9214 502 36 503 644 645 cell_1rw
* cell instance $9215 m0 *1 154.395,49.14
X$9215 504 36 505 644 645 cell_1rw
* cell instance $9216 m0 *1 155.1,49.14
X$9216 506 36 507 644 645 cell_1rw
* cell instance $9217 m0 *1 155.805,49.14
X$9217 508 36 509 644 645 cell_1rw
* cell instance $9218 m0 *1 156.51,49.14
X$9218 510 36 511 644 645 cell_1rw
* cell instance $9219 m0 *1 157.215,49.14
X$9219 512 36 513 644 645 cell_1rw
* cell instance $9220 m0 *1 157.92,49.14
X$9220 514 36 515 644 645 cell_1rw
* cell instance $9221 m0 *1 158.625,49.14
X$9221 516 36 517 644 645 cell_1rw
* cell instance $9222 m0 *1 159.33,49.14
X$9222 518 36 519 644 645 cell_1rw
* cell instance $9223 m0 *1 160.035,49.14
X$9223 520 36 521 644 645 cell_1rw
* cell instance $9224 m0 *1 160.74,49.14
X$9224 522 36 523 644 645 cell_1rw
* cell instance $9225 m0 *1 161.445,49.14
X$9225 524 36 525 644 645 cell_1rw
* cell instance $9226 m0 *1 162.15,49.14
X$9226 526 36 527 644 645 cell_1rw
* cell instance $9227 m0 *1 162.855,49.14
X$9227 528 36 529 644 645 cell_1rw
* cell instance $9228 m0 *1 163.56,49.14
X$9228 530 36 531 644 645 cell_1rw
* cell instance $9229 m0 *1 164.265,49.14
X$9229 532 36 533 644 645 cell_1rw
* cell instance $9230 m0 *1 164.97,49.14
X$9230 534 36 535 644 645 cell_1rw
* cell instance $9231 m0 *1 165.675,49.14
X$9231 536 36 537 644 645 cell_1rw
* cell instance $9232 m0 *1 166.38,49.14
X$9232 538 36 539 644 645 cell_1rw
* cell instance $9233 m0 *1 167.085,49.14
X$9233 540 36 541 644 645 cell_1rw
* cell instance $9234 m0 *1 167.79,49.14
X$9234 542 36 543 644 645 cell_1rw
* cell instance $9235 m0 *1 168.495,49.14
X$9235 544 36 545 644 645 cell_1rw
* cell instance $9236 m0 *1 169.2,49.14
X$9236 546 36 547 644 645 cell_1rw
* cell instance $9237 m0 *1 169.905,49.14
X$9237 548 36 549 644 645 cell_1rw
* cell instance $9238 m0 *1 170.61,49.14
X$9238 550 36 551 644 645 cell_1rw
* cell instance $9239 m0 *1 171.315,49.14
X$9239 552 36 553 644 645 cell_1rw
* cell instance $9240 m0 *1 172.02,49.14
X$9240 554 36 555 644 645 cell_1rw
* cell instance $9241 m0 *1 172.725,49.14
X$9241 556 36 557 644 645 cell_1rw
* cell instance $9242 m0 *1 173.43,49.14
X$9242 558 36 559 644 645 cell_1rw
* cell instance $9243 m0 *1 174.135,49.14
X$9243 560 36 561 644 645 cell_1rw
* cell instance $9244 m0 *1 174.84,49.14
X$9244 562 36 563 644 645 cell_1rw
* cell instance $9245 m0 *1 175.545,49.14
X$9245 564 36 565 644 645 cell_1rw
* cell instance $9246 m0 *1 176.25,49.14
X$9246 566 36 567 644 645 cell_1rw
* cell instance $9247 m0 *1 176.955,49.14
X$9247 568 36 569 644 645 cell_1rw
* cell instance $9248 m0 *1 177.66,49.14
X$9248 570 36 571 644 645 cell_1rw
* cell instance $9249 m0 *1 178.365,49.14
X$9249 572 36 573 644 645 cell_1rw
* cell instance $9250 m0 *1 179.07,49.14
X$9250 574 36 575 644 645 cell_1rw
* cell instance $9251 m0 *1 179.775,49.14
X$9251 576 36 577 644 645 cell_1rw
* cell instance $9252 m0 *1 180.48,49.14
X$9252 578 36 579 644 645 cell_1rw
* cell instance $9253 r0 *1 0.705,49.14
X$9253 67 37 68 644 645 cell_1rw
* cell instance $9254 r0 *1 0,49.14
X$9254 65 37 66 644 645 cell_1rw
* cell instance $9255 r0 *1 1.41,49.14
X$9255 69 37 70 644 645 cell_1rw
* cell instance $9256 r0 *1 2.115,49.14
X$9256 71 37 72 644 645 cell_1rw
* cell instance $9257 r0 *1 2.82,49.14
X$9257 73 37 74 644 645 cell_1rw
* cell instance $9258 r0 *1 3.525,49.14
X$9258 75 37 76 644 645 cell_1rw
* cell instance $9259 r0 *1 4.23,49.14
X$9259 77 37 78 644 645 cell_1rw
* cell instance $9260 r0 *1 4.935,49.14
X$9260 79 37 80 644 645 cell_1rw
* cell instance $9261 r0 *1 5.64,49.14
X$9261 81 37 82 644 645 cell_1rw
* cell instance $9262 r0 *1 6.345,49.14
X$9262 83 37 84 644 645 cell_1rw
* cell instance $9263 r0 *1 7.05,49.14
X$9263 85 37 86 644 645 cell_1rw
* cell instance $9264 r0 *1 7.755,49.14
X$9264 87 37 88 644 645 cell_1rw
* cell instance $9265 r0 *1 8.46,49.14
X$9265 89 37 90 644 645 cell_1rw
* cell instance $9266 r0 *1 9.165,49.14
X$9266 91 37 92 644 645 cell_1rw
* cell instance $9267 r0 *1 9.87,49.14
X$9267 93 37 94 644 645 cell_1rw
* cell instance $9268 r0 *1 10.575,49.14
X$9268 95 37 96 644 645 cell_1rw
* cell instance $9269 r0 *1 11.28,49.14
X$9269 97 37 98 644 645 cell_1rw
* cell instance $9270 r0 *1 11.985,49.14
X$9270 99 37 100 644 645 cell_1rw
* cell instance $9271 r0 *1 12.69,49.14
X$9271 101 37 102 644 645 cell_1rw
* cell instance $9272 r0 *1 13.395,49.14
X$9272 103 37 104 644 645 cell_1rw
* cell instance $9273 r0 *1 14.1,49.14
X$9273 105 37 106 644 645 cell_1rw
* cell instance $9274 r0 *1 14.805,49.14
X$9274 107 37 108 644 645 cell_1rw
* cell instance $9275 r0 *1 15.51,49.14
X$9275 109 37 110 644 645 cell_1rw
* cell instance $9276 r0 *1 16.215,49.14
X$9276 111 37 112 644 645 cell_1rw
* cell instance $9277 r0 *1 16.92,49.14
X$9277 113 37 114 644 645 cell_1rw
* cell instance $9278 r0 *1 17.625,49.14
X$9278 115 37 116 644 645 cell_1rw
* cell instance $9279 r0 *1 18.33,49.14
X$9279 117 37 118 644 645 cell_1rw
* cell instance $9280 r0 *1 19.035,49.14
X$9280 119 37 120 644 645 cell_1rw
* cell instance $9281 r0 *1 19.74,49.14
X$9281 121 37 122 644 645 cell_1rw
* cell instance $9282 r0 *1 20.445,49.14
X$9282 123 37 124 644 645 cell_1rw
* cell instance $9283 r0 *1 21.15,49.14
X$9283 125 37 126 644 645 cell_1rw
* cell instance $9284 r0 *1 21.855,49.14
X$9284 127 37 128 644 645 cell_1rw
* cell instance $9285 r0 *1 22.56,49.14
X$9285 129 37 130 644 645 cell_1rw
* cell instance $9286 r0 *1 23.265,49.14
X$9286 131 37 132 644 645 cell_1rw
* cell instance $9287 r0 *1 23.97,49.14
X$9287 133 37 134 644 645 cell_1rw
* cell instance $9288 r0 *1 24.675,49.14
X$9288 135 37 136 644 645 cell_1rw
* cell instance $9289 r0 *1 25.38,49.14
X$9289 137 37 138 644 645 cell_1rw
* cell instance $9290 r0 *1 26.085,49.14
X$9290 139 37 140 644 645 cell_1rw
* cell instance $9291 r0 *1 26.79,49.14
X$9291 141 37 142 644 645 cell_1rw
* cell instance $9292 r0 *1 27.495,49.14
X$9292 143 37 144 644 645 cell_1rw
* cell instance $9293 r0 *1 28.2,49.14
X$9293 145 37 146 644 645 cell_1rw
* cell instance $9294 r0 *1 28.905,49.14
X$9294 147 37 148 644 645 cell_1rw
* cell instance $9295 r0 *1 29.61,49.14
X$9295 149 37 150 644 645 cell_1rw
* cell instance $9296 r0 *1 30.315,49.14
X$9296 151 37 152 644 645 cell_1rw
* cell instance $9297 r0 *1 31.02,49.14
X$9297 153 37 154 644 645 cell_1rw
* cell instance $9298 r0 *1 31.725,49.14
X$9298 155 37 156 644 645 cell_1rw
* cell instance $9299 r0 *1 32.43,49.14
X$9299 157 37 158 644 645 cell_1rw
* cell instance $9300 r0 *1 33.135,49.14
X$9300 159 37 160 644 645 cell_1rw
* cell instance $9301 r0 *1 33.84,49.14
X$9301 161 37 162 644 645 cell_1rw
* cell instance $9302 r0 *1 34.545,49.14
X$9302 163 37 164 644 645 cell_1rw
* cell instance $9303 r0 *1 35.25,49.14
X$9303 165 37 166 644 645 cell_1rw
* cell instance $9304 r0 *1 35.955,49.14
X$9304 167 37 168 644 645 cell_1rw
* cell instance $9305 r0 *1 36.66,49.14
X$9305 169 37 170 644 645 cell_1rw
* cell instance $9306 r0 *1 37.365,49.14
X$9306 171 37 172 644 645 cell_1rw
* cell instance $9307 r0 *1 38.07,49.14
X$9307 173 37 174 644 645 cell_1rw
* cell instance $9308 r0 *1 38.775,49.14
X$9308 175 37 176 644 645 cell_1rw
* cell instance $9309 r0 *1 39.48,49.14
X$9309 177 37 178 644 645 cell_1rw
* cell instance $9310 r0 *1 40.185,49.14
X$9310 179 37 180 644 645 cell_1rw
* cell instance $9311 r0 *1 40.89,49.14
X$9311 181 37 182 644 645 cell_1rw
* cell instance $9312 r0 *1 41.595,49.14
X$9312 183 37 184 644 645 cell_1rw
* cell instance $9313 r0 *1 42.3,49.14
X$9313 185 37 186 644 645 cell_1rw
* cell instance $9314 r0 *1 43.005,49.14
X$9314 187 37 188 644 645 cell_1rw
* cell instance $9315 r0 *1 43.71,49.14
X$9315 189 37 190 644 645 cell_1rw
* cell instance $9316 r0 *1 44.415,49.14
X$9316 191 37 192 644 645 cell_1rw
* cell instance $9317 r0 *1 45.12,49.14
X$9317 193 37 194 644 645 cell_1rw
* cell instance $9318 r0 *1 45.825,49.14
X$9318 195 37 196 644 645 cell_1rw
* cell instance $9319 r0 *1 46.53,49.14
X$9319 197 37 198 644 645 cell_1rw
* cell instance $9320 r0 *1 47.235,49.14
X$9320 199 37 200 644 645 cell_1rw
* cell instance $9321 r0 *1 47.94,49.14
X$9321 201 37 202 644 645 cell_1rw
* cell instance $9322 r0 *1 48.645,49.14
X$9322 203 37 204 644 645 cell_1rw
* cell instance $9323 r0 *1 49.35,49.14
X$9323 205 37 206 644 645 cell_1rw
* cell instance $9324 r0 *1 50.055,49.14
X$9324 207 37 208 644 645 cell_1rw
* cell instance $9325 r0 *1 50.76,49.14
X$9325 209 37 210 644 645 cell_1rw
* cell instance $9326 r0 *1 51.465,49.14
X$9326 211 37 212 644 645 cell_1rw
* cell instance $9327 r0 *1 52.17,49.14
X$9327 213 37 214 644 645 cell_1rw
* cell instance $9328 r0 *1 52.875,49.14
X$9328 215 37 216 644 645 cell_1rw
* cell instance $9329 r0 *1 53.58,49.14
X$9329 217 37 218 644 645 cell_1rw
* cell instance $9330 r0 *1 54.285,49.14
X$9330 219 37 220 644 645 cell_1rw
* cell instance $9331 r0 *1 54.99,49.14
X$9331 221 37 222 644 645 cell_1rw
* cell instance $9332 r0 *1 55.695,49.14
X$9332 223 37 224 644 645 cell_1rw
* cell instance $9333 r0 *1 56.4,49.14
X$9333 225 37 226 644 645 cell_1rw
* cell instance $9334 r0 *1 57.105,49.14
X$9334 227 37 228 644 645 cell_1rw
* cell instance $9335 r0 *1 57.81,49.14
X$9335 229 37 230 644 645 cell_1rw
* cell instance $9336 r0 *1 58.515,49.14
X$9336 231 37 232 644 645 cell_1rw
* cell instance $9337 r0 *1 59.22,49.14
X$9337 233 37 234 644 645 cell_1rw
* cell instance $9338 r0 *1 59.925,49.14
X$9338 235 37 236 644 645 cell_1rw
* cell instance $9339 r0 *1 60.63,49.14
X$9339 237 37 238 644 645 cell_1rw
* cell instance $9340 r0 *1 61.335,49.14
X$9340 239 37 240 644 645 cell_1rw
* cell instance $9341 r0 *1 62.04,49.14
X$9341 241 37 242 644 645 cell_1rw
* cell instance $9342 r0 *1 62.745,49.14
X$9342 243 37 244 644 645 cell_1rw
* cell instance $9343 r0 *1 63.45,49.14
X$9343 245 37 246 644 645 cell_1rw
* cell instance $9344 r0 *1 64.155,49.14
X$9344 247 37 248 644 645 cell_1rw
* cell instance $9345 r0 *1 64.86,49.14
X$9345 249 37 250 644 645 cell_1rw
* cell instance $9346 r0 *1 65.565,49.14
X$9346 251 37 252 644 645 cell_1rw
* cell instance $9347 r0 *1 66.27,49.14
X$9347 253 37 254 644 645 cell_1rw
* cell instance $9348 r0 *1 66.975,49.14
X$9348 255 37 256 644 645 cell_1rw
* cell instance $9349 r0 *1 67.68,49.14
X$9349 257 37 258 644 645 cell_1rw
* cell instance $9350 r0 *1 68.385,49.14
X$9350 259 37 260 644 645 cell_1rw
* cell instance $9351 r0 *1 69.09,49.14
X$9351 261 37 262 644 645 cell_1rw
* cell instance $9352 r0 *1 69.795,49.14
X$9352 263 37 264 644 645 cell_1rw
* cell instance $9353 r0 *1 70.5,49.14
X$9353 265 37 266 644 645 cell_1rw
* cell instance $9354 r0 *1 71.205,49.14
X$9354 267 37 268 644 645 cell_1rw
* cell instance $9355 r0 *1 71.91,49.14
X$9355 269 37 270 644 645 cell_1rw
* cell instance $9356 r0 *1 72.615,49.14
X$9356 271 37 272 644 645 cell_1rw
* cell instance $9357 r0 *1 73.32,49.14
X$9357 273 37 274 644 645 cell_1rw
* cell instance $9358 r0 *1 74.025,49.14
X$9358 275 37 276 644 645 cell_1rw
* cell instance $9359 r0 *1 74.73,49.14
X$9359 277 37 278 644 645 cell_1rw
* cell instance $9360 r0 *1 75.435,49.14
X$9360 279 37 280 644 645 cell_1rw
* cell instance $9361 r0 *1 76.14,49.14
X$9361 281 37 282 644 645 cell_1rw
* cell instance $9362 r0 *1 76.845,49.14
X$9362 283 37 284 644 645 cell_1rw
* cell instance $9363 r0 *1 77.55,49.14
X$9363 285 37 286 644 645 cell_1rw
* cell instance $9364 r0 *1 78.255,49.14
X$9364 287 37 288 644 645 cell_1rw
* cell instance $9365 r0 *1 78.96,49.14
X$9365 289 37 290 644 645 cell_1rw
* cell instance $9366 r0 *1 79.665,49.14
X$9366 291 37 292 644 645 cell_1rw
* cell instance $9367 r0 *1 80.37,49.14
X$9367 293 37 294 644 645 cell_1rw
* cell instance $9368 r0 *1 81.075,49.14
X$9368 295 37 296 644 645 cell_1rw
* cell instance $9369 r0 *1 81.78,49.14
X$9369 297 37 298 644 645 cell_1rw
* cell instance $9370 r0 *1 82.485,49.14
X$9370 299 37 300 644 645 cell_1rw
* cell instance $9371 r0 *1 83.19,49.14
X$9371 301 37 302 644 645 cell_1rw
* cell instance $9372 r0 *1 83.895,49.14
X$9372 303 37 304 644 645 cell_1rw
* cell instance $9373 r0 *1 84.6,49.14
X$9373 305 37 306 644 645 cell_1rw
* cell instance $9374 r0 *1 85.305,49.14
X$9374 307 37 308 644 645 cell_1rw
* cell instance $9375 r0 *1 86.01,49.14
X$9375 309 37 310 644 645 cell_1rw
* cell instance $9376 r0 *1 86.715,49.14
X$9376 311 37 312 644 645 cell_1rw
* cell instance $9377 r0 *1 87.42,49.14
X$9377 313 37 314 644 645 cell_1rw
* cell instance $9378 r0 *1 88.125,49.14
X$9378 315 37 316 644 645 cell_1rw
* cell instance $9379 r0 *1 88.83,49.14
X$9379 317 37 318 644 645 cell_1rw
* cell instance $9380 r0 *1 89.535,49.14
X$9380 319 37 320 644 645 cell_1rw
* cell instance $9381 r0 *1 90.24,49.14
X$9381 321 37 323 644 645 cell_1rw
* cell instance $9382 r0 *1 90.945,49.14
X$9382 324 37 325 644 645 cell_1rw
* cell instance $9383 r0 *1 91.65,49.14
X$9383 326 37 327 644 645 cell_1rw
* cell instance $9384 r0 *1 92.355,49.14
X$9384 328 37 329 644 645 cell_1rw
* cell instance $9385 r0 *1 93.06,49.14
X$9385 330 37 331 644 645 cell_1rw
* cell instance $9386 r0 *1 93.765,49.14
X$9386 332 37 333 644 645 cell_1rw
* cell instance $9387 r0 *1 94.47,49.14
X$9387 334 37 335 644 645 cell_1rw
* cell instance $9388 r0 *1 95.175,49.14
X$9388 336 37 337 644 645 cell_1rw
* cell instance $9389 r0 *1 95.88,49.14
X$9389 338 37 339 644 645 cell_1rw
* cell instance $9390 r0 *1 96.585,49.14
X$9390 340 37 341 644 645 cell_1rw
* cell instance $9391 r0 *1 97.29,49.14
X$9391 342 37 343 644 645 cell_1rw
* cell instance $9392 r0 *1 97.995,49.14
X$9392 344 37 345 644 645 cell_1rw
* cell instance $9393 r0 *1 98.7,49.14
X$9393 346 37 347 644 645 cell_1rw
* cell instance $9394 r0 *1 99.405,49.14
X$9394 348 37 349 644 645 cell_1rw
* cell instance $9395 r0 *1 100.11,49.14
X$9395 350 37 351 644 645 cell_1rw
* cell instance $9396 r0 *1 100.815,49.14
X$9396 352 37 353 644 645 cell_1rw
* cell instance $9397 r0 *1 101.52,49.14
X$9397 354 37 355 644 645 cell_1rw
* cell instance $9398 r0 *1 102.225,49.14
X$9398 356 37 357 644 645 cell_1rw
* cell instance $9399 r0 *1 102.93,49.14
X$9399 358 37 359 644 645 cell_1rw
* cell instance $9400 r0 *1 103.635,49.14
X$9400 360 37 361 644 645 cell_1rw
* cell instance $9401 r0 *1 104.34,49.14
X$9401 362 37 363 644 645 cell_1rw
* cell instance $9402 r0 *1 105.045,49.14
X$9402 364 37 365 644 645 cell_1rw
* cell instance $9403 r0 *1 105.75,49.14
X$9403 366 37 367 644 645 cell_1rw
* cell instance $9404 r0 *1 106.455,49.14
X$9404 368 37 369 644 645 cell_1rw
* cell instance $9405 r0 *1 107.16,49.14
X$9405 370 37 371 644 645 cell_1rw
* cell instance $9406 r0 *1 107.865,49.14
X$9406 372 37 373 644 645 cell_1rw
* cell instance $9407 r0 *1 108.57,49.14
X$9407 374 37 375 644 645 cell_1rw
* cell instance $9408 r0 *1 109.275,49.14
X$9408 376 37 377 644 645 cell_1rw
* cell instance $9409 r0 *1 109.98,49.14
X$9409 378 37 379 644 645 cell_1rw
* cell instance $9410 r0 *1 110.685,49.14
X$9410 380 37 381 644 645 cell_1rw
* cell instance $9411 r0 *1 111.39,49.14
X$9411 382 37 383 644 645 cell_1rw
* cell instance $9412 r0 *1 112.095,49.14
X$9412 384 37 385 644 645 cell_1rw
* cell instance $9413 r0 *1 112.8,49.14
X$9413 386 37 387 644 645 cell_1rw
* cell instance $9414 r0 *1 113.505,49.14
X$9414 388 37 389 644 645 cell_1rw
* cell instance $9415 r0 *1 114.21,49.14
X$9415 390 37 391 644 645 cell_1rw
* cell instance $9416 r0 *1 114.915,49.14
X$9416 392 37 393 644 645 cell_1rw
* cell instance $9417 r0 *1 115.62,49.14
X$9417 394 37 395 644 645 cell_1rw
* cell instance $9418 r0 *1 116.325,49.14
X$9418 396 37 397 644 645 cell_1rw
* cell instance $9419 r0 *1 117.03,49.14
X$9419 398 37 399 644 645 cell_1rw
* cell instance $9420 r0 *1 117.735,49.14
X$9420 400 37 401 644 645 cell_1rw
* cell instance $9421 r0 *1 118.44,49.14
X$9421 402 37 403 644 645 cell_1rw
* cell instance $9422 r0 *1 119.145,49.14
X$9422 404 37 405 644 645 cell_1rw
* cell instance $9423 r0 *1 119.85,49.14
X$9423 406 37 407 644 645 cell_1rw
* cell instance $9424 r0 *1 120.555,49.14
X$9424 408 37 409 644 645 cell_1rw
* cell instance $9425 r0 *1 121.26,49.14
X$9425 410 37 411 644 645 cell_1rw
* cell instance $9426 r0 *1 121.965,49.14
X$9426 412 37 413 644 645 cell_1rw
* cell instance $9427 r0 *1 122.67,49.14
X$9427 414 37 415 644 645 cell_1rw
* cell instance $9428 r0 *1 123.375,49.14
X$9428 416 37 417 644 645 cell_1rw
* cell instance $9429 r0 *1 124.08,49.14
X$9429 418 37 419 644 645 cell_1rw
* cell instance $9430 r0 *1 124.785,49.14
X$9430 420 37 421 644 645 cell_1rw
* cell instance $9431 r0 *1 125.49,49.14
X$9431 422 37 423 644 645 cell_1rw
* cell instance $9432 r0 *1 126.195,49.14
X$9432 424 37 425 644 645 cell_1rw
* cell instance $9433 r0 *1 126.9,49.14
X$9433 426 37 427 644 645 cell_1rw
* cell instance $9434 r0 *1 127.605,49.14
X$9434 428 37 429 644 645 cell_1rw
* cell instance $9435 r0 *1 128.31,49.14
X$9435 430 37 431 644 645 cell_1rw
* cell instance $9436 r0 *1 129.015,49.14
X$9436 432 37 433 644 645 cell_1rw
* cell instance $9437 r0 *1 129.72,49.14
X$9437 434 37 435 644 645 cell_1rw
* cell instance $9438 r0 *1 130.425,49.14
X$9438 436 37 437 644 645 cell_1rw
* cell instance $9439 r0 *1 131.13,49.14
X$9439 438 37 439 644 645 cell_1rw
* cell instance $9440 r0 *1 131.835,49.14
X$9440 440 37 441 644 645 cell_1rw
* cell instance $9441 r0 *1 132.54,49.14
X$9441 442 37 443 644 645 cell_1rw
* cell instance $9442 r0 *1 133.245,49.14
X$9442 444 37 445 644 645 cell_1rw
* cell instance $9443 r0 *1 133.95,49.14
X$9443 446 37 447 644 645 cell_1rw
* cell instance $9444 r0 *1 134.655,49.14
X$9444 448 37 449 644 645 cell_1rw
* cell instance $9445 r0 *1 135.36,49.14
X$9445 450 37 451 644 645 cell_1rw
* cell instance $9446 r0 *1 136.065,49.14
X$9446 452 37 453 644 645 cell_1rw
* cell instance $9447 r0 *1 136.77,49.14
X$9447 454 37 455 644 645 cell_1rw
* cell instance $9448 r0 *1 137.475,49.14
X$9448 456 37 457 644 645 cell_1rw
* cell instance $9449 r0 *1 138.18,49.14
X$9449 458 37 459 644 645 cell_1rw
* cell instance $9450 r0 *1 138.885,49.14
X$9450 460 37 461 644 645 cell_1rw
* cell instance $9451 r0 *1 139.59,49.14
X$9451 462 37 463 644 645 cell_1rw
* cell instance $9452 r0 *1 140.295,49.14
X$9452 464 37 465 644 645 cell_1rw
* cell instance $9453 r0 *1 141,49.14
X$9453 466 37 467 644 645 cell_1rw
* cell instance $9454 r0 *1 141.705,49.14
X$9454 468 37 469 644 645 cell_1rw
* cell instance $9455 r0 *1 142.41,49.14
X$9455 470 37 471 644 645 cell_1rw
* cell instance $9456 r0 *1 143.115,49.14
X$9456 472 37 473 644 645 cell_1rw
* cell instance $9457 r0 *1 143.82,49.14
X$9457 474 37 475 644 645 cell_1rw
* cell instance $9458 r0 *1 144.525,49.14
X$9458 476 37 477 644 645 cell_1rw
* cell instance $9459 r0 *1 145.23,49.14
X$9459 478 37 479 644 645 cell_1rw
* cell instance $9460 r0 *1 145.935,49.14
X$9460 480 37 481 644 645 cell_1rw
* cell instance $9461 r0 *1 146.64,49.14
X$9461 482 37 483 644 645 cell_1rw
* cell instance $9462 r0 *1 147.345,49.14
X$9462 484 37 485 644 645 cell_1rw
* cell instance $9463 r0 *1 148.05,49.14
X$9463 486 37 487 644 645 cell_1rw
* cell instance $9464 r0 *1 148.755,49.14
X$9464 488 37 489 644 645 cell_1rw
* cell instance $9465 r0 *1 149.46,49.14
X$9465 490 37 491 644 645 cell_1rw
* cell instance $9466 r0 *1 150.165,49.14
X$9466 492 37 493 644 645 cell_1rw
* cell instance $9467 r0 *1 150.87,49.14
X$9467 494 37 495 644 645 cell_1rw
* cell instance $9468 r0 *1 151.575,49.14
X$9468 496 37 497 644 645 cell_1rw
* cell instance $9469 r0 *1 152.28,49.14
X$9469 498 37 499 644 645 cell_1rw
* cell instance $9470 r0 *1 152.985,49.14
X$9470 500 37 501 644 645 cell_1rw
* cell instance $9471 r0 *1 153.69,49.14
X$9471 502 37 503 644 645 cell_1rw
* cell instance $9472 r0 *1 154.395,49.14
X$9472 504 37 505 644 645 cell_1rw
* cell instance $9473 r0 *1 155.1,49.14
X$9473 506 37 507 644 645 cell_1rw
* cell instance $9474 r0 *1 155.805,49.14
X$9474 508 37 509 644 645 cell_1rw
* cell instance $9475 r0 *1 156.51,49.14
X$9475 510 37 511 644 645 cell_1rw
* cell instance $9476 r0 *1 157.215,49.14
X$9476 512 37 513 644 645 cell_1rw
* cell instance $9477 r0 *1 157.92,49.14
X$9477 514 37 515 644 645 cell_1rw
* cell instance $9478 r0 *1 158.625,49.14
X$9478 516 37 517 644 645 cell_1rw
* cell instance $9479 r0 *1 159.33,49.14
X$9479 518 37 519 644 645 cell_1rw
* cell instance $9480 r0 *1 160.035,49.14
X$9480 520 37 521 644 645 cell_1rw
* cell instance $9481 r0 *1 160.74,49.14
X$9481 522 37 523 644 645 cell_1rw
* cell instance $9482 r0 *1 161.445,49.14
X$9482 524 37 525 644 645 cell_1rw
* cell instance $9483 r0 *1 162.15,49.14
X$9483 526 37 527 644 645 cell_1rw
* cell instance $9484 r0 *1 162.855,49.14
X$9484 528 37 529 644 645 cell_1rw
* cell instance $9485 r0 *1 163.56,49.14
X$9485 530 37 531 644 645 cell_1rw
* cell instance $9486 r0 *1 164.265,49.14
X$9486 532 37 533 644 645 cell_1rw
* cell instance $9487 r0 *1 164.97,49.14
X$9487 534 37 535 644 645 cell_1rw
* cell instance $9488 r0 *1 165.675,49.14
X$9488 536 37 537 644 645 cell_1rw
* cell instance $9489 r0 *1 166.38,49.14
X$9489 538 37 539 644 645 cell_1rw
* cell instance $9490 r0 *1 167.085,49.14
X$9490 540 37 541 644 645 cell_1rw
* cell instance $9491 r0 *1 167.79,49.14
X$9491 542 37 543 644 645 cell_1rw
* cell instance $9492 r0 *1 168.495,49.14
X$9492 544 37 545 644 645 cell_1rw
* cell instance $9493 r0 *1 169.2,49.14
X$9493 546 37 547 644 645 cell_1rw
* cell instance $9494 r0 *1 169.905,49.14
X$9494 548 37 549 644 645 cell_1rw
* cell instance $9495 r0 *1 170.61,49.14
X$9495 550 37 551 644 645 cell_1rw
* cell instance $9496 r0 *1 171.315,49.14
X$9496 552 37 553 644 645 cell_1rw
* cell instance $9497 r0 *1 172.02,49.14
X$9497 554 37 555 644 645 cell_1rw
* cell instance $9498 r0 *1 172.725,49.14
X$9498 556 37 557 644 645 cell_1rw
* cell instance $9499 r0 *1 173.43,49.14
X$9499 558 37 559 644 645 cell_1rw
* cell instance $9500 r0 *1 174.135,49.14
X$9500 560 37 561 644 645 cell_1rw
* cell instance $9501 r0 *1 174.84,49.14
X$9501 562 37 563 644 645 cell_1rw
* cell instance $9502 r0 *1 175.545,49.14
X$9502 564 37 565 644 645 cell_1rw
* cell instance $9503 r0 *1 176.25,49.14
X$9503 566 37 567 644 645 cell_1rw
* cell instance $9504 r0 *1 176.955,49.14
X$9504 568 37 569 644 645 cell_1rw
* cell instance $9505 r0 *1 177.66,49.14
X$9505 570 37 571 644 645 cell_1rw
* cell instance $9506 r0 *1 178.365,49.14
X$9506 572 37 573 644 645 cell_1rw
* cell instance $9507 r0 *1 179.07,49.14
X$9507 574 37 575 644 645 cell_1rw
* cell instance $9508 r0 *1 179.775,49.14
X$9508 576 37 577 644 645 cell_1rw
* cell instance $9509 r0 *1 180.48,49.14
X$9509 578 37 579 644 645 cell_1rw
* cell instance $9510 m0 *1 0.705,51.87
X$9510 67 38 68 644 645 cell_1rw
* cell instance $9511 m0 *1 0,51.87
X$9511 65 38 66 644 645 cell_1rw
* cell instance $9512 m0 *1 1.41,51.87
X$9512 69 38 70 644 645 cell_1rw
* cell instance $9513 m0 *1 2.115,51.87
X$9513 71 38 72 644 645 cell_1rw
* cell instance $9514 m0 *1 2.82,51.87
X$9514 73 38 74 644 645 cell_1rw
* cell instance $9515 m0 *1 3.525,51.87
X$9515 75 38 76 644 645 cell_1rw
* cell instance $9516 m0 *1 4.23,51.87
X$9516 77 38 78 644 645 cell_1rw
* cell instance $9517 m0 *1 4.935,51.87
X$9517 79 38 80 644 645 cell_1rw
* cell instance $9518 m0 *1 5.64,51.87
X$9518 81 38 82 644 645 cell_1rw
* cell instance $9519 m0 *1 6.345,51.87
X$9519 83 38 84 644 645 cell_1rw
* cell instance $9520 m0 *1 7.05,51.87
X$9520 85 38 86 644 645 cell_1rw
* cell instance $9521 m0 *1 7.755,51.87
X$9521 87 38 88 644 645 cell_1rw
* cell instance $9522 m0 *1 8.46,51.87
X$9522 89 38 90 644 645 cell_1rw
* cell instance $9523 m0 *1 9.165,51.87
X$9523 91 38 92 644 645 cell_1rw
* cell instance $9524 m0 *1 9.87,51.87
X$9524 93 38 94 644 645 cell_1rw
* cell instance $9525 m0 *1 10.575,51.87
X$9525 95 38 96 644 645 cell_1rw
* cell instance $9526 m0 *1 11.28,51.87
X$9526 97 38 98 644 645 cell_1rw
* cell instance $9527 m0 *1 11.985,51.87
X$9527 99 38 100 644 645 cell_1rw
* cell instance $9528 m0 *1 12.69,51.87
X$9528 101 38 102 644 645 cell_1rw
* cell instance $9529 m0 *1 13.395,51.87
X$9529 103 38 104 644 645 cell_1rw
* cell instance $9530 m0 *1 14.1,51.87
X$9530 105 38 106 644 645 cell_1rw
* cell instance $9531 m0 *1 14.805,51.87
X$9531 107 38 108 644 645 cell_1rw
* cell instance $9532 m0 *1 15.51,51.87
X$9532 109 38 110 644 645 cell_1rw
* cell instance $9533 m0 *1 16.215,51.87
X$9533 111 38 112 644 645 cell_1rw
* cell instance $9534 m0 *1 16.92,51.87
X$9534 113 38 114 644 645 cell_1rw
* cell instance $9535 m0 *1 17.625,51.87
X$9535 115 38 116 644 645 cell_1rw
* cell instance $9536 m0 *1 18.33,51.87
X$9536 117 38 118 644 645 cell_1rw
* cell instance $9537 m0 *1 19.035,51.87
X$9537 119 38 120 644 645 cell_1rw
* cell instance $9538 m0 *1 19.74,51.87
X$9538 121 38 122 644 645 cell_1rw
* cell instance $9539 m0 *1 20.445,51.87
X$9539 123 38 124 644 645 cell_1rw
* cell instance $9540 m0 *1 21.15,51.87
X$9540 125 38 126 644 645 cell_1rw
* cell instance $9541 m0 *1 21.855,51.87
X$9541 127 38 128 644 645 cell_1rw
* cell instance $9542 m0 *1 22.56,51.87
X$9542 129 38 130 644 645 cell_1rw
* cell instance $9543 m0 *1 23.265,51.87
X$9543 131 38 132 644 645 cell_1rw
* cell instance $9544 m0 *1 23.97,51.87
X$9544 133 38 134 644 645 cell_1rw
* cell instance $9545 m0 *1 24.675,51.87
X$9545 135 38 136 644 645 cell_1rw
* cell instance $9546 m0 *1 25.38,51.87
X$9546 137 38 138 644 645 cell_1rw
* cell instance $9547 m0 *1 26.085,51.87
X$9547 139 38 140 644 645 cell_1rw
* cell instance $9548 m0 *1 26.79,51.87
X$9548 141 38 142 644 645 cell_1rw
* cell instance $9549 m0 *1 27.495,51.87
X$9549 143 38 144 644 645 cell_1rw
* cell instance $9550 m0 *1 28.2,51.87
X$9550 145 38 146 644 645 cell_1rw
* cell instance $9551 m0 *1 28.905,51.87
X$9551 147 38 148 644 645 cell_1rw
* cell instance $9552 m0 *1 29.61,51.87
X$9552 149 38 150 644 645 cell_1rw
* cell instance $9553 m0 *1 30.315,51.87
X$9553 151 38 152 644 645 cell_1rw
* cell instance $9554 m0 *1 31.02,51.87
X$9554 153 38 154 644 645 cell_1rw
* cell instance $9555 m0 *1 31.725,51.87
X$9555 155 38 156 644 645 cell_1rw
* cell instance $9556 m0 *1 32.43,51.87
X$9556 157 38 158 644 645 cell_1rw
* cell instance $9557 m0 *1 33.135,51.87
X$9557 159 38 160 644 645 cell_1rw
* cell instance $9558 m0 *1 33.84,51.87
X$9558 161 38 162 644 645 cell_1rw
* cell instance $9559 m0 *1 34.545,51.87
X$9559 163 38 164 644 645 cell_1rw
* cell instance $9560 m0 *1 35.25,51.87
X$9560 165 38 166 644 645 cell_1rw
* cell instance $9561 m0 *1 35.955,51.87
X$9561 167 38 168 644 645 cell_1rw
* cell instance $9562 m0 *1 36.66,51.87
X$9562 169 38 170 644 645 cell_1rw
* cell instance $9563 m0 *1 37.365,51.87
X$9563 171 38 172 644 645 cell_1rw
* cell instance $9564 m0 *1 38.07,51.87
X$9564 173 38 174 644 645 cell_1rw
* cell instance $9565 m0 *1 38.775,51.87
X$9565 175 38 176 644 645 cell_1rw
* cell instance $9566 m0 *1 39.48,51.87
X$9566 177 38 178 644 645 cell_1rw
* cell instance $9567 m0 *1 40.185,51.87
X$9567 179 38 180 644 645 cell_1rw
* cell instance $9568 m0 *1 40.89,51.87
X$9568 181 38 182 644 645 cell_1rw
* cell instance $9569 m0 *1 41.595,51.87
X$9569 183 38 184 644 645 cell_1rw
* cell instance $9570 m0 *1 42.3,51.87
X$9570 185 38 186 644 645 cell_1rw
* cell instance $9571 m0 *1 43.005,51.87
X$9571 187 38 188 644 645 cell_1rw
* cell instance $9572 m0 *1 43.71,51.87
X$9572 189 38 190 644 645 cell_1rw
* cell instance $9573 m0 *1 44.415,51.87
X$9573 191 38 192 644 645 cell_1rw
* cell instance $9574 m0 *1 45.12,51.87
X$9574 193 38 194 644 645 cell_1rw
* cell instance $9575 m0 *1 45.825,51.87
X$9575 195 38 196 644 645 cell_1rw
* cell instance $9576 m0 *1 46.53,51.87
X$9576 197 38 198 644 645 cell_1rw
* cell instance $9577 m0 *1 47.235,51.87
X$9577 199 38 200 644 645 cell_1rw
* cell instance $9578 m0 *1 47.94,51.87
X$9578 201 38 202 644 645 cell_1rw
* cell instance $9579 m0 *1 48.645,51.87
X$9579 203 38 204 644 645 cell_1rw
* cell instance $9580 m0 *1 49.35,51.87
X$9580 205 38 206 644 645 cell_1rw
* cell instance $9581 m0 *1 50.055,51.87
X$9581 207 38 208 644 645 cell_1rw
* cell instance $9582 m0 *1 50.76,51.87
X$9582 209 38 210 644 645 cell_1rw
* cell instance $9583 m0 *1 51.465,51.87
X$9583 211 38 212 644 645 cell_1rw
* cell instance $9584 m0 *1 52.17,51.87
X$9584 213 38 214 644 645 cell_1rw
* cell instance $9585 m0 *1 52.875,51.87
X$9585 215 38 216 644 645 cell_1rw
* cell instance $9586 m0 *1 53.58,51.87
X$9586 217 38 218 644 645 cell_1rw
* cell instance $9587 m0 *1 54.285,51.87
X$9587 219 38 220 644 645 cell_1rw
* cell instance $9588 m0 *1 54.99,51.87
X$9588 221 38 222 644 645 cell_1rw
* cell instance $9589 m0 *1 55.695,51.87
X$9589 223 38 224 644 645 cell_1rw
* cell instance $9590 m0 *1 56.4,51.87
X$9590 225 38 226 644 645 cell_1rw
* cell instance $9591 m0 *1 57.105,51.87
X$9591 227 38 228 644 645 cell_1rw
* cell instance $9592 m0 *1 57.81,51.87
X$9592 229 38 230 644 645 cell_1rw
* cell instance $9593 m0 *1 58.515,51.87
X$9593 231 38 232 644 645 cell_1rw
* cell instance $9594 m0 *1 59.22,51.87
X$9594 233 38 234 644 645 cell_1rw
* cell instance $9595 m0 *1 59.925,51.87
X$9595 235 38 236 644 645 cell_1rw
* cell instance $9596 m0 *1 60.63,51.87
X$9596 237 38 238 644 645 cell_1rw
* cell instance $9597 m0 *1 61.335,51.87
X$9597 239 38 240 644 645 cell_1rw
* cell instance $9598 m0 *1 62.04,51.87
X$9598 241 38 242 644 645 cell_1rw
* cell instance $9599 m0 *1 62.745,51.87
X$9599 243 38 244 644 645 cell_1rw
* cell instance $9600 m0 *1 63.45,51.87
X$9600 245 38 246 644 645 cell_1rw
* cell instance $9601 m0 *1 64.155,51.87
X$9601 247 38 248 644 645 cell_1rw
* cell instance $9602 m0 *1 64.86,51.87
X$9602 249 38 250 644 645 cell_1rw
* cell instance $9603 m0 *1 65.565,51.87
X$9603 251 38 252 644 645 cell_1rw
* cell instance $9604 m0 *1 66.27,51.87
X$9604 253 38 254 644 645 cell_1rw
* cell instance $9605 m0 *1 66.975,51.87
X$9605 255 38 256 644 645 cell_1rw
* cell instance $9606 m0 *1 67.68,51.87
X$9606 257 38 258 644 645 cell_1rw
* cell instance $9607 m0 *1 68.385,51.87
X$9607 259 38 260 644 645 cell_1rw
* cell instance $9608 m0 *1 69.09,51.87
X$9608 261 38 262 644 645 cell_1rw
* cell instance $9609 m0 *1 69.795,51.87
X$9609 263 38 264 644 645 cell_1rw
* cell instance $9610 m0 *1 70.5,51.87
X$9610 265 38 266 644 645 cell_1rw
* cell instance $9611 m0 *1 71.205,51.87
X$9611 267 38 268 644 645 cell_1rw
* cell instance $9612 m0 *1 71.91,51.87
X$9612 269 38 270 644 645 cell_1rw
* cell instance $9613 m0 *1 72.615,51.87
X$9613 271 38 272 644 645 cell_1rw
* cell instance $9614 m0 *1 73.32,51.87
X$9614 273 38 274 644 645 cell_1rw
* cell instance $9615 m0 *1 74.025,51.87
X$9615 275 38 276 644 645 cell_1rw
* cell instance $9616 m0 *1 74.73,51.87
X$9616 277 38 278 644 645 cell_1rw
* cell instance $9617 m0 *1 75.435,51.87
X$9617 279 38 280 644 645 cell_1rw
* cell instance $9618 m0 *1 76.14,51.87
X$9618 281 38 282 644 645 cell_1rw
* cell instance $9619 m0 *1 76.845,51.87
X$9619 283 38 284 644 645 cell_1rw
* cell instance $9620 m0 *1 77.55,51.87
X$9620 285 38 286 644 645 cell_1rw
* cell instance $9621 m0 *1 78.255,51.87
X$9621 287 38 288 644 645 cell_1rw
* cell instance $9622 m0 *1 78.96,51.87
X$9622 289 38 290 644 645 cell_1rw
* cell instance $9623 m0 *1 79.665,51.87
X$9623 291 38 292 644 645 cell_1rw
* cell instance $9624 m0 *1 80.37,51.87
X$9624 293 38 294 644 645 cell_1rw
* cell instance $9625 m0 *1 81.075,51.87
X$9625 295 38 296 644 645 cell_1rw
* cell instance $9626 m0 *1 81.78,51.87
X$9626 297 38 298 644 645 cell_1rw
* cell instance $9627 m0 *1 82.485,51.87
X$9627 299 38 300 644 645 cell_1rw
* cell instance $9628 m0 *1 83.19,51.87
X$9628 301 38 302 644 645 cell_1rw
* cell instance $9629 m0 *1 83.895,51.87
X$9629 303 38 304 644 645 cell_1rw
* cell instance $9630 m0 *1 84.6,51.87
X$9630 305 38 306 644 645 cell_1rw
* cell instance $9631 m0 *1 85.305,51.87
X$9631 307 38 308 644 645 cell_1rw
* cell instance $9632 m0 *1 86.01,51.87
X$9632 309 38 310 644 645 cell_1rw
* cell instance $9633 m0 *1 86.715,51.87
X$9633 311 38 312 644 645 cell_1rw
* cell instance $9634 m0 *1 87.42,51.87
X$9634 313 38 314 644 645 cell_1rw
* cell instance $9635 m0 *1 88.125,51.87
X$9635 315 38 316 644 645 cell_1rw
* cell instance $9636 m0 *1 88.83,51.87
X$9636 317 38 318 644 645 cell_1rw
* cell instance $9637 m0 *1 89.535,51.87
X$9637 319 38 320 644 645 cell_1rw
* cell instance $9638 m0 *1 90.24,51.87
X$9638 321 38 323 644 645 cell_1rw
* cell instance $9639 m0 *1 90.945,51.87
X$9639 324 38 325 644 645 cell_1rw
* cell instance $9640 m0 *1 91.65,51.87
X$9640 326 38 327 644 645 cell_1rw
* cell instance $9641 m0 *1 92.355,51.87
X$9641 328 38 329 644 645 cell_1rw
* cell instance $9642 m0 *1 93.06,51.87
X$9642 330 38 331 644 645 cell_1rw
* cell instance $9643 m0 *1 93.765,51.87
X$9643 332 38 333 644 645 cell_1rw
* cell instance $9644 m0 *1 94.47,51.87
X$9644 334 38 335 644 645 cell_1rw
* cell instance $9645 m0 *1 95.175,51.87
X$9645 336 38 337 644 645 cell_1rw
* cell instance $9646 m0 *1 95.88,51.87
X$9646 338 38 339 644 645 cell_1rw
* cell instance $9647 m0 *1 96.585,51.87
X$9647 340 38 341 644 645 cell_1rw
* cell instance $9648 m0 *1 97.29,51.87
X$9648 342 38 343 644 645 cell_1rw
* cell instance $9649 m0 *1 97.995,51.87
X$9649 344 38 345 644 645 cell_1rw
* cell instance $9650 m0 *1 98.7,51.87
X$9650 346 38 347 644 645 cell_1rw
* cell instance $9651 m0 *1 99.405,51.87
X$9651 348 38 349 644 645 cell_1rw
* cell instance $9652 m0 *1 100.11,51.87
X$9652 350 38 351 644 645 cell_1rw
* cell instance $9653 m0 *1 100.815,51.87
X$9653 352 38 353 644 645 cell_1rw
* cell instance $9654 m0 *1 101.52,51.87
X$9654 354 38 355 644 645 cell_1rw
* cell instance $9655 m0 *1 102.225,51.87
X$9655 356 38 357 644 645 cell_1rw
* cell instance $9656 m0 *1 102.93,51.87
X$9656 358 38 359 644 645 cell_1rw
* cell instance $9657 m0 *1 103.635,51.87
X$9657 360 38 361 644 645 cell_1rw
* cell instance $9658 m0 *1 104.34,51.87
X$9658 362 38 363 644 645 cell_1rw
* cell instance $9659 m0 *1 105.045,51.87
X$9659 364 38 365 644 645 cell_1rw
* cell instance $9660 m0 *1 105.75,51.87
X$9660 366 38 367 644 645 cell_1rw
* cell instance $9661 m0 *1 106.455,51.87
X$9661 368 38 369 644 645 cell_1rw
* cell instance $9662 m0 *1 107.16,51.87
X$9662 370 38 371 644 645 cell_1rw
* cell instance $9663 m0 *1 107.865,51.87
X$9663 372 38 373 644 645 cell_1rw
* cell instance $9664 m0 *1 108.57,51.87
X$9664 374 38 375 644 645 cell_1rw
* cell instance $9665 m0 *1 109.275,51.87
X$9665 376 38 377 644 645 cell_1rw
* cell instance $9666 m0 *1 109.98,51.87
X$9666 378 38 379 644 645 cell_1rw
* cell instance $9667 m0 *1 110.685,51.87
X$9667 380 38 381 644 645 cell_1rw
* cell instance $9668 m0 *1 111.39,51.87
X$9668 382 38 383 644 645 cell_1rw
* cell instance $9669 m0 *1 112.095,51.87
X$9669 384 38 385 644 645 cell_1rw
* cell instance $9670 m0 *1 112.8,51.87
X$9670 386 38 387 644 645 cell_1rw
* cell instance $9671 m0 *1 113.505,51.87
X$9671 388 38 389 644 645 cell_1rw
* cell instance $9672 m0 *1 114.21,51.87
X$9672 390 38 391 644 645 cell_1rw
* cell instance $9673 m0 *1 114.915,51.87
X$9673 392 38 393 644 645 cell_1rw
* cell instance $9674 m0 *1 115.62,51.87
X$9674 394 38 395 644 645 cell_1rw
* cell instance $9675 m0 *1 116.325,51.87
X$9675 396 38 397 644 645 cell_1rw
* cell instance $9676 m0 *1 117.03,51.87
X$9676 398 38 399 644 645 cell_1rw
* cell instance $9677 m0 *1 117.735,51.87
X$9677 400 38 401 644 645 cell_1rw
* cell instance $9678 m0 *1 118.44,51.87
X$9678 402 38 403 644 645 cell_1rw
* cell instance $9679 m0 *1 119.145,51.87
X$9679 404 38 405 644 645 cell_1rw
* cell instance $9680 m0 *1 119.85,51.87
X$9680 406 38 407 644 645 cell_1rw
* cell instance $9681 m0 *1 120.555,51.87
X$9681 408 38 409 644 645 cell_1rw
* cell instance $9682 m0 *1 121.26,51.87
X$9682 410 38 411 644 645 cell_1rw
* cell instance $9683 m0 *1 121.965,51.87
X$9683 412 38 413 644 645 cell_1rw
* cell instance $9684 m0 *1 122.67,51.87
X$9684 414 38 415 644 645 cell_1rw
* cell instance $9685 m0 *1 123.375,51.87
X$9685 416 38 417 644 645 cell_1rw
* cell instance $9686 m0 *1 124.08,51.87
X$9686 418 38 419 644 645 cell_1rw
* cell instance $9687 m0 *1 124.785,51.87
X$9687 420 38 421 644 645 cell_1rw
* cell instance $9688 m0 *1 125.49,51.87
X$9688 422 38 423 644 645 cell_1rw
* cell instance $9689 m0 *1 126.195,51.87
X$9689 424 38 425 644 645 cell_1rw
* cell instance $9690 m0 *1 126.9,51.87
X$9690 426 38 427 644 645 cell_1rw
* cell instance $9691 m0 *1 127.605,51.87
X$9691 428 38 429 644 645 cell_1rw
* cell instance $9692 m0 *1 128.31,51.87
X$9692 430 38 431 644 645 cell_1rw
* cell instance $9693 m0 *1 129.015,51.87
X$9693 432 38 433 644 645 cell_1rw
* cell instance $9694 m0 *1 129.72,51.87
X$9694 434 38 435 644 645 cell_1rw
* cell instance $9695 m0 *1 130.425,51.87
X$9695 436 38 437 644 645 cell_1rw
* cell instance $9696 m0 *1 131.13,51.87
X$9696 438 38 439 644 645 cell_1rw
* cell instance $9697 m0 *1 131.835,51.87
X$9697 440 38 441 644 645 cell_1rw
* cell instance $9698 m0 *1 132.54,51.87
X$9698 442 38 443 644 645 cell_1rw
* cell instance $9699 m0 *1 133.245,51.87
X$9699 444 38 445 644 645 cell_1rw
* cell instance $9700 m0 *1 133.95,51.87
X$9700 446 38 447 644 645 cell_1rw
* cell instance $9701 m0 *1 134.655,51.87
X$9701 448 38 449 644 645 cell_1rw
* cell instance $9702 m0 *1 135.36,51.87
X$9702 450 38 451 644 645 cell_1rw
* cell instance $9703 m0 *1 136.065,51.87
X$9703 452 38 453 644 645 cell_1rw
* cell instance $9704 m0 *1 136.77,51.87
X$9704 454 38 455 644 645 cell_1rw
* cell instance $9705 m0 *1 137.475,51.87
X$9705 456 38 457 644 645 cell_1rw
* cell instance $9706 m0 *1 138.18,51.87
X$9706 458 38 459 644 645 cell_1rw
* cell instance $9707 m0 *1 138.885,51.87
X$9707 460 38 461 644 645 cell_1rw
* cell instance $9708 m0 *1 139.59,51.87
X$9708 462 38 463 644 645 cell_1rw
* cell instance $9709 m0 *1 140.295,51.87
X$9709 464 38 465 644 645 cell_1rw
* cell instance $9710 m0 *1 141,51.87
X$9710 466 38 467 644 645 cell_1rw
* cell instance $9711 m0 *1 141.705,51.87
X$9711 468 38 469 644 645 cell_1rw
* cell instance $9712 m0 *1 142.41,51.87
X$9712 470 38 471 644 645 cell_1rw
* cell instance $9713 m0 *1 143.115,51.87
X$9713 472 38 473 644 645 cell_1rw
* cell instance $9714 m0 *1 143.82,51.87
X$9714 474 38 475 644 645 cell_1rw
* cell instance $9715 m0 *1 144.525,51.87
X$9715 476 38 477 644 645 cell_1rw
* cell instance $9716 m0 *1 145.23,51.87
X$9716 478 38 479 644 645 cell_1rw
* cell instance $9717 m0 *1 145.935,51.87
X$9717 480 38 481 644 645 cell_1rw
* cell instance $9718 m0 *1 146.64,51.87
X$9718 482 38 483 644 645 cell_1rw
* cell instance $9719 m0 *1 147.345,51.87
X$9719 484 38 485 644 645 cell_1rw
* cell instance $9720 m0 *1 148.05,51.87
X$9720 486 38 487 644 645 cell_1rw
* cell instance $9721 m0 *1 148.755,51.87
X$9721 488 38 489 644 645 cell_1rw
* cell instance $9722 m0 *1 149.46,51.87
X$9722 490 38 491 644 645 cell_1rw
* cell instance $9723 m0 *1 150.165,51.87
X$9723 492 38 493 644 645 cell_1rw
* cell instance $9724 m0 *1 150.87,51.87
X$9724 494 38 495 644 645 cell_1rw
* cell instance $9725 m0 *1 151.575,51.87
X$9725 496 38 497 644 645 cell_1rw
* cell instance $9726 m0 *1 152.28,51.87
X$9726 498 38 499 644 645 cell_1rw
* cell instance $9727 m0 *1 152.985,51.87
X$9727 500 38 501 644 645 cell_1rw
* cell instance $9728 m0 *1 153.69,51.87
X$9728 502 38 503 644 645 cell_1rw
* cell instance $9729 m0 *1 154.395,51.87
X$9729 504 38 505 644 645 cell_1rw
* cell instance $9730 m0 *1 155.1,51.87
X$9730 506 38 507 644 645 cell_1rw
* cell instance $9731 m0 *1 155.805,51.87
X$9731 508 38 509 644 645 cell_1rw
* cell instance $9732 m0 *1 156.51,51.87
X$9732 510 38 511 644 645 cell_1rw
* cell instance $9733 m0 *1 157.215,51.87
X$9733 512 38 513 644 645 cell_1rw
* cell instance $9734 m0 *1 157.92,51.87
X$9734 514 38 515 644 645 cell_1rw
* cell instance $9735 m0 *1 158.625,51.87
X$9735 516 38 517 644 645 cell_1rw
* cell instance $9736 m0 *1 159.33,51.87
X$9736 518 38 519 644 645 cell_1rw
* cell instance $9737 m0 *1 160.035,51.87
X$9737 520 38 521 644 645 cell_1rw
* cell instance $9738 m0 *1 160.74,51.87
X$9738 522 38 523 644 645 cell_1rw
* cell instance $9739 m0 *1 161.445,51.87
X$9739 524 38 525 644 645 cell_1rw
* cell instance $9740 m0 *1 162.15,51.87
X$9740 526 38 527 644 645 cell_1rw
* cell instance $9741 m0 *1 162.855,51.87
X$9741 528 38 529 644 645 cell_1rw
* cell instance $9742 m0 *1 163.56,51.87
X$9742 530 38 531 644 645 cell_1rw
* cell instance $9743 m0 *1 164.265,51.87
X$9743 532 38 533 644 645 cell_1rw
* cell instance $9744 m0 *1 164.97,51.87
X$9744 534 38 535 644 645 cell_1rw
* cell instance $9745 m0 *1 165.675,51.87
X$9745 536 38 537 644 645 cell_1rw
* cell instance $9746 m0 *1 166.38,51.87
X$9746 538 38 539 644 645 cell_1rw
* cell instance $9747 m0 *1 167.085,51.87
X$9747 540 38 541 644 645 cell_1rw
* cell instance $9748 m0 *1 167.79,51.87
X$9748 542 38 543 644 645 cell_1rw
* cell instance $9749 m0 *1 168.495,51.87
X$9749 544 38 545 644 645 cell_1rw
* cell instance $9750 m0 *1 169.2,51.87
X$9750 546 38 547 644 645 cell_1rw
* cell instance $9751 m0 *1 169.905,51.87
X$9751 548 38 549 644 645 cell_1rw
* cell instance $9752 m0 *1 170.61,51.87
X$9752 550 38 551 644 645 cell_1rw
* cell instance $9753 m0 *1 171.315,51.87
X$9753 552 38 553 644 645 cell_1rw
* cell instance $9754 m0 *1 172.02,51.87
X$9754 554 38 555 644 645 cell_1rw
* cell instance $9755 m0 *1 172.725,51.87
X$9755 556 38 557 644 645 cell_1rw
* cell instance $9756 m0 *1 173.43,51.87
X$9756 558 38 559 644 645 cell_1rw
* cell instance $9757 m0 *1 174.135,51.87
X$9757 560 38 561 644 645 cell_1rw
* cell instance $9758 m0 *1 174.84,51.87
X$9758 562 38 563 644 645 cell_1rw
* cell instance $9759 m0 *1 175.545,51.87
X$9759 564 38 565 644 645 cell_1rw
* cell instance $9760 m0 *1 176.25,51.87
X$9760 566 38 567 644 645 cell_1rw
* cell instance $9761 m0 *1 176.955,51.87
X$9761 568 38 569 644 645 cell_1rw
* cell instance $9762 m0 *1 177.66,51.87
X$9762 570 38 571 644 645 cell_1rw
* cell instance $9763 m0 *1 178.365,51.87
X$9763 572 38 573 644 645 cell_1rw
* cell instance $9764 m0 *1 179.07,51.87
X$9764 574 38 575 644 645 cell_1rw
* cell instance $9765 m0 *1 179.775,51.87
X$9765 576 38 577 644 645 cell_1rw
* cell instance $9766 m0 *1 180.48,51.87
X$9766 578 38 579 644 645 cell_1rw
* cell instance $9767 m0 *1 0.705,54.6
X$9767 67 39 68 644 645 cell_1rw
* cell instance $9768 m0 *1 0,54.6
X$9768 65 39 66 644 645 cell_1rw
* cell instance $9769 m0 *1 1.41,54.6
X$9769 69 39 70 644 645 cell_1rw
* cell instance $9770 m0 *1 2.115,54.6
X$9770 71 39 72 644 645 cell_1rw
* cell instance $9771 m0 *1 2.82,54.6
X$9771 73 39 74 644 645 cell_1rw
* cell instance $9772 m0 *1 3.525,54.6
X$9772 75 39 76 644 645 cell_1rw
* cell instance $9773 m0 *1 4.23,54.6
X$9773 77 39 78 644 645 cell_1rw
* cell instance $9774 m0 *1 4.935,54.6
X$9774 79 39 80 644 645 cell_1rw
* cell instance $9775 m0 *1 5.64,54.6
X$9775 81 39 82 644 645 cell_1rw
* cell instance $9776 m0 *1 6.345,54.6
X$9776 83 39 84 644 645 cell_1rw
* cell instance $9777 m0 *1 7.05,54.6
X$9777 85 39 86 644 645 cell_1rw
* cell instance $9778 m0 *1 7.755,54.6
X$9778 87 39 88 644 645 cell_1rw
* cell instance $9779 m0 *1 8.46,54.6
X$9779 89 39 90 644 645 cell_1rw
* cell instance $9780 m0 *1 9.165,54.6
X$9780 91 39 92 644 645 cell_1rw
* cell instance $9781 m0 *1 9.87,54.6
X$9781 93 39 94 644 645 cell_1rw
* cell instance $9782 m0 *1 10.575,54.6
X$9782 95 39 96 644 645 cell_1rw
* cell instance $9783 m0 *1 11.28,54.6
X$9783 97 39 98 644 645 cell_1rw
* cell instance $9784 m0 *1 11.985,54.6
X$9784 99 39 100 644 645 cell_1rw
* cell instance $9785 m0 *1 12.69,54.6
X$9785 101 39 102 644 645 cell_1rw
* cell instance $9786 m0 *1 13.395,54.6
X$9786 103 39 104 644 645 cell_1rw
* cell instance $9787 m0 *1 14.1,54.6
X$9787 105 39 106 644 645 cell_1rw
* cell instance $9788 m0 *1 14.805,54.6
X$9788 107 39 108 644 645 cell_1rw
* cell instance $9789 m0 *1 15.51,54.6
X$9789 109 39 110 644 645 cell_1rw
* cell instance $9790 m0 *1 16.215,54.6
X$9790 111 39 112 644 645 cell_1rw
* cell instance $9791 m0 *1 16.92,54.6
X$9791 113 39 114 644 645 cell_1rw
* cell instance $9792 m0 *1 17.625,54.6
X$9792 115 39 116 644 645 cell_1rw
* cell instance $9793 m0 *1 18.33,54.6
X$9793 117 39 118 644 645 cell_1rw
* cell instance $9794 m0 *1 19.035,54.6
X$9794 119 39 120 644 645 cell_1rw
* cell instance $9795 m0 *1 19.74,54.6
X$9795 121 39 122 644 645 cell_1rw
* cell instance $9796 m0 *1 20.445,54.6
X$9796 123 39 124 644 645 cell_1rw
* cell instance $9797 m0 *1 21.15,54.6
X$9797 125 39 126 644 645 cell_1rw
* cell instance $9798 m0 *1 21.855,54.6
X$9798 127 39 128 644 645 cell_1rw
* cell instance $9799 m0 *1 22.56,54.6
X$9799 129 39 130 644 645 cell_1rw
* cell instance $9800 m0 *1 23.265,54.6
X$9800 131 39 132 644 645 cell_1rw
* cell instance $9801 m0 *1 23.97,54.6
X$9801 133 39 134 644 645 cell_1rw
* cell instance $9802 m0 *1 24.675,54.6
X$9802 135 39 136 644 645 cell_1rw
* cell instance $9803 m0 *1 25.38,54.6
X$9803 137 39 138 644 645 cell_1rw
* cell instance $9804 m0 *1 26.085,54.6
X$9804 139 39 140 644 645 cell_1rw
* cell instance $9805 m0 *1 26.79,54.6
X$9805 141 39 142 644 645 cell_1rw
* cell instance $9806 m0 *1 27.495,54.6
X$9806 143 39 144 644 645 cell_1rw
* cell instance $9807 m0 *1 28.2,54.6
X$9807 145 39 146 644 645 cell_1rw
* cell instance $9808 m0 *1 28.905,54.6
X$9808 147 39 148 644 645 cell_1rw
* cell instance $9809 m0 *1 29.61,54.6
X$9809 149 39 150 644 645 cell_1rw
* cell instance $9810 m0 *1 30.315,54.6
X$9810 151 39 152 644 645 cell_1rw
* cell instance $9811 m0 *1 31.02,54.6
X$9811 153 39 154 644 645 cell_1rw
* cell instance $9812 m0 *1 31.725,54.6
X$9812 155 39 156 644 645 cell_1rw
* cell instance $9813 m0 *1 32.43,54.6
X$9813 157 39 158 644 645 cell_1rw
* cell instance $9814 m0 *1 33.135,54.6
X$9814 159 39 160 644 645 cell_1rw
* cell instance $9815 m0 *1 33.84,54.6
X$9815 161 39 162 644 645 cell_1rw
* cell instance $9816 m0 *1 34.545,54.6
X$9816 163 39 164 644 645 cell_1rw
* cell instance $9817 m0 *1 35.25,54.6
X$9817 165 39 166 644 645 cell_1rw
* cell instance $9818 m0 *1 35.955,54.6
X$9818 167 39 168 644 645 cell_1rw
* cell instance $9819 m0 *1 36.66,54.6
X$9819 169 39 170 644 645 cell_1rw
* cell instance $9820 m0 *1 37.365,54.6
X$9820 171 39 172 644 645 cell_1rw
* cell instance $9821 m0 *1 38.07,54.6
X$9821 173 39 174 644 645 cell_1rw
* cell instance $9822 m0 *1 38.775,54.6
X$9822 175 39 176 644 645 cell_1rw
* cell instance $9823 m0 *1 39.48,54.6
X$9823 177 39 178 644 645 cell_1rw
* cell instance $9824 m0 *1 40.185,54.6
X$9824 179 39 180 644 645 cell_1rw
* cell instance $9825 m0 *1 40.89,54.6
X$9825 181 39 182 644 645 cell_1rw
* cell instance $9826 m0 *1 41.595,54.6
X$9826 183 39 184 644 645 cell_1rw
* cell instance $9827 m0 *1 42.3,54.6
X$9827 185 39 186 644 645 cell_1rw
* cell instance $9828 m0 *1 43.005,54.6
X$9828 187 39 188 644 645 cell_1rw
* cell instance $9829 m0 *1 43.71,54.6
X$9829 189 39 190 644 645 cell_1rw
* cell instance $9830 m0 *1 44.415,54.6
X$9830 191 39 192 644 645 cell_1rw
* cell instance $9831 m0 *1 45.12,54.6
X$9831 193 39 194 644 645 cell_1rw
* cell instance $9832 m0 *1 45.825,54.6
X$9832 195 39 196 644 645 cell_1rw
* cell instance $9833 m0 *1 46.53,54.6
X$9833 197 39 198 644 645 cell_1rw
* cell instance $9834 m0 *1 47.235,54.6
X$9834 199 39 200 644 645 cell_1rw
* cell instance $9835 m0 *1 47.94,54.6
X$9835 201 39 202 644 645 cell_1rw
* cell instance $9836 m0 *1 48.645,54.6
X$9836 203 39 204 644 645 cell_1rw
* cell instance $9837 m0 *1 49.35,54.6
X$9837 205 39 206 644 645 cell_1rw
* cell instance $9838 m0 *1 50.055,54.6
X$9838 207 39 208 644 645 cell_1rw
* cell instance $9839 m0 *1 50.76,54.6
X$9839 209 39 210 644 645 cell_1rw
* cell instance $9840 m0 *1 51.465,54.6
X$9840 211 39 212 644 645 cell_1rw
* cell instance $9841 m0 *1 52.17,54.6
X$9841 213 39 214 644 645 cell_1rw
* cell instance $9842 m0 *1 52.875,54.6
X$9842 215 39 216 644 645 cell_1rw
* cell instance $9843 m0 *1 53.58,54.6
X$9843 217 39 218 644 645 cell_1rw
* cell instance $9844 m0 *1 54.285,54.6
X$9844 219 39 220 644 645 cell_1rw
* cell instance $9845 m0 *1 54.99,54.6
X$9845 221 39 222 644 645 cell_1rw
* cell instance $9846 m0 *1 55.695,54.6
X$9846 223 39 224 644 645 cell_1rw
* cell instance $9847 m0 *1 56.4,54.6
X$9847 225 39 226 644 645 cell_1rw
* cell instance $9848 m0 *1 57.105,54.6
X$9848 227 39 228 644 645 cell_1rw
* cell instance $9849 m0 *1 57.81,54.6
X$9849 229 39 230 644 645 cell_1rw
* cell instance $9850 m0 *1 58.515,54.6
X$9850 231 39 232 644 645 cell_1rw
* cell instance $9851 m0 *1 59.22,54.6
X$9851 233 39 234 644 645 cell_1rw
* cell instance $9852 m0 *1 59.925,54.6
X$9852 235 39 236 644 645 cell_1rw
* cell instance $9853 m0 *1 60.63,54.6
X$9853 237 39 238 644 645 cell_1rw
* cell instance $9854 m0 *1 61.335,54.6
X$9854 239 39 240 644 645 cell_1rw
* cell instance $9855 m0 *1 62.04,54.6
X$9855 241 39 242 644 645 cell_1rw
* cell instance $9856 m0 *1 62.745,54.6
X$9856 243 39 244 644 645 cell_1rw
* cell instance $9857 m0 *1 63.45,54.6
X$9857 245 39 246 644 645 cell_1rw
* cell instance $9858 m0 *1 64.155,54.6
X$9858 247 39 248 644 645 cell_1rw
* cell instance $9859 m0 *1 64.86,54.6
X$9859 249 39 250 644 645 cell_1rw
* cell instance $9860 m0 *1 65.565,54.6
X$9860 251 39 252 644 645 cell_1rw
* cell instance $9861 m0 *1 66.27,54.6
X$9861 253 39 254 644 645 cell_1rw
* cell instance $9862 m0 *1 66.975,54.6
X$9862 255 39 256 644 645 cell_1rw
* cell instance $9863 m0 *1 67.68,54.6
X$9863 257 39 258 644 645 cell_1rw
* cell instance $9864 m0 *1 68.385,54.6
X$9864 259 39 260 644 645 cell_1rw
* cell instance $9865 m0 *1 69.09,54.6
X$9865 261 39 262 644 645 cell_1rw
* cell instance $9866 m0 *1 69.795,54.6
X$9866 263 39 264 644 645 cell_1rw
* cell instance $9867 m0 *1 70.5,54.6
X$9867 265 39 266 644 645 cell_1rw
* cell instance $9868 m0 *1 71.205,54.6
X$9868 267 39 268 644 645 cell_1rw
* cell instance $9869 m0 *1 71.91,54.6
X$9869 269 39 270 644 645 cell_1rw
* cell instance $9870 m0 *1 72.615,54.6
X$9870 271 39 272 644 645 cell_1rw
* cell instance $9871 m0 *1 73.32,54.6
X$9871 273 39 274 644 645 cell_1rw
* cell instance $9872 m0 *1 74.025,54.6
X$9872 275 39 276 644 645 cell_1rw
* cell instance $9873 m0 *1 74.73,54.6
X$9873 277 39 278 644 645 cell_1rw
* cell instance $9874 m0 *1 75.435,54.6
X$9874 279 39 280 644 645 cell_1rw
* cell instance $9875 m0 *1 76.14,54.6
X$9875 281 39 282 644 645 cell_1rw
* cell instance $9876 m0 *1 76.845,54.6
X$9876 283 39 284 644 645 cell_1rw
* cell instance $9877 m0 *1 77.55,54.6
X$9877 285 39 286 644 645 cell_1rw
* cell instance $9878 m0 *1 78.255,54.6
X$9878 287 39 288 644 645 cell_1rw
* cell instance $9879 m0 *1 78.96,54.6
X$9879 289 39 290 644 645 cell_1rw
* cell instance $9880 m0 *1 79.665,54.6
X$9880 291 39 292 644 645 cell_1rw
* cell instance $9881 m0 *1 80.37,54.6
X$9881 293 39 294 644 645 cell_1rw
* cell instance $9882 m0 *1 81.075,54.6
X$9882 295 39 296 644 645 cell_1rw
* cell instance $9883 m0 *1 81.78,54.6
X$9883 297 39 298 644 645 cell_1rw
* cell instance $9884 m0 *1 82.485,54.6
X$9884 299 39 300 644 645 cell_1rw
* cell instance $9885 m0 *1 83.19,54.6
X$9885 301 39 302 644 645 cell_1rw
* cell instance $9886 m0 *1 83.895,54.6
X$9886 303 39 304 644 645 cell_1rw
* cell instance $9887 m0 *1 84.6,54.6
X$9887 305 39 306 644 645 cell_1rw
* cell instance $9888 m0 *1 85.305,54.6
X$9888 307 39 308 644 645 cell_1rw
* cell instance $9889 m0 *1 86.01,54.6
X$9889 309 39 310 644 645 cell_1rw
* cell instance $9890 m0 *1 86.715,54.6
X$9890 311 39 312 644 645 cell_1rw
* cell instance $9891 m0 *1 87.42,54.6
X$9891 313 39 314 644 645 cell_1rw
* cell instance $9892 m0 *1 88.125,54.6
X$9892 315 39 316 644 645 cell_1rw
* cell instance $9893 m0 *1 88.83,54.6
X$9893 317 39 318 644 645 cell_1rw
* cell instance $9894 m0 *1 89.535,54.6
X$9894 319 39 320 644 645 cell_1rw
* cell instance $9895 m0 *1 90.24,54.6
X$9895 321 39 323 644 645 cell_1rw
* cell instance $9896 m0 *1 90.945,54.6
X$9896 324 39 325 644 645 cell_1rw
* cell instance $9897 m0 *1 91.65,54.6
X$9897 326 39 327 644 645 cell_1rw
* cell instance $9898 m0 *1 92.355,54.6
X$9898 328 39 329 644 645 cell_1rw
* cell instance $9899 m0 *1 93.06,54.6
X$9899 330 39 331 644 645 cell_1rw
* cell instance $9900 m0 *1 93.765,54.6
X$9900 332 39 333 644 645 cell_1rw
* cell instance $9901 m0 *1 94.47,54.6
X$9901 334 39 335 644 645 cell_1rw
* cell instance $9902 m0 *1 95.175,54.6
X$9902 336 39 337 644 645 cell_1rw
* cell instance $9903 m0 *1 95.88,54.6
X$9903 338 39 339 644 645 cell_1rw
* cell instance $9904 m0 *1 96.585,54.6
X$9904 340 39 341 644 645 cell_1rw
* cell instance $9905 m0 *1 97.29,54.6
X$9905 342 39 343 644 645 cell_1rw
* cell instance $9906 m0 *1 97.995,54.6
X$9906 344 39 345 644 645 cell_1rw
* cell instance $9907 m0 *1 98.7,54.6
X$9907 346 39 347 644 645 cell_1rw
* cell instance $9908 m0 *1 99.405,54.6
X$9908 348 39 349 644 645 cell_1rw
* cell instance $9909 m0 *1 100.11,54.6
X$9909 350 39 351 644 645 cell_1rw
* cell instance $9910 m0 *1 100.815,54.6
X$9910 352 39 353 644 645 cell_1rw
* cell instance $9911 m0 *1 101.52,54.6
X$9911 354 39 355 644 645 cell_1rw
* cell instance $9912 m0 *1 102.225,54.6
X$9912 356 39 357 644 645 cell_1rw
* cell instance $9913 m0 *1 102.93,54.6
X$9913 358 39 359 644 645 cell_1rw
* cell instance $9914 m0 *1 103.635,54.6
X$9914 360 39 361 644 645 cell_1rw
* cell instance $9915 m0 *1 104.34,54.6
X$9915 362 39 363 644 645 cell_1rw
* cell instance $9916 m0 *1 105.045,54.6
X$9916 364 39 365 644 645 cell_1rw
* cell instance $9917 m0 *1 105.75,54.6
X$9917 366 39 367 644 645 cell_1rw
* cell instance $9918 m0 *1 106.455,54.6
X$9918 368 39 369 644 645 cell_1rw
* cell instance $9919 m0 *1 107.16,54.6
X$9919 370 39 371 644 645 cell_1rw
* cell instance $9920 m0 *1 107.865,54.6
X$9920 372 39 373 644 645 cell_1rw
* cell instance $9921 m0 *1 108.57,54.6
X$9921 374 39 375 644 645 cell_1rw
* cell instance $9922 m0 *1 109.275,54.6
X$9922 376 39 377 644 645 cell_1rw
* cell instance $9923 m0 *1 109.98,54.6
X$9923 378 39 379 644 645 cell_1rw
* cell instance $9924 m0 *1 110.685,54.6
X$9924 380 39 381 644 645 cell_1rw
* cell instance $9925 m0 *1 111.39,54.6
X$9925 382 39 383 644 645 cell_1rw
* cell instance $9926 m0 *1 112.095,54.6
X$9926 384 39 385 644 645 cell_1rw
* cell instance $9927 m0 *1 112.8,54.6
X$9927 386 39 387 644 645 cell_1rw
* cell instance $9928 m0 *1 113.505,54.6
X$9928 388 39 389 644 645 cell_1rw
* cell instance $9929 m0 *1 114.21,54.6
X$9929 390 39 391 644 645 cell_1rw
* cell instance $9930 m0 *1 114.915,54.6
X$9930 392 39 393 644 645 cell_1rw
* cell instance $9931 m0 *1 115.62,54.6
X$9931 394 39 395 644 645 cell_1rw
* cell instance $9932 m0 *1 116.325,54.6
X$9932 396 39 397 644 645 cell_1rw
* cell instance $9933 m0 *1 117.03,54.6
X$9933 398 39 399 644 645 cell_1rw
* cell instance $9934 m0 *1 117.735,54.6
X$9934 400 39 401 644 645 cell_1rw
* cell instance $9935 m0 *1 118.44,54.6
X$9935 402 39 403 644 645 cell_1rw
* cell instance $9936 m0 *1 119.145,54.6
X$9936 404 39 405 644 645 cell_1rw
* cell instance $9937 m0 *1 119.85,54.6
X$9937 406 39 407 644 645 cell_1rw
* cell instance $9938 m0 *1 120.555,54.6
X$9938 408 39 409 644 645 cell_1rw
* cell instance $9939 m0 *1 121.26,54.6
X$9939 410 39 411 644 645 cell_1rw
* cell instance $9940 m0 *1 121.965,54.6
X$9940 412 39 413 644 645 cell_1rw
* cell instance $9941 m0 *1 122.67,54.6
X$9941 414 39 415 644 645 cell_1rw
* cell instance $9942 m0 *1 123.375,54.6
X$9942 416 39 417 644 645 cell_1rw
* cell instance $9943 m0 *1 124.08,54.6
X$9943 418 39 419 644 645 cell_1rw
* cell instance $9944 m0 *1 124.785,54.6
X$9944 420 39 421 644 645 cell_1rw
* cell instance $9945 m0 *1 125.49,54.6
X$9945 422 39 423 644 645 cell_1rw
* cell instance $9946 m0 *1 126.195,54.6
X$9946 424 39 425 644 645 cell_1rw
* cell instance $9947 m0 *1 126.9,54.6
X$9947 426 39 427 644 645 cell_1rw
* cell instance $9948 m0 *1 127.605,54.6
X$9948 428 39 429 644 645 cell_1rw
* cell instance $9949 m0 *1 128.31,54.6
X$9949 430 39 431 644 645 cell_1rw
* cell instance $9950 m0 *1 129.015,54.6
X$9950 432 39 433 644 645 cell_1rw
* cell instance $9951 m0 *1 129.72,54.6
X$9951 434 39 435 644 645 cell_1rw
* cell instance $9952 m0 *1 130.425,54.6
X$9952 436 39 437 644 645 cell_1rw
* cell instance $9953 m0 *1 131.13,54.6
X$9953 438 39 439 644 645 cell_1rw
* cell instance $9954 m0 *1 131.835,54.6
X$9954 440 39 441 644 645 cell_1rw
* cell instance $9955 m0 *1 132.54,54.6
X$9955 442 39 443 644 645 cell_1rw
* cell instance $9956 m0 *1 133.245,54.6
X$9956 444 39 445 644 645 cell_1rw
* cell instance $9957 m0 *1 133.95,54.6
X$9957 446 39 447 644 645 cell_1rw
* cell instance $9958 m0 *1 134.655,54.6
X$9958 448 39 449 644 645 cell_1rw
* cell instance $9959 m0 *1 135.36,54.6
X$9959 450 39 451 644 645 cell_1rw
* cell instance $9960 m0 *1 136.065,54.6
X$9960 452 39 453 644 645 cell_1rw
* cell instance $9961 m0 *1 136.77,54.6
X$9961 454 39 455 644 645 cell_1rw
* cell instance $9962 m0 *1 137.475,54.6
X$9962 456 39 457 644 645 cell_1rw
* cell instance $9963 m0 *1 138.18,54.6
X$9963 458 39 459 644 645 cell_1rw
* cell instance $9964 m0 *1 138.885,54.6
X$9964 460 39 461 644 645 cell_1rw
* cell instance $9965 m0 *1 139.59,54.6
X$9965 462 39 463 644 645 cell_1rw
* cell instance $9966 m0 *1 140.295,54.6
X$9966 464 39 465 644 645 cell_1rw
* cell instance $9967 m0 *1 141,54.6
X$9967 466 39 467 644 645 cell_1rw
* cell instance $9968 m0 *1 141.705,54.6
X$9968 468 39 469 644 645 cell_1rw
* cell instance $9969 m0 *1 142.41,54.6
X$9969 470 39 471 644 645 cell_1rw
* cell instance $9970 m0 *1 143.115,54.6
X$9970 472 39 473 644 645 cell_1rw
* cell instance $9971 m0 *1 143.82,54.6
X$9971 474 39 475 644 645 cell_1rw
* cell instance $9972 m0 *1 144.525,54.6
X$9972 476 39 477 644 645 cell_1rw
* cell instance $9973 m0 *1 145.23,54.6
X$9973 478 39 479 644 645 cell_1rw
* cell instance $9974 m0 *1 145.935,54.6
X$9974 480 39 481 644 645 cell_1rw
* cell instance $9975 m0 *1 146.64,54.6
X$9975 482 39 483 644 645 cell_1rw
* cell instance $9976 m0 *1 147.345,54.6
X$9976 484 39 485 644 645 cell_1rw
* cell instance $9977 m0 *1 148.05,54.6
X$9977 486 39 487 644 645 cell_1rw
* cell instance $9978 m0 *1 148.755,54.6
X$9978 488 39 489 644 645 cell_1rw
* cell instance $9979 m0 *1 149.46,54.6
X$9979 490 39 491 644 645 cell_1rw
* cell instance $9980 m0 *1 150.165,54.6
X$9980 492 39 493 644 645 cell_1rw
* cell instance $9981 m0 *1 150.87,54.6
X$9981 494 39 495 644 645 cell_1rw
* cell instance $9982 m0 *1 151.575,54.6
X$9982 496 39 497 644 645 cell_1rw
* cell instance $9983 m0 *1 152.28,54.6
X$9983 498 39 499 644 645 cell_1rw
* cell instance $9984 m0 *1 152.985,54.6
X$9984 500 39 501 644 645 cell_1rw
* cell instance $9985 m0 *1 153.69,54.6
X$9985 502 39 503 644 645 cell_1rw
* cell instance $9986 m0 *1 154.395,54.6
X$9986 504 39 505 644 645 cell_1rw
* cell instance $9987 m0 *1 155.1,54.6
X$9987 506 39 507 644 645 cell_1rw
* cell instance $9988 m0 *1 155.805,54.6
X$9988 508 39 509 644 645 cell_1rw
* cell instance $9989 m0 *1 156.51,54.6
X$9989 510 39 511 644 645 cell_1rw
* cell instance $9990 m0 *1 157.215,54.6
X$9990 512 39 513 644 645 cell_1rw
* cell instance $9991 m0 *1 157.92,54.6
X$9991 514 39 515 644 645 cell_1rw
* cell instance $9992 m0 *1 158.625,54.6
X$9992 516 39 517 644 645 cell_1rw
* cell instance $9993 m0 *1 159.33,54.6
X$9993 518 39 519 644 645 cell_1rw
* cell instance $9994 m0 *1 160.035,54.6
X$9994 520 39 521 644 645 cell_1rw
* cell instance $9995 m0 *1 160.74,54.6
X$9995 522 39 523 644 645 cell_1rw
* cell instance $9996 m0 *1 161.445,54.6
X$9996 524 39 525 644 645 cell_1rw
* cell instance $9997 m0 *1 162.15,54.6
X$9997 526 39 527 644 645 cell_1rw
* cell instance $9998 m0 *1 162.855,54.6
X$9998 528 39 529 644 645 cell_1rw
* cell instance $9999 m0 *1 163.56,54.6
X$9999 530 39 531 644 645 cell_1rw
* cell instance $10000 m0 *1 164.265,54.6
X$10000 532 39 533 644 645 cell_1rw
* cell instance $10001 m0 *1 164.97,54.6
X$10001 534 39 535 644 645 cell_1rw
* cell instance $10002 m0 *1 165.675,54.6
X$10002 536 39 537 644 645 cell_1rw
* cell instance $10003 m0 *1 166.38,54.6
X$10003 538 39 539 644 645 cell_1rw
* cell instance $10004 m0 *1 167.085,54.6
X$10004 540 39 541 644 645 cell_1rw
* cell instance $10005 m0 *1 167.79,54.6
X$10005 542 39 543 644 645 cell_1rw
* cell instance $10006 m0 *1 168.495,54.6
X$10006 544 39 545 644 645 cell_1rw
* cell instance $10007 m0 *1 169.2,54.6
X$10007 546 39 547 644 645 cell_1rw
* cell instance $10008 m0 *1 169.905,54.6
X$10008 548 39 549 644 645 cell_1rw
* cell instance $10009 m0 *1 170.61,54.6
X$10009 550 39 551 644 645 cell_1rw
* cell instance $10010 m0 *1 171.315,54.6
X$10010 552 39 553 644 645 cell_1rw
* cell instance $10011 m0 *1 172.02,54.6
X$10011 554 39 555 644 645 cell_1rw
* cell instance $10012 m0 *1 172.725,54.6
X$10012 556 39 557 644 645 cell_1rw
* cell instance $10013 m0 *1 173.43,54.6
X$10013 558 39 559 644 645 cell_1rw
* cell instance $10014 m0 *1 174.135,54.6
X$10014 560 39 561 644 645 cell_1rw
* cell instance $10015 m0 *1 174.84,54.6
X$10015 562 39 563 644 645 cell_1rw
* cell instance $10016 m0 *1 175.545,54.6
X$10016 564 39 565 644 645 cell_1rw
* cell instance $10017 m0 *1 176.25,54.6
X$10017 566 39 567 644 645 cell_1rw
* cell instance $10018 m0 *1 176.955,54.6
X$10018 568 39 569 644 645 cell_1rw
* cell instance $10019 m0 *1 177.66,54.6
X$10019 570 39 571 644 645 cell_1rw
* cell instance $10020 m0 *1 178.365,54.6
X$10020 572 39 573 644 645 cell_1rw
* cell instance $10021 m0 *1 179.07,54.6
X$10021 574 39 575 644 645 cell_1rw
* cell instance $10022 m0 *1 179.775,54.6
X$10022 576 39 577 644 645 cell_1rw
* cell instance $10023 m0 *1 180.48,54.6
X$10023 578 39 579 644 645 cell_1rw
* cell instance $10024 r0 *1 0.705,51.87
X$10024 67 40 68 644 645 cell_1rw
* cell instance $10025 r0 *1 0,51.87
X$10025 65 40 66 644 645 cell_1rw
* cell instance $10026 r0 *1 1.41,51.87
X$10026 69 40 70 644 645 cell_1rw
* cell instance $10027 r0 *1 2.115,51.87
X$10027 71 40 72 644 645 cell_1rw
* cell instance $10028 r0 *1 2.82,51.87
X$10028 73 40 74 644 645 cell_1rw
* cell instance $10029 r0 *1 3.525,51.87
X$10029 75 40 76 644 645 cell_1rw
* cell instance $10030 r0 *1 4.23,51.87
X$10030 77 40 78 644 645 cell_1rw
* cell instance $10031 r0 *1 4.935,51.87
X$10031 79 40 80 644 645 cell_1rw
* cell instance $10032 r0 *1 5.64,51.87
X$10032 81 40 82 644 645 cell_1rw
* cell instance $10033 r0 *1 6.345,51.87
X$10033 83 40 84 644 645 cell_1rw
* cell instance $10034 r0 *1 7.05,51.87
X$10034 85 40 86 644 645 cell_1rw
* cell instance $10035 r0 *1 7.755,51.87
X$10035 87 40 88 644 645 cell_1rw
* cell instance $10036 r0 *1 8.46,51.87
X$10036 89 40 90 644 645 cell_1rw
* cell instance $10037 r0 *1 9.165,51.87
X$10037 91 40 92 644 645 cell_1rw
* cell instance $10038 r0 *1 9.87,51.87
X$10038 93 40 94 644 645 cell_1rw
* cell instance $10039 r0 *1 10.575,51.87
X$10039 95 40 96 644 645 cell_1rw
* cell instance $10040 r0 *1 11.28,51.87
X$10040 97 40 98 644 645 cell_1rw
* cell instance $10041 r0 *1 11.985,51.87
X$10041 99 40 100 644 645 cell_1rw
* cell instance $10042 r0 *1 12.69,51.87
X$10042 101 40 102 644 645 cell_1rw
* cell instance $10043 r0 *1 13.395,51.87
X$10043 103 40 104 644 645 cell_1rw
* cell instance $10044 r0 *1 14.1,51.87
X$10044 105 40 106 644 645 cell_1rw
* cell instance $10045 r0 *1 14.805,51.87
X$10045 107 40 108 644 645 cell_1rw
* cell instance $10046 r0 *1 15.51,51.87
X$10046 109 40 110 644 645 cell_1rw
* cell instance $10047 r0 *1 16.215,51.87
X$10047 111 40 112 644 645 cell_1rw
* cell instance $10048 r0 *1 16.92,51.87
X$10048 113 40 114 644 645 cell_1rw
* cell instance $10049 r0 *1 17.625,51.87
X$10049 115 40 116 644 645 cell_1rw
* cell instance $10050 r0 *1 18.33,51.87
X$10050 117 40 118 644 645 cell_1rw
* cell instance $10051 r0 *1 19.035,51.87
X$10051 119 40 120 644 645 cell_1rw
* cell instance $10052 r0 *1 19.74,51.87
X$10052 121 40 122 644 645 cell_1rw
* cell instance $10053 r0 *1 20.445,51.87
X$10053 123 40 124 644 645 cell_1rw
* cell instance $10054 r0 *1 21.15,51.87
X$10054 125 40 126 644 645 cell_1rw
* cell instance $10055 r0 *1 21.855,51.87
X$10055 127 40 128 644 645 cell_1rw
* cell instance $10056 r0 *1 22.56,51.87
X$10056 129 40 130 644 645 cell_1rw
* cell instance $10057 r0 *1 23.265,51.87
X$10057 131 40 132 644 645 cell_1rw
* cell instance $10058 r0 *1 23.97,51.87
X$10058 133 40 134 644 645 cell_1rw
* cell instance $10059 r0 *1 24.675,51.87
X$10059 135 40 136 644 645 cell_1rw
* cell instance $10060 r0 *1 25.38,51.87
X$10060 137 40 138 644 645 cell_1rw
* cell instance $10061 r0 *1 26.085,51.87
X$10061 139 40 140 644 645 cell_1rw
* cell instance $10062 r0 *1 26.79,51.87
X$10062 141 40 142 644 645 cell_1rw
* cell instance $10063 r0 *1 27.495,51.87
X$10063 143 40 144 644 645 cell_1rw
* cell instance $10064 r0 *1 28.2,51.87
X$10064 145 40 146 644 645 cell_1rw
* cell instance $10065 r0 *1 28.905,51.87
X$10065 147 40 148 644 645 cell_1rw
* cell instance $10066 r0 *1 29.61,51.87
X$10066 149 40 150 644 645 cell_1rw
* cell instance $10067 r0 *1 30.315,51.87
X$10067 151 40 152 644 645 cell_1rw
* cell instance $10068 r0 *1 31.02,51.87
X$10068 153 40 154 644 645 cell_1rw
* cell instance $10069 r0 *1 31.725,51.87
X$10069 155 40 156 644 645 cell_1rw
* cell instance $10070 r0 *1 32.43,51.87
X$10070 157 40 158 644 645 cell_1rw
* cell instance $10071 r0 *1 33.135,51.87
X$10071 159 40 160 644 645 cell_1rw
* cell instance $10072 r0 *1 33.84,51.87
X$10072 161 40 162 644 645 cell_1rw
* cell instance $10073 r0 *1 34.545,51.87
X$10073 163 40 164 644 645 cell_1rw
* cell instance $10074 r0 *1 35.25,51.87
X$10074 165 40 166 644 645 cell_1rw
* cell instance $10075 r0 *1 35.955,51.87
X$10075 167 40 168 644 645 cell_1rw
* cell instance $10076 r0 *1 36.66,51.87
X$10076 169 40 170 644 645 cell_1rw
* cell instance $10077 r0 *1 37.365,51.87
X$10077 171 40 172 644 645 cell_1rw
* cell instance $10078 r0 *1 38.07,51.87
X$10078 173 40 174 644 645 cell_1rw
* cell instance $10079 r0 *1 38.775,51.87
X$10079 175 40 176 644 645 cell_1rw
* cell instance $10080 r0 *1 39.48,51.87
X$10080 177 40 178 644 645 cell_1rw
* cell instance $10081 r0 *1 40.185,51.87
X$10081 179 40 180 644 645 cell_1rw
* cell instance $10082 r0 *1 40.89,51.87
X$10082 181 40 182 644 645 cell_1rw
* cell instance $10083 r0 *1 41.595,51.87
X$10083 183 40 184 644 645 cell_1rw
* cell instance $10084 r0 *1 42.3,51.87
X$10084 185 40 186 644 645 cell_1rw
* cell instance $10085 r0 *1 43.005,51.87
X$10085 187 40 188 644 645 cell_1rw
* cell instance $10086 r0 *1 43.71,51.87
X$10086 189 40 190 644 645 cell_1rw
* cell instance $10087 r0 *1 44.415,51.87
X$10087 191 40 192 644 645 cell_1rw
* cell instance $10088 r0 *1 45.12,51.87
X$10088 193 40 194 644 645 cell_1rw
* cell instance $10089 r0 *1 45.825,51.87
X$10089 195 40 196 644 645 cell_1rw
* cell instance $10090 r0 *1 46.53,51.87
X$10090 197 40 198 644 645 cell_1rw
* cell instance $10091 r0 *1 47.235,51.87
X$10091 199 40 200 644 645 cell_1rw
* cell instance $10092 r0 *1 47.94,51.87
X$10092 201 40 202 644 645 cell_1rw
* cell instance $10093 r0 *1 48.645,51.87
X$10093 203 40 204 644 645 cell_1rw
* cell instance $10094 r0 *1 49.35,51.87
X$10094 205 40 206 644 645 cell_1rw
* cell instance $10095 r0 *1 50.055,51.87
X$10095 207 40 208 644 645 cell_1rw
* cell instance $10096 r0 *1 50.76,51.87
X$10096 209 40 210 644 645 cell_1rw
* cell instance $10097 r0 *1 51.465,51.87
X$10097 211 40 212 644 645 cell_1rw
* cell instance $10098 r0 *1 52.17,51.87
X$10098 213 40 214 644 645 cell_1rw
* cell instance $10099 r0 *1 52.875,51.87
X$10099 215 40 216 644 645 cell_1rw
* cell instance $10100 r0 *1 53.58,51.87
X$10100 217 40 218 644 645 cell_1rw
* cell instance $10101 r0 *1 54.285,51.87
X$10101 219 40 220 644 645 cell_1rw
* cell instance $10102 r0 *1 54.99,51.87
X$10102 221 40 222 644 645 cell_1rw
* cell instance $10103 r0 *1 55.695,51.87
X$10103 223 40 224 644 645 cell_1rw
* cell instance $10104 r0 *1 56.4,51.87
X$10104 225 40 226 644 645 cell_1rw
* cell instance $10105 r0 *1 57.105,51.87
X$10105 227 40 228 644 645 cell_1rw
* cell instance $10106 r0 *1 57.81,51.87
X$10106 229 40 230 644 645 cell_1rw
* cell instance $10107 r0 *1 58.515,51.87
X$10107 231 40 232 644 645 cell_1rw
* cell instance $10108 r0 *1 59.22,51.87
X$10108 233 40 234 644 645 cell_1rw
* cell instance $10109 r0 *1 59.925,51.87
X$10109 235 40 236 644 645 cell_1rw
* cell instance $10110 r0 *1 60.63,51.87
X$10110 237 40 238 644 645 cell_1rw
* cell instance $10111 r0 *1 61.335,51.87
X$10111 239 40 240 644 645 cell_1rw
* cell instance $10112 r0 *1 62.04,51.87
X$10112 241 40 242 644 645 cell_1rw
* cell instance $10113 r0 *1 62.745,51.87
X$10113 243 40 244 644 645 cell_1rw
* cell instance $10114 r0 *1 63.45,51.87
X$10114 245 40 246 644 645 cell_1rw
* cell instance $10115 r0 *1 64.155,51.87
X$10115 247 40 248 644 645 cell_1rw
* cell instance $10116 r0 *1 64.86,51.87
X$10116 249 40 250 644 645 cell_1rw
* cell instance $10117 r0 *1 65.565,51.87
X$10117 251 40 252 644 645 cell_1rw
* cell instance $10118 r0 *1 66.27,51.87
X$10118 253 40 254 644 645 cell_1rw
* cell instance $10119 r0 *1 66.975,51.87
X$10119 255 40 256 644 645 cell_1rw
* cell instance $10120 r0 *1 67.68,51.87
X$10120 257 40 258 644 645 cell_1rw
* cell instance $10121 r0 *1 68.385,51.87
X$10121 259 40 260 644 645 cell_1rw
* cell instance $10122 r0 *1 69.09,51.87
X$10122 261 40 262 644 645 cell_1rw
* cell instance $10123 r0 *1 69.795,51.87
X$10123 263 40 264 644 645 cell_1rw
* cell instance $10124 r0 *1 70.5,51.87
X$10124 265 40 266 644 645 cell_1rw
* cell instance $10125 r0 *1 71.205,51.87
X$10125 267 40 268 644 645 cell_1rw
* cell instance $10126 r0 *1 71.91,51.87
X$10126 269 40 270 644 645 cell_1rw
* cell instance $10127 r0 *1 72.615,51.87
X$10127 271 40 272 644 645 cell_1rw
* cell instance $10128 r0 *1 73.32,51.87
X$10128 273 40 274 644 645 cell_1rw
* cell instance $10129 r0 *1 74.025,51.87
X$10129 275 40 276 644 645 cell_1rw
* cell instance $10130 r0 *1 74.73,51.87
X$10130 277 40 278 644 645 cell_1rw
* cell instance $10131 r0 *1 75.435,51.87
X$10131 279 40 280 644 645 cell_1rw
* cell instance $10132 r0 *1 76.14,51.87
X$10132 281 40 282 644 645 cell_1rw
* cell instance $10133 r0 *1 76.845,51.87
X$10133 283 40 284 644 645 cell_1rw
* cell instance $10134 r0 *1 77.55,51.87
X$10134 285 40 286 644 645 cell_1rw
* cell instance $10135 r0 *1 78.255,51.87
X$10135 287 40 288 644 645 cell_1rw
* cell instance $10136 r0 *1 78.96,51.87
X$10136 289 40 290 644 645 cell_1rw
* cell instance $10137 r0 *1 79.665,51.87
X$10137 291 40 292 644 645 cell_1rw
* cell instance $10138 r0 *1 80.37,51.87
X$10138 293 40 294 644 645 cell_1rw
* cell instance $10139 r0 *1 81.075,51.87
X$10139 295 40 296 644 645 cell_1rw
* cell instance $10140 r0 *1 81.78,51.87
X$10140 297 40 298 644 645 cell_1rw
* cell instance $10141 r0 *1 82.485,51.87
X$10141 299 40 300 644 645 cell_1rw
* cell instance $10142 r0 *1 83.19,51.87
X$10142 301 40 302 644 645 cell_1rw
* cell instance $10143 r0 *1 83.895,51.87
X$10143 303 40 304 644 645 cell_1rw
* cell instance $10144 r0 *1 84.6,51.87
X$10144 305 40 306 644 645 cell_1rw
* cell instance $10145 r0 *1 85.305,51.87
X$10145 307 40 308 644 645 cell_1rw
* cell instance $10146 r0 *1 86.01,51.87
X$10146 309 40 310 644 645 cell_1rw
* cell instance $10147 r0 *1 86.715,51.87
X$10147 311 40 312 644 645 cell_1rw
* cell instance $10148 r0 *1 87.42,51.87
X$10148 313 40 314 644 645 cell_1rw
* cell instance $10149 r0 *1 88.125,51.87
X$10149 315 40 316 644 645 cell_1rw
* cell instance $10150 r0 *1 88.83,51.87
X$10150 317 40 318 644 645 cell_1rw
* cell instance $10151 r0 *1 89.535,51.87
X$10151 319 40 320 644 645 cell_1rw
* cell instance $10152 r0 *1 90.24,51.87
X$10152 321 40 323 644 645 cell_1rw
* cell instance $10153 r0 *1 90.945,51.87
X$10153 324 40 325 644 645 cell_1rw
* cell instance $10154 r0 *1 91.65,51.87
X$10154 326 40 327 644 645 cell_1rw
* cell instance $10155 r0 *1 92.355,51.87
X$10155 328 40 329 644 645 cell_1rw
* cell instance $10156 r0 *1 93.06,51.87
X$10156 330 40 331 644 645 cell_1rw
* cell instance $10157 r0 *1 93.765,51.87
X$10157 332 40 333 644 645 cell_1rw
* cell instance $10158 r0 *1 94.47,51.87
X$10158 334 40 335 644 645 cell_1rw
* cell instance $10159 r0 *1 95.175,51.87
X$10159 336 40 337 644 645 cell_1rw
* cell instance $10160 r0 *1 95.88,51.87
X$10160 338 40 339 644 645 cell_1rw
* cell instance $10161 r0 *1 96.585,51.87
X$10161 340 40 341 644 645 cell_1rw
* cell instance $10162 r0 *1 97.29,51.87
X$10162 342 40 343 644 645 cell_1rw
* cell instance $10163 r0 *1 97.995,51.87
X$10163 344 40 345 644 645 cell_1rw
* cell instance $10164 r0 *1 98.7,51.87
X$10164 346 40 347 644 645 cell_1rw
* cell instance $10165 r0 *1 99.405,51.87
X$10165 348 40 349 644 645 cell_1rw
* cell instance $10166 r0 *1 100.11,51.87
X$10166 350 40 351 644 645 cell_1rw
* cell instance $10167 r0 *1 100.815,51.87
X$10167 352 40 353 644 645 cell_1rw
* cell instance $10168 r0 *1 101.52,51.87
X$10168 354 40 355 644 645 cell_1rw
* cell instance $10169 r0 *1 102.225,51.87
X$10169 356 40 357 644 645 cell_1rw
* cell instance $10170 r0 *1 102.93,51.87
X$10170 358 40 359 644 645 cell_1rw
* cell instance $10171 r0 *1 103.635,51.87
X$10171 360 40 361 644 645 cell_1rw
* cell instance $10172 r0 *1 104.34,51.87
X$10172 362 40 363 644 645 cell_1rw
* cell instance $10173 r0 *1 105.045,51.87
X$10173 364 40 365 644 645 cell_1rw
* cell instance $10174 r0 *1 105.75,51.87
X$10174 366 40 367 644 645 cell_1rw
* cell instance $10175 r0 *1 106.455,51.87
X$10175 368 40 369 644 645 cell_1rw
* cell instance $10176 r0 *1 107.16,51.87
X$10176 370 40 371 644 645 cell_1rw
* cell instance $10177 r0 *1 107.865,51.87
X$10177 372 40 373 644 645 cell_1rw
* cell instance $10178 r0 *1 108.57,51.87
X$10178 374 40 375 644 645 cell_1rw
* cell instance $10179 r0 *1 109.275,51.87
X$10179 376 40 377 644 645 cell_1rw
* cell instance $10180 r0 *1 109.98,51.87
X$10180 378 40 379 644 645 cell_1rw
* cell instance $10181 r0 *1 110.685,51.87
X$10181 380 40 381 644 645 cell_1rw
* cell instance $10182 r0 *1 111.39,51.87
X$10182 382 40 383 644 645 cell_1rw
* cell instance $10183 r0 *1 112.095,51.87
X$10183 384 40 385 644 645 cell_1rw
* cell instance $10184 r0 *1 112.8,51.87
X$10184 386 40 387 644 645 cell_1rw
* cell instance $10185 r0 *1 113.505,51.87
X$10185 388 40 389 644 645 cell_1rw
* cell instance $10186 r0 *1 114.21,51.87
X$10186 390 40 391 644 645 cell_1rw
* cell instance $10187 r0 *1 114.915,51.87
X$10187 392 40 393 644 645 cell_1rw
* cell instance $10188 r0 *1 115.62,51.87
X$10188 394 40 395 644 645 cell_1rw
* cell instance $10189 r0 *1 116.325,51.87
X$10189 396 40 397 644 645 cell_1rw
* cell instance $10190 r0 *1 117.03,51.87
X$10190 398 40 399 644 645 cell_1rw
* cell instance $10191 r0 *1 117.735,51.87
X$10191 400 40 401 644 645 cell_1rw
* cell instance $10192 r0 *1 118.44,51.87
X$10192 402 40 403 644 645 cell_1rw
* cell instance $10193 r0 *1 119.145,51.87
X$10193 404 40 405 644 645 cell_1rw
* cell instance $10194 r0 *1 119.85,51.87
X$10194 406 40 407 644 645 cell_1rw
* cell instance $10195 r0 *1 120.555,51.87
X$10195 408 40 409 644 645 cell_1rw
* cell instance $10196 r0 *1 121.26,51.87
X$10196 410 40 411 644 645 cell_1rw
* cell instance $10197 r0 *1 121.965,51.87
X$10197 412 40 413 644 645 cell_1rw
* cell instance $10198 r0 *1 122.67,51.87
X$10198 414 40 415 644 645 cell_1rw
* cell instance $10199 r0 *1 123.375,51.87
X$10199 416 40 417 644 645 cell_1rw
* cell instance $10200 r0 *1 124.08,51.87
X$10200 418 40 419 644 645 cell_1rw
* cell instance $10201 r0 *1 124.785,51.87
X$10201 420 40 421 644 645 cell_1rw
* cell instance $10202 r0 *1 125.49,51.87
X$10202 422 40 423 644 645 cell_1rw
* cell instance $10203 r0 *1 126.195,51.87
X$10203 424 40 425 644 645 cell_1rw
* cell instance $10204 r0 *1 126.9,51.87
X$10204 426 40 427 644 645 cell_1rw
* cell instance $10205 r0 *1 127.605,51.87
X$10205 428 40 429 644 645 cell_1rw
* cell instance $10206 r0 *1 128.31,51.87
X$10206 430 40 431 644 645 cell_1rw
* cell instance $10207 r0 *1 129.015,51.87
X$10207 432 40 433 644 645 cell_1rw
* cell instance $10208 r0 *1 129.72,51.87
X$10208 434 40 435 644 645 cell_1rw
* cell instance $10209 r0 *1 130.425,51.87
X$10209 436 40 437 644 645 cell_1rw
* cell instance $10210 r0 *1 131.13,51.87
X$10210 438 40 439 644 645 cell_1rw
* cell instance $10211 r0 *1 131.835,51.87
X$10211 440 40 441 644 645 cell_1rw
* cell instance $10212 r0 *1 132.54,51.87
X$10212 442 40 443 644 645 cell_1rw
* cell instance $10213 r0 *1 133.245,51.87
X$10213 444 40 445 644 645 cell_1rw
* cell instance $10214 r0 *1 133.95,51.87
X$10214 446 40 447 644 645 cell_1rw
* cell instance $10215 r0 *1 134.655,51.87
X$10215 448 40 449 644 645 cell_1rw
* cell instance $10216 r0 *1 135.36,51.87
X$10216 450 40 451 644 645 cell_1rw
* cell instance $10217 r0 *1 136.065,51.87
X$10217 452 40 453 644 645 cell_1rw
* cell instance $10218 r0 *1 136.77,51.87
X$10218 454 40 455 644 645 cell_1rw
* cell instance $10219 r0 *1 137.475,51.87
X$10219 456 40 457 644 645 cell_1rw
* cell instance $10220 r0 *1 138.18,51.87
X$10220 458 40 459 644 645 cell_1rw
* cell instance $10221 r0 *1 138.885,51.87
X$10221 460 40 461 644 645 cell_1rw
* cell instance $10222 r0 *1 139.59,51.87
X$10222 462 40 463 644 645 cell_1rw
* cell instance $10223 r0 *1 140.295,51.87
X$10223 464 40 465 644 645 cell_1rw
* cell instance $10224 r0 *1 141,51.87
X$10224 466 40 467 644 645 cell_1rw
* cell instance $10225 r0 *1 141.705,51.87
X$10225 468 40 469 644 645 cell_1rw
* cell instance $10226 r0 *1 142.41,51.87
X$10226 470 40 471 644 645 cell_1rw
* cell instance $10227 r0 *1 143.115,51.87
X$10227 472 40 473 644 645 cell_1rw
* cell instance $10228 r0 *1 143.82,51.87
X$10228 474 40 475 644 645 cell_1rw
* cell instance $10229 r0 *1 144.525,51.87
X$10229 476 40 477 644 645 cell_1rw
* cell instance $10230 r0 *1 145.23,51.87
X$10230 478 40 479 644 645 cell_1rw
* cell instance $10231 r0 *1 145.935,51.87
X$10231 480 40 481 644 645 cell_1rw
* cell instance $10232 r0 *1 146.64,51.87
X$10232 482 40 483 644 645 cell_1rw
* cell instance $10233 r0 *1 147.345,51.87
X$10233 484 40 485 644 645 cell_1rw
* cell instance $10234 r0 *1 148.05,51.87
X$10234 486 40 487 644 645 cell_1rw
* cell instance $10235 r0 *1 148.755,51.87
X$10235 488 40 489 644 645 cell_1rw
* cell instance $10236 r0 *1 149.46,51.87
X$10236 490 40 491 644 645 cell_1rw
* cell instance $10237 r0 *1 150.165,51.87
X$10237 492 40 493 644 645 cell_1rw
* cell instance $10238 r0 *1 150.87,51.87
X$10238 494 40 495 644 645 cell_1rw
* cell instance $10239 r0 *1 151.575,51.87
X$10239 496 40 497 644 645 cell_1rw
* cell instance $10240 r0 *1 152.28,51.87
X$10240 498 40 499 644 645 cell_1rw
* cell instance $10241 r0 *1 152.985,51.87
X$10241 500 40 501 644 645 cell_1rw
* cell instance $10242 r0 *1 153.69,51.87
X$10242 502 40 503 644 645 cell_1rw
* cell instance $10243 r0 *1 154.395,51.87
X$10243 504 40 505 644 645 cell_1rw
* cell instance $10244 r0 *1 155.1,51.87
X$10244 506 40 507 644 645 cell_1rw
* cell instance $10245 r0 *1 155.805,51.87
X$10245 508 40 509 644 645 cell_1rw
* cell instance $10246 r0 *1 156.51,51.87
X$10246 510 40 511 644 645 cell_1rw
* cell instance $10247 r0 *1 157.215,51.87
X$10247 512 40 513 644 645 cell_1rw
* cell instance $10248 r0 *1 157.92,51.87
X$10248 514 40 515 644 645 cell_1rw
* cell instance $10249 r0 *1 158.625,51.87
X$10249 516 40 517 644 645 cell_1rw
* cell instance $10250 r0 *1 159.33,51.87
X$10250 518 40 519 644 645 cell_1rw
* cell instance $10251 r0 *1 160.035,51.87
X$10251 520 40 521 644 645 cell_1rw
* cell instance $10252 r0 *1 160.74,51.87
X$10252 522 40 523 644 645 cell_1rw
* cell instance $10253 r0 *1 161.445,51.87
X$10253 524 40 525 644 645 cell_1rw
* cell instance $10254 r0 *1 162.15,51.87
X$10254 526 40 527 644 645 cell_1rw
* cell instance $10255 r0 *1 162.855,51.87
X$10255 528 40 529 644 645 cell_1rw
* cell instance $10256 r0 *1 163.56,51.87
X$10256 530 40 531 644 645 cell_1rw
* cell instance $10257 r0 *1 164.265,51.87
X$10257 532 40 533 644 645 cell_1rw
* cell instance $10258 r0 *1 164.97,51.87
X$10258 534 40 535 644 645 cell_1rw
* cell instance $10259 r0 *1 165.675,51.87
X$10259 536 40 537 644 645 cell_1rw
* cell instance $10260 r0 *1 166.38,51.87
X$10260 538 40 539 644 645 cell_1rw
* cell instance $10261 r0 *1 167.085,51.87
X$10261 540 40 541 644 645 cell_1rw
* cell instance $10262 r0 *1 167.79,51.87
X$10262 542 40 543 644 645 cell_1rw
* cell instance $10263 r0 *1 168.495,51.87
X$10263 544 40 545 644 645 cell_1rw
* cell instance $10264 r0 *1 169.2,51.87
X$10264 546 40 547 644 645 cell_1rw
* cell instance $10265 r0 *1 169.905,51.87
X$10265 548 40 549 644 645 cell_1rw
* cell instance $10266 r0 *1 170.61,51.87
X$10266 550 40 551 644 645 cell_1rw
* cell instance $10267 r0 *1 171.315,51.87
X$10267 552 40 553 644 645 cell_1rw
* cell instance $10268 r0 *1 172.02,51.87
X$10268 554 40 555 644 645 cell_1rw
* cell instance $10269 r0 *1 172.725,51.87
X$10269 556 40 557 644 645 cell_1rw
* cell instance $10270 r0 *1 173.43,51.87
X$10270 558 40 559 644 645 cell_1rw
* cell instance $10271 r0 *1 174.135,51.87
X$10271 560 40 561 644 645 cell_1rw
* cell instance $10272 r0 *1 174.84,51.87
X$10272 562 40 563 644 645 cell_1rw
* cell instance $10273 r0 *1 175.545,51.87
X$10273 564 40 565 644 645 cell_1rw
* cell instance $10274 r0 *1 176.25,51.87
X$10274 566 40 567 644 645 cell_1rw
* cell instance $10275 r0 *1 176.955,51.87
X$10275 568 40 569 644 645 cell_1rw
* cell instance $10276 r0 *1 177.66,51.87
X$10276 570 40 571 644 645 cell_1rw
* cell instance $10277 r0 *1 178.365,51.87
X$10277 572 40 573 644 645 cell_1rw
* cell instance $10278 r0 *1 179.07,51.87
X$10278 574 40 575 644 645 cell_1rw
* cell instance $10279 r0 *1 179.775,51.87
X$10279 576 40 577 644 645 cell_1rw
* cell instance $10280 r0 *1 180.48,51.87
X$10280 578 40 579 644 645 cell_1rw
* cell instance $10281 m0 *1 0.705,57.33
X$10281 67 41 68 644 645 cell_1rw
* cell instance $10282 m0 *1 0,57.33
X$10282 65 41 66 644 645 cell_1rw
* cell instance $10283 m0 *1 1.41,57.33
X$10283 69 41 70 644 645 cell_1rw
* cell instance $10284 m0 *1 2.115,57.33
X$10284 71 41 72 644 645 cell_1rw
* cell instance $10285 m0 *1 2.82,57.33
X$10285 73 41 74 644 645 cell_1rw
* cell instance $10286 m0 *1 3.525,57.33
X$10286 75 41 76 644 645 cell_1rw
* cell instance $10287 m0 *1 4.23,57.33
X$10287 77 41 78 644 645 cell_1rw
* cell instance $10288 m0 *1 4.935,57.33
X$10288 79 41 80 644 645 cell_1rw
* cell instance $10289 m0 *1 5.64,57.33
X$10289 81 41 82 644 645 cell_1rw
* cell instance $10290 m0 *1 6.345,57.33
X$10290 83 41 84 644 645 cell_1rw
* cell instance $10291 m0 *1 7.05,57.33
X$10291 85 41 86 644 645 cell_1rw
* cell instance $10292 m0 *1 7.755,57.33
X$10292 87 41 88 644 645 cell_1rw
* cell instance $10293 m0 *1 8.46,57.33
X$10293 89 41 90 644 645 cell_1rw
* cell instance $10294 m0 *1 9.165,57.33
X$10294 91 41 92 644 645 cell_1rw
* cell instance $10295 m0 *1 9.87,57.33
X$10295 93 41 94 644 645 cell_1rw
* cell instance $10296 m0 *1 10.575,57.33
X$10296 95 41 96 644 645 cell_1rw
* cell instance $10297 m0 *1 11.28,57.33
X$10297 97 41 98 644 645 cell_1rw
* cell instance $10298 m0 *1 11.985,57.33
X$10298 99 41 100 644 645 cell_1rw
* cell instance $10299 m0 *1 12.69,57.33
X$10299 101 41 102 644 645 cell_1rw
* cell instance $10300 m0 *1 13.395,57.33
X$10300 103 41 104 644 645 cell_1rw
* cell instance $10301 m0 *1 14.1,57.33
X$10301 105 41 106 644 645 cell_1rw
* cell instance $10302 m0 *1 14.805,57.33
X$10302 107 41 108 644 645 cell_1rw
* cell instance $10303 m0 *1 15.51,57.33
X$10303 109 41 110 644 645 cell_1rw
* cell instance $10304 m0 *1 16.215,57.33
X$10304 111 41 112 644 645 cell_1rw
* cell instance $10305 m0 *1 16.92,57.33
X$10305 113 41 114 644 645 cell_1rw
* cell instance $10306 m0 *1 17.625,57.33
X$10306 115 41 116 644 645 cell_1rw
* cell instance $10307 m0 *1 18.33,57.33
X$10307 117 41 118 644 645 cell_1rw
* cell instance $10308 m0 *1 19.035,57.33
X$10308 119 41 120 644 645 cell_1rw
* cell instance $10309 m0 *1 19.74,57.33
X$10309 121 41 122 644 645 cell_1rw
* cell instance $10310 m0 *1 20.445,57.33
X$10310 123 41 124 644 645 cell_1rw
* cell instance $10311 m0 *1 21.15,57.33
X$10311 125 41 126 644 645 cell_1rw
* cell instance $10312 m0 *1 21.855,57.33
X$10312 127 41 128 644 645 cell_1rw
* cell instance $10313 m0 *1 22.56,57.33
X$10313 129 41 130 644 645 cell_1rw
* cell instance $10314 m0 *1 23.265,57.33
X$10314 131 41 132 644 645 cell_1rw
* cell instance $10315 m0 *1 23.97,57.33
X$10315 133 41 134 644 645 cell_1rw
* cell instance $10316 m0 *1 24.675,57.33
X$10316 135 41 136 644 645 cell_1rw
* cell instance $10317 m0 *1 25.38,57.33
X$10317 137 41 138 644 645 cell_1rw
* cell instance $10318 m0 *1 26.085,57.33
X$10318 139 41 140 644 645 cell_1rw
* cell instance $10319 m0 *1 26.79,57.33
X$10319 141 41 142 644 645 cell_1rw
* cell instance $10320 m0 *1 27.495,57.33
X$10320 143 41 144 644 645 cell_1rw
* cell instance $10321 m0 *1 28.2,57.33
X$10321 145 41 146 644 645 cell_1rw
* cell instance $10322 m0 *1 28.905,57.33
X$10322 147 41 148 644 645 cell_1rw
* cell instance $10323 m0 *1 29.61,57.33
X$10323 149 41 150 644 645 cell_1rw
* cell instance $10324 m0 *1 30.315,57.33
X$10324 151 41 152 644 645 cell_1rw
* cell instance $10325 m0 *1 31.02,57.33
X$10325 153 41 154 644 645 cell_1rw
* cell instance $10326 m0 *1 31.725,57.33
X$10326 155 41 156 644 645 cell_1rw
* cell instance $10327 m0 *1 32.43,57.33
X$10327 157 41 158 644 645 cell_1rw
* cell instance $10328 m0 *1 33.135,57.33
X$10328 159 41 160 644 645 cell_1rw
* cell instance $10329 m0 *1 33.84,57.33
X$10329 161 41 162 644 645 cell_1rw
* cell instance $10330 m0 *1 34.545,57.33
X$10330 163 41 164 644 645 cell_1rw
* cell instance $10331 m0 *1 35.25,57.33
X$10331 165 41 166 644 645 cell_1rw
* cell instance $10332 m0 *1 35.955,57.33
X$10332 167 41 168 644 645 cell_1rw
* cell instance $10333 m0 *1 36.66,57.33
X$10333 169 41 170 644 645 cell_1rw
* cell instance $10334 m0 *1 37.365,57.33
X$10334 171 41 172 644 645 cell_1rw
* cell instance $10335 m0 *1 38.07,57.33
X$10335 173 41 174 644 645 cell_1rw
* cell instance $10336 m0 *1 38.775,57.33
X$10336 175 41 176 644 645 cell_1rw
* cell instance $10337 m0 *1 39.48,57.33
X$10337 177 41 178 644 645 cell_1rw
* cell instance $10338 m0 *1 40.185,57.33
X$10338 179 41 180 644 645 cell_1rw
* cell instance $10339 m0 *1 40.89,57.33
X$10339 181 41 182 644 645 cell_1rw
* cell instance $10340 m0 *1 41.595,57.33
X$10340 183 41 184 644 645 cell_1rw
* cell instance $10341 m0 *1 42.3,57.33
X$10341 185 41 186 644 645 cell_1rw
* cell instance $10342 m0 *1 43.005,57.33
X$10342 187 41 188 644 645 cell_1rw
* cell instance $10343 m0 *1 43.71,57.33
X$10343 189 41 190 644 645 cell_1rw
* cell instance $10344 m0 *1 44.415,57.33
X$10344 191 41 192 644 645 cell_1rw
* cell instance $10345 m0 *1 45.12,57.33
X$10345 193 41 194 644 645 cell_1rw
* cell instance $10346 m0 *1 45.825,57.33
X$10346 195 41 196 644 645 cell_1rw
* cell instance $10347 m0 *1 46.53,57.33
X$10347 197 41 198 644 645 cell_1rw
* cell instance $10348 m0 *1 47.235,57.33
X$10348 199 41 200 644 645 cell_1rw
* cell instance $10349 m0 *1 47.94,57.33
X$10349 201 41 202 644 645 cell_1rw
* cell instance $10350 m0 *1 48.645,57.33
X$10350 203 41 204 644 645 cell_1rw
* cell instance $10351 m0 *1 49.35,57.33
X$10351 205 41 206 644 645 cell_1rw
* cell instance $10352 m0 *1 50.055,57.33
X$10352 207 41 208 644 645 cell_1rw
* cell instance $10353 m0 *1 50.76,57.33
X$10353 209 41 210 644 645 cell_1rw
* cell instance $10354 m0 *1 51.465,57.33
X$10354 211 41 212 644 645 cell_1rw
* cell instance $10355 m0 *1 52.17,57.33
X$10355 213 41 214 644 645 cell_1rw
* cell instance $10356 m0 *1 52.875,57.33
X$10356 215 41 216 644 645 cell_1rw
* cell instance $10357 m0 *1 53.58,57.33
X$10357 217 41 218 644 645 cell_1rw
* cell instance $10358 m0 *1 54.285,57.33
X$10358 219 41 220 644 645 cell_1rw
* cell instance $10359 m0 *1 54.99,57.33
X$10359 221 41 222 644 645 cell_1rw
* cell instance $10360 m0 *1 55.695,57.33
X$10360 223 41 224 644 645 cell_1rw
* cell instance $10361 m0 *1 56.4,57.33
X$10361 225 41 226 644 645 cell_1rw
* cell instance $10362 m0 *1 57.105,57.33
X$10362 227 41 228 644 645 cell_1rw
* cell instance $10363 m0 *1 57.81,57.33
X$10363 229 41 230 644 645 cell_1rw
* cell instance $10364 m0 *1 58.515,57.33
X$10364 231 41 232 644 645 cell_1rw
* cell instance $10365 m0 *1 59.22,57.33
X$10365 233 41 234 644 645 cell_1rw
* cell instance $10366 m0 *1 59.925,57.33
X$10366 235 41 236 644 645 cell_1rw
* cell instance $10367 m0 *1 60.63,57.33
X$10367 237 41 238 644 645 cell_1rw
* cell instance $10368 m0 *1 61.335,57.33
X$10368 239 41 240 644 645 cell_1rw
* cell instance $10369 m0 *1 62.04,57.33
X$10369 241 41 242 644 645 cell_1rw
* cell instance $10370 m0 *1 62.745,57.33
X$10370 243 41 244 644 645 cell_1rw
* cell instance $10371 m0 *1 63.45,57.33
X$10371 245 41 246 644 645 cell_1rw
* cell instance $10372 m0 *1 64.155,57.33
X$10372 247 41 248 644 645 cell_1rw
* cell instance $10373 m0 *1 64.86,57.33
X$10373 249 41 250 644 645 cell_1rw
* cell instance $10374 m0 *1 65.565,57.33
X$10374 251 41 252 644 645 cell_1rw
* cell instance $10375 m0 *1 66.27,57.33
X$10375 253 41 254 644 645 cell_1rw
* cell instance $10376 m0 *1 66.975,57.33
X$10376 255 41 256 644 645 cell_1rw
* cell instance $10377 m0 *1 67.68,57.33
X$10377 257 41 258 644 645 cell_1rw
* cell instance $10378 m0 *1 68.385,57.33
X$10378 259 41 260 644 645 cell_1rw
* cell instance $10379 m0 *1 69.09,57.33
X$10379 261 41 262 644 645 cell_1rw
* cell instance $10380 m0 *1 69.795,57.33
X$10380 263 41 264 644 645 cell_1rw
* cell instance $10381 m0 *1 70.5,57.33
X$10381 265 41 266 644 645 cell_1rw
* cell instance $10382 m0 *1 71.205,57.33
X$10382 267 41 268 644 645 cell_1rw
* cell instance $10383 m0 *1 71.91,57.33
X$10383 269 41 270 644 645 cell_1rw
* cell instance $10384 m0 *1 72.615,57.33
X$10384 271 41 272 644 645 cell_1rw
* cell instance $10385 m0 *1 73.32,57.33
X$10385 273 41 274 644 645 cell_1rw
* cell instance $10386 m0 *1 74.025,57.33
X$10386 275 41 276 644 645 cell_1rw
* cell instance $10387 m0 *1 74.73,57.33
X$10387 277 41 278 644 645 cell_1rw
* cell instance $10388 m0 *1 75.435,57.33
X$10388 279 41 280 644 645 cell_1rw
* cell instance $10389 m0 *1 76.14,57.33
X$10389 281 41 282 644 645 cell_1rw
* cell instance $10390 m0 *1 76.845,57.33
X$10390 283 41 284 644 645 cell_1rw
* cell instance $10391 m0 *1 77.55,57.33
X$10391 285 41 286 644 645 cell_1rw
* cell instance $10392 m0 *1 78.255,57.33
X$10392 287 41 288 644 645 cell_1rw
* cell instance $10393 m0 *1 78.96,57.33
X$10393 289 41 290 644 645 cell_1rw
* cell instance $10394 m0 *1 79.665,57.33
X$10394 291 41 292 644 645 cell_1rw
* cell instance $10395 m0 *1 80.37,57.33
X$10395 293 41 294 644 645 cell_1rw
* cell instance $10396 m0 *1 81.075,57.33
X$10396 295 41 296 644 645 cell_1rw
* cell instance $10397 m0 *1 81.78,57.33
X$10397 297 41 298 644 645 cell_1rw
* cell instance $10398 m0 *1 82.485,57.33
X$10398 299 41 300 644 645 cell_1rw
* cell instance $10399 m0 *1 83.19,57.33
X$10399 301 41 302 644 645 cell_1rw
* cell instance $10400 m0 *1 83.895,57.33
X$10400 303 41 304 644 645 cell_1rw
* cell instance $10401 m0 *1 84.6,57.33
X$10401 305 41 306 644 645 cell_1rw
* cell instance $10402 m0 *1 85.305,57.33
X$10402 307 41 308 644 645 cell_1rw
* cell instance $10403 m0 *1 86.01,57.33
X$10403 309 41 310 644 645 cell_1rw
* cell instance $10404 m0 *1 86.715,57.33
X$10404 311 41 312 644 645 cell_1rw
* cell instance $10405 m0 *1 87.42,57.33
X$10405 313 41 314 644 645 cell_1rw
* cell instance $10406 m0 *1 88.125,57.33
X$10406 315 41 316 644 645 cell_1rw
* cell instance $10407 m0 *1 88.83,57.33
X$10407 317 41 318 644 645 cell_1rw
* cell instance $10408 m0 *1 89.535,57.33
X$10408 319 41 320 644 645 cell_1rw
* cell instance $10409 m0 *1 90.24,57.33
X$10409 321 41 323 644 645 cell_1rw
* cell instance $10410 m0 *1 90.945,57.33
X$10410 324 41 325 644 645 cell_1rw
* cell instance $10411 m0 *1 91.65,57.33
X$10411 326 41 327 644 645 cell_1rw
* cell instance $10412 m0 *1 92.355,57.33
X$10412 328 41 329 644 645 cell_1rw
* cell instance $10413 m0 *1 93.06,57.33
X$10413 330 41 331 644 645 cell_1rw
* cell instance $10414 m0 *1 93.765,57.33
X$10414 332 41 333 644 645 cell_1rw
* cell instance $10415 m0 *1 94.47,57.33
X$10415 334 41 335 644 645 cell_1rw
* cell instance $10416 m0 *1 95.175,57.33
X$10416 336 41 337 644 645 cell_1rw
* cell instance $10417 m0 *1 95.88,57.33
X$10417 338 41 339 644 645 cell_1rw
* cell instance $10418 m0 *1 96.585,57.33
X$10418 340 41 341 644 645 cell_1rw
* cell instance $10419 m0 *1 97.29,57.33
X$10419 342 41 343 644 645 cell_1rw
* cell instance $10420 m0 *1 97.995,57.33
X$10420 344 41 345 644 645 cell_1rw
* cell instance $10421 m0 *1 98.7,57.33
X$10421 346 41 347 644 645 cell_1rw
* cell instance $10422 m0 *1 99.405,57.33
X$10422 348 41 349 644 645 cell_1rw
* cell instance $10423 m0 *1 100.11,57.33
X$10423 350 41 351 644 645 cell_1rw
* cell instance $10424 m0 *1 100.815,57.33
X$10424 352 41 353 644 645 cell_1rw
* cell instance $10425 m0 *1 101.52,57.33
X$10425 354 41 355 644 645 cell_1rw
* cell instance $10426 m0 *1 102.225,57.33
X$10426 356 41 357 644 645 cell_1rw
* cell instance $10427 m0 *1 102.93,57.33
X$10427 358 41 359 644 645 cell_1rw
* cell instance $10428 m0 *1 103.635,57.33
X$10428 360 41 361 644 645 cell_1rw
* cell instance $10429 m0 *1 104.34,57.33
X$10429 362 41 363 644 645 cell_1rw
* cell instance $10430 m0 *1 105.045,57.33
X$10430 364 41 365 644 645 cell_1rw
* cell instance $10431 m0 *1 105.75,57.33
X$10431 366 41 367 644 645 cell_1rw
* cell instance $10432 m0 *1 106.455,57.33
X$10432 368 41 369 644 645 cell_1rw
* cell instance $10433 m0 *1 107.16,57.33
X$10433 370 41 371 644 645 cell_1rw
* cell instance $10434 m0 *1 107.865,57.33
X$10434 372 41 373 644 645 cell_1rw
* cell instance $10435 m0 *1 108.57,57.33
X$10435 374 41 375 644 645 cell_1rw
* cell instance $10436 m0 *1 109.275,57.33
X$10436 376 41 377 644 645 cell_1rw
* cell instance $10437 m0 *1 109.98,57.33
X$10437 378 41 379 644 645 cell_1rw
* cell instance $10438 m0 *1 110.685,57.33
X$10438 380 41 381 644 645 cell_1rw
* cell instance $10439 m0 *1 111.39,57.33
X$10439 382 41 383 644 645 cell_1rw
* cell instance $10440 m0 *1 112.095,57.33
X$10440 384 41 385 644 645 cell_1rw
* cell instance $10441 m0 *1 112.8,57.33
X$10441 386 41 387 644 645 cell_1rw
* cell instance $10442 m0 *1 113.505,57.33
X$10442 388 41 389 644 645 cell_1rw
* cell instance $10443 m0 *1 114.21,57.33
X$10443 390 41 391 644 645 cell_1rw
* cell instance $10444 m0 *1 114.915,57.33
X$10444 392 41 393 644 645 cell_1rw
* cell instance $10445 m0 *1 115.62,57.33
X$10445 394 41 395 644 645 cell_1rw
* cell instance $10446 m0 *1 116.325,57.33
X$10446 396 41 397 644 645 cell_1rw
* cell instance $10447 m0 *1 117.03,57.33
X$10447 398 41 399 644 645 cell_1rw
* cell instance $10448 m0 *1 117.735,57.33
X$10448 400 41 401 644 645 cell_1rw
* cell instance $10449 m0 *1 118.44,57.33
X$10449 402 41 403 644 645 cell_1rw
* cell instance $10450 m0 *1 119.145,57.33
X$10450 404 41 405 644 645 cell_1rw
* cell instance $10451 m0 *1 119.85,57.33
X$10451 406 41 407 644 645 cell_1rw
* cell instance $10452 m0 *1 120.555,57.33
X$10452 408 41 409 644 645 cell_1rw
* cell instance $10453 m0 *1 121.26,57.33
X$10453 410 41 411 644 645 cell_1rw
* cell instance $10454 m0 *1 121.965,57.33
X$10454 412 41 413 644 645 cell_1rw
* cell instance $10455 m0 *1 122.67,57.33
X$10455 414 41 415 644 645 cell_1rw
* cell instance $10456 m0 *1 123.375,57.33
X$10456 416 41 417 644 645 cell_1rw
* cell instance $10457 m0 *1 124.08,57.33
X$10457 418 41 419 644 645 cell_1rw
* cell instance $10458 m0 *1 124.785,57.33
X$10458 420 41 421 644 645 cell_1rw
* cell instance $10459 m0 *1 125.49,57.33
X$10459 422 41 423 644 645 cell_1rw
* cell instance $10460 m0 *1 126.195,57.33
X$10460 424 41 425 644 645 cell_1rw
* cell instance $10461 m0 *1 126.9,57.33
X$10461 426 41 427 644 645 cell_1rw
* cell instance $10462 m0 *1 127.605,57.33
X$10462 428 41 429 644 645 cell_1rw
* cell instance $10463 m0 *1 128.31,57.33
X$10463 430 41 431 644 645 cell_1rw
* cell instance $10464 m0 *1 129.015,57.33
X$10464 432 41 433 644 645 cell_1rw
* cell instance $10465 m0 *1 129.72,57.33
X$10465 434 41 435 644 645 cell_1rw
* cell instance $10466 m0 *1 130.425,57.33
X$10466 436 41 437 644 645 cell_1rw
* cell instance $10467 m0 *1 131.13,57.33
X$10467 438 41 439 644 645 cell_1rw
* cell instance $10468 m0 *1 131.835,57.33
X$10468 440 41 441 644 645 cell_1rw
* cell instance $10469 m0 *1 132.54,57.33
X$10469 442 41 443 644 645 cell_1rw
* cell instance $10470 m0 *1 133.245,57.33
X$10470 444 41 445 644 645 cell_1rw
* cell instance $10471 m0 *1 133.95,57.33
X$10471 446 41 447 644 645 cell_1rw
* cell instance $10472 m0 *1 134.655,57.33
X$10472 448 41 449 644 645 cell_1rw
* cell instance $10473 m0 *1 135.36,57.33
X$10473 450 41 451 644 645 cell_1rw
* cell instance $10474 m0 *1 136.065,57.33
X$10474 452 41 453 644 645 cell_1rw
* cell instance $10475 m0 *1 136.77,57.33
X$10475 454 41 455 644 645 cell_1rw
* cell instance $10476 m0 *1 137.475,57.33
X$10476 456 41 457 644 645 cell_1rw
* cell instance $10477 m0 *1 138.18,57.33
X$10477 458 41 459 644 645 cell_1rw
* cell instance $10478 m0 *1 138.885,57.33
X$10478 460 41 461 644 645 cell_1rw
* cell instance $10479 m0 *1 139.59,57.33
X$10479 462 41 463 644 645 cell_1rw
* cell instance $10480 m0 *1 140.295,57.33
X$10480 464 41 465 644 645 cell_1rw
* cell instance $10481 m0 *1 141,57.33
X$10481 466 41 467 644 645 cell_1rw
* cell instance $10482 m0 *1 141.705,57.33
X$10482 468 41 469 644 645 cell_1rw
* cell instance $10483 m0 *1 142.41,57.33
X$10483 470 41 471 644 645 cell_1rw
* cell instance $10484 m0 *1 143.115,57.33
X$10484 472 41 473 644 645 cell_1rw
* cell instance $10485 m0 *1 143.82,57.33
X$10485 474 41 475 644 645 cell_1rw
* cell instance $10486 m0 *1 144.525,57.33
X$10486 476 41 477 644 645 cell_1rw
* cell instance $10487 m0 *1 145.23,57.33
X$10487 478 41 479 644 645 cell_1rw
* cell instance $10488 m0 *1 145.935,57.33
X$10488 480 41 481 644 645 cell_1rw
* cell instance $10489 m0 *1 146.64,57.33
X$10489 482 41 483 644 645 cell_1rw
* cell instance $10490 m0 *1 147.345,57.33
X$10490 484 41 485 644 645 cell_1rw
* cell instance $10491 m0 *1 148.05,57.33
X$10491 486 41 487 644 645 cell_1rw
* cell instance $10492 m0 *1 148.755,57.33
X$10492 488 41 489 644 645 cell_1rw
* cell instance $10493 m0 *1 149.46,57.33
X$10493 490 41 491 644 645 cell_1rw
* cell instance $10494 m0 *1 150.165,57.33
X$10494 492 41 493 644 645 cell_1rw
* cell instance $10495 m0 *1 150.87,57.33
X$10495 494 41 495 644 645 cell_1rw
* cell instance $10496 m0 *1 151.575,57.33
X$10496 496 41 497 644 645 cell_1rw
* cell instance $10497 m0 *1 152.28,57.33
X$10497 498 41 499 644 645 cell_1rw
* cell instance $10498 m0 *1 152.985,57.33
X$10498 500 41 501 644 645 cell_1rw
* cell instance $10499 m0 *1 153.69,57.33
X$10499 502 41 503 644 645 cell_1rw
* cell instance $10500 m0 *1 154.395,57.33
X$10500 504 41 505 644 645 cell_1rw
* cell instance $10501 m0 *1 155.1,57.33
X$10501 506 41 507 644 645 cell_1rw
* cell instance $10502 m0 *1 155.805,57.33
X$10502 508 41 509 644 645 cell_1rw
* cell instance $10503 m0 *1 156.51,57.33
X$10503 510 41 511 644 645 cell_1rw
* cell instance $10504 m0 *1 157.215,57.33
X$10504 512 41 513 644 645 cell_1rw
* cell instance $10505 m0 *1 157.92,57.33
X$10505 514 41 515 644 645 cell_1rw
* cell instance $10506 m0 *1 158.625,57.33
X$10506 516 41 517 644 645 cell_1rw
* cell instance $10507 m0 *1 159.33,57.33
X$10507 518 41 519 644 645 cell_1rw
* cell instance $10508 m0 *1 160.035,57.33
X$10508 520 41 521 644 645 cell_1rw
* cell instance $10509 m0 *1 160.74,57.33
X$10509 522 41 523 644 645 cell_1rw
* cell instance $10510 m0 *1 161.445,57.33
X$10510 524 41 525 644 645 cell_1rw
* cell instance $10511 m0 *1 162.15,57.33
X$10511 526 41 527 644 645 cell_1rw
* cell instance $10512 m0 *1 162.855,57.33
X$10512 528 41 529 644 645 cell_1rw
* cell instance $10513 m0 *1 163.56,57.33
X$10513 530 41 531 644 645 cell_1rw
* cell instance $10514 m0 *1 164.265,57.33
X$10514 532 41 533 644 645 cell_1rw
* cell instance $10515 m0 *1 164.97,57.33
X$10515 534 41 535 644 645 cell_1rw
* cell instance $10516 m0 *1 165.675,57.33
X$10516 536 41 537 644 645 cell_1rw
* cell instance $10517 m0 *1 166.38,57.33
X$10517 538 41 539 644 645 cell_1rw
* cell instance $10518 m0 *1 167.085,57.33
X$10518 540 41 541 644 645 cell_1rw
* cell instance $10519 m0 *1 167.79,57.33
X$10519 542 41 543 644 645 cell_1rw
* cell instance $10520 m0 *1 168.495,57.33
X$10520 544 41 545 644 645 cell_1rw
* cell instance $10521 m0 *1 169.2,57.33
X$10521 546 41 547 644 645 cell_1rw
* cell instance $10522 m0 *1 169.905,57.33
X$10522 548 41 549 644 645 cell_1rw
* cell instance $10523 m0 *1 170.61,57.33
X$10523 550 41 551 644 645 cell_1rw
* cell instance $10524 m0 *1 171.315,57.33
X$10524 552 41 553 644 645 cell_1rw
* cell instance $10525 m0 *1 172.02,57.33
X$10525 554 41 555 644 645 cell_1rw
* cell instance $10526 m0 *1 172.725,57.33
X$10526 556 41 557 644 645 cell_1rw
* cell instance $10527 m0 *1 173.43,57.33
X$10527 558 41 559 644 645 cell_1rw
* cell instance $10528 m0 *1 174.135,57.33
X$10528 560 41 561 644 645 cell_1rw
* cell instance $10529 m0 *1 174.84,57.33
X$10529 562 41 563 644 645 cell_1rw
* cell instance $10530 m0 *1 175.545,57.33
X$10530 564 41 565 644 645 cell_1rw
* cell instance $10531 m0 *1 176.25,57.33
X$10531 566 41 567 644 645 cell_1rw
* cell instance $10532 m0 *1 176.955,57.33
X$10532 568 41 569 644 645 cell_1rw
* cell instance $10533 m0 *1 177.66,57.33
X$10533 570 41 571 644 645 cell_1rw
* cell instance $10534 m0 *1 178.365,57.33
X$10534 572 41 573 644 645 cell_1rw
* cell instance $10535 m0 *1 179.07,57.33
X$10535 574 41 575 644 645 cell_1rw
* cell instance $10536 m0 *1 179.775,57.33
X$10536 576 41 577 644 645 cell_1rw
* cell instance $10537 m0 *1 180.48,57.33
X$10537 578 41 579 644 645 cell_1rw
* cell instance $10538 r0 *1 0.705,54.6
X$10538 67 42 68 644 645 cell_1rw
* cell instance $10539 r0 *1 0,54.6
X$10539 65 42 66 644 645 cell_1rw
* cell instance $10540 r0 *1 1.41,54.6
X$10540 69 42 70 644 645 cell_1rw
* cell instance $10541 r0 *1 2.115,54.6
X$10541 71 42 72 644 645 cell_1rw
* cell instance $10542 r0 *1 2.82,54.6
X$10542 73 42 74 644 645 cell_1rw
* cell instance $10543 r0 *1 3.525,54.6
X$10543 75 42 76 644 645 cell_1rw
* cell instance $10544 r0 *1 4.23,54.6
X$10544 77 42 78 644 645 cell_1rw
* cell instance $10545 r0 *1 4.935,54.6
X$10545 79 42 80 644 645 cell_1rw
* cell instance $10546 r0 *1 5.64,54.6
X$10546 81 42 82 644 645 cell_1rw
* cell instance $10547 r0 *1 6.345,54.6
X$10547 83 42 84 644 645 cell_1rw
* cell instance $10548 r0 *1 7.05,54.6
X$10548 85 42 86 644 645 cell_1rw
* cell instance $10549 r0 *1 7.755,54.6
X$10549 87 42 88 644 645 cell_1rw
* cell instance $10550 r0 *1 8.46,54.6
X$10550 89 42 90 644 645 cell_1rw
* cell instance $10551 r0 *1 9.165,54.6
X$10551 91 42 92 644 645 cell_1rw
* cell instance $10552 r0 *1 9.87,54.6
X$10552 93 42 94 644 645 cell_1rw
* cell instance $10553 r0 *1 10.575,54.6
X$10553 95 42 96 644 645 cell_1rw
* cell instance $10554 r0 *1 11.28,54.6
X$10554 97 42 98 644 645 cell_1rw
* cell instance $10555 r0 *1 11.985,54.6
X$10555 99 42 100 644 645 cell_1rw
* cell instance $10556 r0 *1 12.69,54.6
X$10556 101 42 102 644 645 cell_1rw
* cell instance $10557 r0 *1 13.395,54.6
X$10557 103 42 104 644 645 cell_1rw
* cell instance $10558 r0 *1 14.1,54.6
X$10558 105 42 106 644 645 cell_1rw
* cell instance $10559 r0 *1 14.805,54.6
X$10559 107 42 108 644 645 cell_1rw
* cell instance $10560 r0 *1 15.51,54.6
X$10560 109 42 110 644 645 cell_1rw
* cell instance $10561 r0 *1 16.215,54.6
X$10561 111 42 112 644 645 cell_1rw
* cell instance $10562 r0 *1 16.92,54.6
X$10562 113 42 114 644 645 cell_1rw
* cell instance $10563 r0 *1 17.625,54.6
X$10563 115 42 116 644 645 cell_1rw
* cell instance $10564 r0 *1 18.33,54.6
X$10564 117 42 118 644 645 cell_1rw
* cell instance $10565 r0 *1 19.035,54.6
X$10565 119 42 120 644 645 cell_1rw
* cell instance $10566 r0 *1 19.74,54.6
X$10566 121 42 122 644 645 cell_1rw
* cell instance $10567 r0 *1 20.445,54.6
X$10567 123 42 124 644 645 cell_1rw
* cell instance $10568 r0 *1 21.15,54.6
X$10568 125 42 126 644 645 cell_1rw
* cell instance $10569 r0 *1 21.855,54.6
X$10569 127 42 128 644 645 cell_1rw
* cell instance $10570 r0 *1 22.56,54.6
X$10570 129 42 130 644 645 cell_1rw
* cell instance $10571 r0 *1 23.265,54.6
X$10571 131 42 132 644 645 cell_1rw
* cell instance $10572 r0 *1 23.97,54.6
X$10572 133 42 134 644 645 cell_1rw
* cell instance $10573 r0 *1 24.675,54.6
X$10573 135 42 136 644 645 cell_1rw
* cell instance $10574 r0 *1 25.38,54.6
X$10574 137 42 138 644 645 cell_1rw
* cell instance $10575 r0 *1 26.085,54.6
X$10575 139 42 140 644 645 cell_1rw
* cell instance $10576 r0 *1 26.79,54.6
X$10576 141 42 142 644 645 cell_1rw
* cell instance $10577 r0 *1 27.495,54.6
X$10577 143 42 144 644 645 cell_1rw
* cell instance $10578 r0 *1 28.2,54.6
X$10578 145 42 146 644 645 cell_1rw
* cell instance $10579 r0 *1 28.905,54.6
X$10579 147 42 148 644 645 cell_1rw
* cell instance $10580 r0 *1 29.61,54.6
X$10580 149 42 150 644 645 cell_1rw
* cell instance $10581 r0 *1 30.315,54.6
X$10581 151 42 152 644 645 cell_1rw
* cell instance $10582 r0 *1 31.02,54.6
X$10582 153 42 154 644 645 cell_1rw
* cell instance $10583 r0 *1 31.725,54.6
X$10583 155 42 156 644 645 cell_1rw
* cell instance $10584 r0 *1 32.43,54.6
X$10584 157 42 158 644 645 cell_1rw
* cell instance $10585 r0 *1 33.135,54.6
X$10585 159 42 160 644 645 cell_1rw
* cell instance $10586 r0 *1 33.84,54.6
X$10586 161 42 162 644 645 cell_1rw
* cell instance $10587 r0 *1 34.545,54.6
X$10587 163 42 164 644 645 cell_1rw
* cell instance $10588 r0 *1 35.25,54.6
X$10588 165 42 166 644 645 cell_1rw
* cell instance $10589 r0 *1 35.955,54.6
X$10589 167 42 168 644 645 cell_1rw
* cell instance $10590 r0 *1 36.66,54.6
X$10590 169 42 170 644 645 cell_1rw
* cell instance $10591 r0 *1 37.365,54.6
X$10591 171 42 172 644 645 cell_1rw
* cell instance $10592 r0 *1 38.07,54.6
X$10592 173 42 174 644 645 cell_1rw
* cell instance $10593 r0 *1 38.775,54.6
X$10593 175 42 176 644 645 cell_1rw
* cell instance $10594 r0 *1 39.48,54.6
X$10594 177 42 178 644 645 cell_1rw
* cell instance $10595 r0 *1 40.185,54.6
X$10595 179 42 180 644 645 cell_1rw
* cell instance $10596 r0 *1 40.89,54.6
X$10596 181 42 182 644 645 cell_1rw
* cell instance $10597 r0 *1 41.595,54.6
X$10597 183 42 184 644 645 cell_1rw
* cell instance $10598 r0 *1 42.3,54.6
X$10598 185 42 186 644 645 cell_1rw
* cell instance $10599 r0 *1 43.005,54.6
X$10599 187 42 188 644 645 cell_1rw
* cell instance $10600 r0 *1 43.71,54.6
X$10600 189 42 190 644 645 cell_1rw
* cell instance $10601 r0 *1 44.415,54.6
X$10601 191 42 192 644 645 cell_1rw
* cell instance $10602 r0 *1 45.12,54.6
X$10602 193 42 194 644 645 cell_1rw
* cell instance $10603 r0 *1 45.825,54.6
X$10603 195 42 196 644 645 cell_1rw
* cell instance $10604 r0 *1 46.53,54.6
X$10604 197 42 198 644 645 cell_1rw
* cell instance $10605 r0 *1 47.235,54.6
X$10605 199 42 200 644 645 cell_1rw
* cell instance $10606 r0 *1 47.94,54.6
X$10606 201 42 202 644 645 cell_1rw
* cell instance $10607 r0 *1 48.645,54.6
X$10607 203 42 204 644 645 cell_1rw
* cell instance $10608 r0 *1 49.35,54.6
X$10608 205 42 206 644 645 cell_1rw
* cell instance $10609 r0 *1 50.055,54.6
X$10609 207 42 208 644 645 cell_1rw
* cell instance $10610 r0 *1 50.76,54.6
X$10610 209 42 210 644 645 cell_1rw
* cell instance $10611 r0 *1 51.465,54.6
X$10611 211 42 212 644 645 cell_1rw
* cell instance $10612 r0 *1 52.17,54.6
X$10612 213 42 214 644 645 cell_1rw
* cell instance $10613 r0 *1 52.875,54.6
X$10613 215 42 216 644 645 cell_1rw
* cell instance $10614 r0 *1 53.58,54.6
X$10614 217 42 218 644 645 cell_1rw
* cell instance $10615 r0 *1 54.285,54.6
X$10615 219 42 220 644 645 cell_1rw
* cell instance $10616 r0 *1 54.99,54.6
X$10616 221 42 222 644 645 cell_1rw
* cell instance $10617 r0 *1 55.695,54.6
X$10617 223 42 224 644 645 cell_1rw
* cell instance $10618 r0 *1 56.4,54.6
X$10618 225 42 226 644 645 cell_1rw
* cell instance $10619 r0 *1 57.105,54.6
X$10619 227 42 228 644 645 cell_1rw
* cell instance $10620 r0 *1 57.81,54.6
X$10620 229 42 230 644 645 cell_1rw
* cell instance $10621 r0 *1 58.515,54.6
X$10621 231 42 232 644 645 cell_1rw
* cell instance $10622 r0 *1 59.22,54.6
X$10622 233 42 234 644 645 cell_1rw
* cell instance $10623 r0 *1 59.925,54.6
X$10623 235 42 236 644 645 cell_1rw
* cell instance $10624 r0 *1 60.63,54.6
X$10624 237 42 238 644 645 cell_1rw
* cell instance $10625 r0 *1 61.335,54.6
X$10625 239 42 240 644 645 cell_1rw
* cell instance $10626 r0 *1 62.04,54.6
X$10626 241 42 242 644 645 cell_1rw
* cell instance $10627 r0 *1 62.745,54.6
X$10627 243 42 244 644 645 cell_1rw
* cell instance $10628 r0 *1 63.45,54.6
X$10628 245 42 246 644 645 cell_1rw
* cell instance $10629 r0 *1 64.155,54.6
X$10629 247 42 248 644 645 cell_1rw
* cell instance $10630 r0 *1 64.86,54.6
X$10630 249 42 250 644 645 cell_1rw
* cell instance $10631 r0 *1 65.565,54.6
X$10631 251 42 252 644 645 cell_1rw
* cell instance $10632 r0 *1 66.27,54.6
X$10632 253 42 254 644 645 cell_1rw
* cell instance $10633 r0 *1 66.975,54.6
X$10633 255 42 256 644 645 cell_1rw
* cell instance $10634 r0 *1 67.68,54.6
X$10634 257 42 258 644 645 cell_1rw
* cell instance $10635 r0 *1 68.385,54.6
X$10635 259 42 260 644 645 cell_1rw
* cell instance $10636 r0 *1 69.09,54.6
X$10636 261 42 262 644 645 cell_1rw
* cell instance $10637 r0 *1 69.795,54.6
X$10637 263 42 264 644 645 cell_1rw
* cell instance $10638 r0 *1 70.5,54.6
X$10638 265 42 266 644 645 cell_1rw
* cell instance $10639 r0 *1 71.205,54.6
X$10639 267 42 268 644 645 cell_1rw
* cell instance $10640 r0 *1 71.91,54.6
X$10640 269 42 270 644 645 cell_1rw
* cell instance $10641 r0 *1 72.615,54.6
X$10641 271 42 272 644 645 cell_1rw
* cell instance $10642 r0 *1 73.32,54.6
X$10642 273 42 274 644 645 cell_1rw
* cell instance $10643 r0 *1 74.025,54.6
X$10643 275 42 276 644 645 cell_1rw
* cell instance $10644 r0 *1 74.73,54.6
X$10644 277 42 278 644 645 cell_1rw
* cell instance $10645 r0 *1 75.435,54.6
X$10645 279 42 280 644 645 cell_1rw
* cell instance $10646 r0 *1 76.14,54.6
X$10646 281 42 282 644 645 cell_1rw
* cell instance $10647 r0 *1 76.845,54.6
X$10647 283 42 284 644 645 cell_1rw
* cell instance $10648 r0 *1 77.55,54.6
X$10648 285 42 286 644 645 cell_1rw
* cell instance $10649 r0 *1 78.255,54.6
X$10649 287 42 288 644 645 cell_1rw
* cell instance $10650 r0 *1 78.96,54.6
X$10650 289 42 290 644 645 cell_1rw
* cell instance $10651 r0 *1 79.665,54.6
X$10651 291 42 292 644 645 cell_1rw
* cell instance $10652 r0 *1 80.37,54.6
X$10652 293 42 294 644 645 cell_1rw
* cell instance $10653 r0 *1 81.075,54.6
X$10653 295 42 296 644 645 cell_1rw
* cell instance $10654 r0 *1 81.78,54.6
X$10654 297 42 298 644 645 cell_1rw
* cell instance $10655 r0 *1 82.485,54.6
X$10655 299 42 300 644 645 cell_1rw
* cell instance $10656 r0 *1 83.19,54.6
X$10656 301 42 302 644 645 cell_1rw
* cell instance $10657 r0 *1 83.895,54.6
X$10657 303 42 304 644 645 cell_1rw
* cell instance $10658 r0 *1 84.6,54.6
X$10658 305 42 306 644 645 cell_1rw
* cell instance $10659 r0 *1 85.305,54.6
X$10659 307 42 308 644 645 cell_1rw
* cell instance $10660 r0 *1 86.01,54.6
X$10660 309 42 310 644 645 cell_1rw
* cell instance $10661 r0 *1 86.715,54.6
X$10661 311 42 312 644 645 cell_1rw
* cell instance $10662 r0 *1 87.42,54.6
X$10662 313 42 314 644 645 cell_1rw
* cell instance $10663 r0 *1 88.125,54.6
X$10663 315 42 316 644 645 cell_1rw
* cell instance $10664 r0 *1 88.83,54.6
X$10664 317 42 318 644 645 cell_1rw
* cell instance $10665 r0 *1 89.535,54.6
X$10665 319 42 320 644 645 cell_1rw
* cell instance $10666 r0 *1 90.24,54.6
X$10666 321 42 323 644 645 cell_1rw
* cell instance $10667 r0 *1 90.945,54.6
X$10667 324 42 325 644 645 cell_1rw
* cell instance $10668 r0 *1 91.65,54.6
X$10668 326 42 327 644 645 cell_1rw
* cell instance $10669 r0 *1 92.355,54.6
X$10669 328 42 329 644 645 cell_1rw
* cell instance $10670 r0 *1 93.06,54.6
X$10670 330 42 331 644 645 cell_1rw
* cell instance $10671 r0 *1 93.765,54.6
X$10671 332 42 333 644 645 cell_1rw
* cell instance $10672 r0 *1 94.47,54.6
X$10672 334 42 335 644 645 cell_1rw
* cell instance $10673 r0 *1 95.175,54.6
X$10673 336 42 337 644 645 cell_1rw
* cell instance $10674 r0 *1 95.88,54.6
X$10674 338 42 339 644 645 cell_1rw
* cell instance $10675 r0 *1 96.585,54.6
X$10675 340 42 341 644 645 cell_1rw
* cell instance $10676 r0 *1 97.29,54.6
X$10676 342 42 343 644 645 cell_1rw
* cell instance $10677 r0 *1 97.995,54.6
X$10677 344 42 345 644 645 cell_1rw
* cell instance $10678 r0 *1 98.7,54.6
X$10678 346 42 347 644 645 cell_1rw
* cell instance $10679 r0 *1 99.405,54.6
X$10679 348 42 349 644 645 cell_1rw
* cell instance $10680 r0 *1 100.11,54.6
X$10680 350 42 351 644 645 cell_1rw
* cell instance $10681 r0 *1 100.815,54.6
X$10681 352 42 353 644 645 cell_1rw
* cell instance $10682 r0 *1 101.52,54.6
X$10682 354 42 355 644 645 cell_1rw
* cell instance $10683 r0 *1 102.225,54.6
X$10683 356 42 357 644 645 cell_1rw
* cell instance $10684 r0 *1 102.93,54.6
X$10684 358 42 359 644 645 cell_1rw
* cell instance $10685 r0 *1 103.635,54.6
X$10685 360 42 361 644 645 cell_1rw
* cell instance $10686 r0 *1 104.34,54.6
X$10686 362 42 363 644 645 cell_1rw
* cell instance $10687 r0 *1 105.045,54.6
X$10687 364 42 365 644 645 cell_1rw
* cell instance $10688 r0 *1 105.75,54.6
X$10688 366 42 367 644 645 cell_1rw
* cell instance $10689 r0 *1 106.455,54.6
X$10689 368 42 369 644 645 cell_1rw
* cell instance $10690 r0 *1 107.16,54.6
X$10690 370 42 371 644 645 cell_1rw
* cell instance $10691 r0 *1 107.865,54.6
X$10691 372 42 373 644 645 cell_1rw
* cell instance $10692 r0 *1 108.57,54.6
X$10692 374 42 375 644 645 cell_1rw
* cell instance $10693 r0 *1 109.275,54.6
X$10693 376 42 377 644 645 cell_1rw
* cell instance $10694 r0 *1 109.98,54.6
X$10694 378 42 379 644 645 cell_1rw
* cell instance $10695 r0 *1 110.685,54.6
X$10695 380 42 381 644 645 cell_1rw
* cell instance $10696 r0 *1 111.39,54.6
X$10696 382 42 383 644 645 cell_1rw
* cell instance $10697 r0 *1 112.095,54.6
X$10697 384 42 385 644 645 cell_1rw
* cell instance $10698 r0 *1 112.8,54.6
X$10698 386 42 387 644 645 cell_1rw
* cell instance $10699 r0 *1 113.505,54.6
X$10699 388 42 389 644 645 cell_1rw
* cell instance $10700 r0 *1 114.21,54.6
X$10700 390 42 391 644 645 cell_1rw
* cell instance $10701 r0 *1 114.915,54.6
X$10701 392 42 393 644 645 cell_1rw
* cell instance $10702 r0 *1 115.62,54.6
X$10702 394 42 395 644 645 cell_1rw
* cell instance $10703 r0 *1 116.325,54.6
X$10703 396 42 397 644 645 cell_1rw
* cell instance $10704 r0 *1 117.03,54.6
X$10704 398 42 399 644 645 cell_1rw
* cell instance $10705 r0 *1 117.735,54.6
X$10705 400 42 401 644 645 cell_1rw
* cell instance $10706 r0 *1 118.44,54.6
X$10706 402 42 403 644 645 cell_1rw
* cell instance $10707 r0 *1 119.145,54.6
X$10707 404 42 405 644 645 cell_1rw
* cell instance $10708 r0 *1 119.85,54.6
X$10708 406 42 407 644 645 cell_1rw
* cell instance $10709 r0 *1 120.555,54.6
X$10709 408 42 409 644 645 cell_1rw
* cell instance $10710 r0 *1 121.26,54.6
X$10710 410 42 411 644 645 cell_1rw
* cell instance $10711 r0 *1 121.965,54.6
X$10711 412 42 413 644 645 cell_1rw
* cell instance $10712 r0 *1 122.67,54.6
X$10712 414 42 415 644 645 cell_1rw
* cell instance $10713 r0 *1 123.375,54.6
X$10713 416 42 417 644 645 cell_1rw
* cell instance $10714 r0 *1 124.08,54.6
X$10714 418 42 419 644 645 cell_1rw
* cell instance $10715 r0 *1 124.785,54.6
X$10715 420 42 421 644 645 cell_1rw
* cell instance $10716 r0 *1 125.49,54.6
X$10716 422 42 423 644 645 cell_1rw
* cell instance $10717 r0 *1 126.195,54.6
X$10717 424 42 425 644 645 cell_1rw
* cell instance $10718 r0 *1 126.9,54.6
X$10718 426 42 427 644 645 cell_1rw
* cell instance $10719 r0 *1 127.605,54.6
X$10719 428 42 429 644 645 cell_1rw
* cell instance $10720 r0 *1 128.31,54.6
X$10720 430 42 431 644 645 cell_1rw
* cell instance $10721 r0 *1 129.015,54.6
X$10721 432 42 433 644 645 cell_1rw
* cell instance $10722 r0 *1 129.72,54.6
X$10722 434 42 435 644 645 cell_1rw
* cell instance $10723 r0 *1 130.425,54.6
X$10723 436 42 437 644 645 cell_1rw
* cell instance $10724 r0 *1 131.13,54.6
X$10724 438 42 439 644 645 cell_1rw
* cell instance $10725 r0 *1 131.835,54.6
X$10725 440 42 441 644 645 cell_1rw
* cell instance $10726 r0 *1 132.54,54.6
X$10726 442 42 443 644 645 cell_1rw
* cell instance $10727 r0 *1 133.245,54.6
X$10727 444 42 445 644 645 cell_1rw
* cell instance $10728 r0 *1 133.95,54.6
X$10728 446 42 447 644 645 cell_1rw
* cell instance $10729 r0 *1 134.655,54.6
X$10729 448 42 449 644 645 cell_1rw
* cell instance $10730 r0 *1 135.36,54.6
X$10730 450 42 451 644 645 cell_1rw
* cell instance $10731 r0 *1 136.065,54.6
X$10731 452 42 453 644 645 cell_1rw
* cell instance $10732 r0 *1 136.77,54.6
X$10732 454 42 455 644 645 cell_1rw
* cell instance $10733 r0 *1 137.475,54.6
X$10733 456 42 457 644 645 cell_1rw
* cell instance $10734 r0 *1 138.18,54.6
X$10734 458 42 459 644 645 cell_1rw
* cell instance $10735 r0 *1 138.885,54.6
X$10735 460 42 461 644 645 cell_1rw
* cell instance $10736 r0 *1 139.59,54.6
X$10736 462 42 463 644 645 cell_1rw
* cell instance $10737 r0 *1 140.295,54.6
X$10737 464 42 465 644 645 cell_1rw
* cell instance $10738 r0 *1 141,54.6
X$10738 466 42 467 644 645 cell_1rw
* cell instance $10739 r0 *1 141.705,54.6
X$10739 468 42 469 644 645 cell_1rw
* cell instance $10740 r0 *1 142.41,54.6
X$10740 470 42 471 644 645 cell_1rw
* cell instance $10741 r0 *1 143.115,54.6
X$10741 472 42 473 644 645 cell_1rw
* cell instance $10742 r0 *1 143.82,54.6
X$10742 474 42 475 644 645 cell_1rw
* cell instance $10743 r0 *1 144.525,54.6
X$10743 476 42 477 644 645 cell_1rw
* cell instance $10744 r0 *1 145.23,54.6
X$10744 478 42 479 644 645 cell_1rw
* cell instance $10745 r0 *1 145.935,54.6
X$10745 480 42 481 644 645 cell_1rw
* cell instance $10746 r0 *1 146.64,54.6
X$10746 482 42 483 644 645 cell_1rw
* cell instance $10747 r0 *1 147.345,54.6
X$10747 484 42 485 644 645 cell_1rw
* cell instance $10748 r0 *1 148.05,54.6
X$10748 486 42 487 644 645 cell_1rw
* cell instance $10749 r0 *1 148.755,54.6
X$10749 488 42 489 644 645 cell_1rw
* cell instance $10750 r0 *1 149.46,54.6
X$10750 490 42 491 644 645 cell_1rw
* cell instance $10751 r0 *1 150.165,54.6
X$10751 492 42 493 644 645 cell_1rw
* cell instance $10752 r0 *1 150.87,54.6
X$10752 494 42 495 644 645 cell_1rw
* cell instance $10753 r0 *1 151.575,54.6
X$10753 496 42 497 644 645 cell_1rw
* cell instance $10754 r0 *1 152.28,54.6
X$10754 498 42 499 644 645 cell_1rw
* cell instance $10755 r0 *1 152.985,54.6
X$10755 500 42 501 644 645 cell_1rw
* cell instance $10756 r0 *1 153.69,54.6
X$10756 502 42 503 644 645 cell_1rw
* cell instance $10757 r0 *1 154.395,54.6
X$10757 504 42 505 644 645 cell_1rw
* cell instance $10758 r0 *1 155.1,54.6
X$10758 506 42 507 644 645 cell_1rw
* cell instance $10759 r0 *1 155.805,54.6
X$10759 508 42 509 644 645 cell_1rw
* cell instance $10760 r0 *1 156.51,54.6
X$10760 510 42 511 644 645 cell_1rw
* cell instance $10761 r0 *1 157.215,54.6
X$10761 512 42 513 644 645 cell_1rw
* cell instance $10762 r0 *1 157.92,54.6
X$10762 514 42 515 644 645 cell_1rw
* cell instance $10763 r0 *1 158.625,54.6
X$10763 516 42 517 644 645 cell_1rw
* cell instance $10764 r0 *1 159.33,54.6
X$10764 518 42 519 644 645 cell_1rw
* cell instance $10765 r0 *1 160.035,54.6
X$10765 520 42 521 644 645 cell_1rw
* cell instance $10766 r0 *1 160.74,54.6
X$10766 522 42 523 644 645 cell_1rw
* cell instance $10767 r0 *1 161.445,54.6
X$10767 524 42 525 644 645 cell_1rw
* cell instance $10768 r0 *1 162.15,54.6
X$10768 526 42 527 644 645 cell_1rw
* cell instance $10769 r0 *1 162.855,54.6
X$10769 528 42 529 644 645 cell_1rw
* cell instance $10770 r0 *1 163.56,54.6
X$10770 530 42 531 644 645 cell_1rw
* cell instance $10771 r0 *1 164.265,54.6
X$10771 532 42 533 644 645 cell_1rw
* cell instance $10772 r0 *1 164.97,54.6
X$10772 534 42 535 644 645 cell_1rw
* cell instance $10773 r0 *1 165.675,54.6
X$10773 536 42 537 644 645 cell_1rw
* cell instance $10774 r0 *1 166.38,54.6
X$10774 538 42 539 644 645 cell_1rw
* cell instance $10775 r0 *1 167.085,54.6
X$10775 540 42 541 644 645 cell_1rw
* cell instance $10776 r0 *1 167.79,54.6
X$10776 542 42 543 644 645 cell_1rw
* cell instance $10777 r0 *1 168.495,54.6
X$10777 544 42 545 644 645 cell_1rw
* cell instance $10778 r0 *1 169.2,54.6
X$10778 546 42 547 644 645 cell_1rw
* cell instance $10779 r0 *1 169.905,54.6
X$10779 548 42 549 644 645 cell_1rw
* cell instance $10780 r0 *1 170.61,54.6
X$10780 550 42 551 644 645 cell_1rw
* cell instance $10781 r0 *1 171.315,54.6
X$10781 552 42 553 644 645 cell_1rw
* cell instance $10782 r0 *1 172.02,54.6
X$10782 554 42 555 644 645 cell_1rw
* cell instance $10783 r0 *1 172.725,54.6
X$10783 556 42 557 644 645 cell_1rw
* cell instance $10784 r0 *1 173.43,54.6
X$10784 558 42 559 644 645 cell_1rw
* cell instance $10785 r0 *1 174.135,54.6
X$10785 560 42 561 644 645 cell_1rw
* cell instance $10786 r0 *1 174.84,54.6
X$10786 562 42 563 644 645 cell_1rw
* cell instance $10787 r0 *1 175.545,54.6
X$10787 564 42 565 644 645 cell_1rw
* cell instance $10788 r0 *1 176.25,54.6
X$10788 566 42 567 644 645 cell_1rw
* cell instance $10789 r0 *1 176.955,54.6
X$10789 568 42 569 644 645 cell_1rw
* cell instance $10790 r0 *1 177.66,54.6
X$10790 570 42 571 644 645 cell_1rw
* cell instance $10791 r0 *1 178.365,54.6
X$10791 572 42 573 644 645 cell_1rw
* cell instance $10792 r0 *1 179.07,54.6
X$10792 574 42 575 644 645 cell_1rw
* cell instance $10793 r0 *1 179.775,54.6
X$10793 576 42 577 644 645 cell_1rw
* cell instance $10794 r0 *1 180.48,54.6
X$10794 578 42 579 644 645 cell_1rw
* cell instance $10795 m0 *1 0.705,60.06
X$10795 67 43 68 644 645 cell_1rw
* cell instance $10796 m0 *1 0,60.06
X$10796 65 43 66 644 645 cell_1rw
* cell instance $10797 m0 *1 1.41,60.06
X$10797 69 43 70 644 645 cell_1rw
* cell instance $10798 m0 *1 2.115,60.06
X$10798 71 43 72 644 645 cell_1rw
* cell instance $10799 m0 *1 2.82,60.06
X$10799 73 43 74 644 645 cell_1rw
* cell instance $10800 m0 *1 3.525,60.06
X$10800 75 43 76 644 645 cell_1rw
* cell instance $10801 m0 *1 4.23,60.06
X$10801 77 43 78 644 645 cell_1rw
* cell instance $10802 m0 *1 4.935,60.06
X$10802 79 43 80 644 645 cell_1rw
* cell instance $10803 m0 *1 5.64,60.06
X$10803 81 43 82 644 645 cell_1rw
* cell instance $10804 m0 *1 6.345,60.06
X$10804 83 43 84 644 645 cell_1rw
* cell instance $10805 m0 *1 7.05,60.06
X$10805 85 43 86 644 645 cell_1rw
* cell instance $10806 m0 *1 7.755,60.06
X$10806 87 43 88 644 645 cell_1rw
* cell instance $10807 m0 *1 8.46,60.06
X$10807 89 43 90 644 645 cell_1rw
* cell instance $10808 m0 *1 9.165,60.06
X$10808 91 43 92 644 645 cell_1rw
* cell instance $10809 m0 *1 9.87,60.06
X$10809 93 43 94 644 645 cell_1rw
* cell instance $10810 m0 *1 10.575,60.06
X$10810 95 43 96 644 645 cell_1rw
* cell instance $10811 m0 *1 11.28,60.06
X$10811 97 43 98 644 645 cell_1rw
* cell instance $10812 m0 *1 11.985,60.06
X$10812 99 43 100 644 645 cell_1rw
* cell instance $10813 m0 *1 12.69,60.06
X$10813 101 43 102 644 645 cell_1rw
* cell instance $10814 m0 *1 13.395,60.06
X$10814 103 43 104 644 645 cell_1rw
* cell instance $10815 m0 *1 14.1,60.06
X$10815 105 43 106 644 645 cell_1rw
* cell instance $10816 m0 *1 14.805,60.06
X$10816 107 43 108 644 645 cell_1rw
* cell instance $10817 m0 *1 15.51,60.06
X$10817 109 43 110 644 645 cell_1rw
* cell instance $10818 m0 *1 16.215,60.06
X$10818 111 43 112 644 645 cell_1rw
* cell instance $10819 m0 *1 16.92,60.06
X$10819 113 43 114 644 645 cell_1rw
* cell instance $10820 m0 *1 17.625,60.06
X$10820 115 43 116 644 645 cell_1rw
* cell instance $10821 m0 *1 18.33,60.06
X$10821 117 43 118 644 645 cell_1rw
* cell instance $10822 m0 *1 19.035,60.06
X$10822 119 43 120 644 645 cell_1rw
* cell instance $10823 m0 *1 19.74,60.06
X$10823 121 43 122 644 645 cell_1rw
* cell instance $10824 m0 *1 20.445,60.06
X$10824 123 43 124 644 645 cell_1rw
* cell instance $10825 m0 *1 21.15,60.06
X$10825 125 43 126 644 645 cell_1rw
* cell instance $10826 m0 *1 21.855,60.06
X$10826 127 43 128 644 645 cell_1rw
* cell instance $10827 m0 *1 22.56,60.06
X$10827 129 43 130 644 645 cell_1rw
* cell instance $10828 m0 *1 23.265,60.06
X$10828 131 43 132 644 645 cell_1rw
* cell instance $10829 m0 *1 23.97,60.06
X$10829 133 43 134 644 645 cell_1rw
* cell instance $10830 m0 *1 24.675,60.06
X$10830 135 43 136 644 645 cell_1rw
* cell instance $10831 m0 *1 25.38,60.06
X$10831 137 43 138 644 645 cell_1rw
* cell instance $10832 m0 *1 26.085,60.06
X$10832 139 43 140 644 645 cell_1rw
* cell instance $10833 m0 *1 26.79,60.06
X$10833 141 43 142 644 645 cell_1rw
* cell instance $10834 m0 *1 27.495,60.06
X$10834 143 43 144 644 645 cell_1rw
* cell instance $10835 m0 *1 28.2,60.06
X$10835 145 43 146 644 645 cell_1rw
* cell instance $10836 m0 *1 28.905,60.06
X$10836 147 43 148 644 645 cell_1rw
* cell instance $10837 m0 *1 29.61,60.06
X$10837 149 43 150 644 645 cell_1rw
* cell instance $10838 m0 *1 30.315,60.06
X$10838 151 43 152 644 645 cell_1rw
* cell instance $10839 m0 *1 31.02,60.06
X$10839 153 43 154 644 645 cell_1rw
* cell instance $10840 m0 *1 31.725,60.06
X$10840 155 43 156 644 645 cell_1rw
* cell instance $10841 m0 *1 32.43,60.06
X$10841 157 43 158 644 645 cell_1rw
* cell instance $10842 m0 *1 33.135,60.06
X$10842 159 43 160 644 645 cell_1rw
* cell instance $10843 m0 *1 33.84,60.06
X$10843 161 43 162 644 645 cell_1rw
* cell instance $10844 m0 *1 34.545,60.06
X$10844 163 43 164 644 645 cell_1rw
* cell instance $10845 m0 *1 35.25,60.06
X$10845 165 43 166 644 645 cell_1rw
* cell instance $10846 m0 *1 35.955,60.06
X$10846 167 43 168 644 645 cell_1rw
* cell instance $10847 m0 *1 36.66,60.06
X$10847 169 43 170 644 645 cell_1rw
* cell instance $10848 m0 *1 37.365,60.06
X$10848 171 43 172 644 645 cell_1rw
* cell instance $10849 m0 *1 38.07,60.06
X$10849 173 43 174 644 645 cell_1rw
* cell instance $10850 m0 *1 38.775,60.06
X$10850 175 43 176 644 645 cell_1rw
* cell instance $10851 m0 *1 39.48,60.06
X$10851 177 43 178 644 645 cell_1rw
* cell instance $10852 m0 *1 40.185,60.06
X$10852 179 43 180 644 645 cell_1rw
* cell instance $10853 m0 *1 40.89,60.06
X$10853 181 43 182 644 645 cell_1rw
* cell instance $10854 m0 *1 41.595,60.06
X$10854 183 43 184 644 645 cell_1rw
* cell instance $10855 m0 *1 42.3,60.06
X$10855 185 43 186 644 645 cell_1rw
* cell instance $10856 m0 *1 43.005,60.06
X$10856 187 43 188 644 645 cell_1rw
* cell instance $10857 m0 *1 43.71,60.06
X$10857 189 43 190 644 645 cell_1rw
* cell instance $10858 m0 *1 44.415,60.06
X$10858 191 43 192 644 645 cell_1rw
* cell instance $10859 m0 *1 45.12,60.06
X$10859 193 43 194 644 645 cell_1rw
* cell instance $10860 m0 *1 45.825,60.06
X$10860 195 43 196 644 645 cell_1rw
* cell instance $10861 m0 *1 46.53,60.06
X$10861 197 43 198 644 645 cell_1rw
* cell instance $10862 m0 *1 47.235,60.06
X$10862 199 43 200 644 645 cell_1rw
* cell instance $10863 m0 *1 47.94,60.06
X$10863 201 43 202 644 645 cell_1rw
* cell instance $10864 m0 *1 48.645,60.06
X$10864 203 43 204 644 645 cell_1rw
* cell instance $10865 m0 *1 49.35,60.06
X$10865 205 43 206 644 645 cell_1rw
* cell instance $10866 m0 *1 50.055,60.06
X$10866 207 43 208 644 645 cell_1rw
* cell instance $10867 m0 *1 50.76,60.06
X$10867 209 43 210 644 645 cell_1rw
* cell instance $10868 m0 *1 51.465,60.06
X$10868 211 43 212 644 645 cell_1rw
* cell instance $10869 m0 *1 52.17,60.06
X$10869 213 43 214 644 645 cell_1rw
* cell instance $10870 m0 *1 52.875,60.06
X$10870 215 43 216 644 645 cell_1rw
* cell instance $10871 m0 *1 53.58,60.06
X$10871 217 43 218 644 645 cell_1rw
* cell instance $10872 m0 *1 54.285,60.06
X$10872 219 43 220 644 645 cell_1rw
* cell instance $10873 m0 *1 54.99,60.06
X$10873 221 43 222 644 645 cell_1rw
* cell instance $10874 m0 *1 55.695,60.06
X$10874 223 43 224 644 645 cell_1rw
* cell instance $10875 m0 *1 56.4,60.06
X$10875 225 43 226 644 645 cell_1rw
* cell instance $10876 m0 *1 57.105,60.06
X$10876 227 43 228 644 645 cell_1rw
* cell instance $10877 m0 *1 57.81,60.06
X$10877 229 43 230 644 645 cell_1rw
* cell instance $10878 m0 *1 58.515,60.06
X$10878 231 43 232 644 645 cell_1rw
* cell instance $10879 m0 *1 59.22,60.06
X$10879 233 43 234 644 645 cell_1rw
* cell instance $10880 m0 *1 59.925,60.06
X$10880 235 43 236 644 645 cell_1rw
* cell instance $10881 m0 *1 60.63,60.06
X$10881 237 43 238 644 645 cell_1rw
* cell instance $10882 m0 *1 61.335,60.06
X$10882 239 43 240 644 645 cell_1rw
* cell instance $10883 m0 *1 62.04,60.06
X$10883 241 43 242 644 645 cell_1rw
* cell instance $10884 m0 *1 62.745,60.06
X$10884 243 43 244 644 645 cell_1rw
* cell instance $10885 m0 *1 63.45,60.06
X$10885 245 43 246 644 645 cell_1rw
* cell instance $10886 m0 *1 64.155,60.06
X$10886 247 43 248 644 645 cell_1rw
* cell instance $10887 m0 *1 64.86,60.06
X$10887 249 43 250 644 645 cell_1rw
* cell instance $10888 m0 *1 65.565,60.06
X$10888 251 43 252 644 645 cell_1rw
* cell instance $10889 m0 *1 66.27,60.06
X$10889 253 43 254 644 645 cell_1rw
* cell instance $10890 m0 *1 66.975,60.06
X$10890 255 43 256 644 645 cell_1rw
* cell instance $10891 m0 *1 67.68,60.06
X$10891 257 43 258 644 645 cell_1rw
* cell instance $10892 m0 *1 68.385,60.06
X$10892 259 43 260 644 645 cell_1rw
* cell instance $10893 m0 *1 69.09,60.06
X$10893 261 43 262 644 645 cell_1rw
* cell instance $10894 m0 *1 69.795,60.06
X$10894 263 43 264 644 645 cell_1rw
* cell instance $10895 m0 *1 70.5,60.06
X$10895 265 43 266 644 645 cell_1rw
* cell instance $10896 m0 *1 71.205,60.06
X$10896 267 43 268 644 645 cell_1rw
* cell instance $10897 m0 *1 71.91,60.06
X$10897 269 43 270 644 645 cell_1rw
* cell instance $10898 m0 *1 72.615,60.06
X$10898 271 43 272 644 645 cell_1rw
* cell instance $10899 m0 *1 73.32,60.06
X$10899 273 43 274 644 645 cell_1rw
* cell instance $10900 m0 *1 74.025,60.06
X$10900 275 43 276 644 645 cell_1rw
* cell instance $10901 m0 *1 74.73,60.06
X$10901 277 43 278 644 645 cell_1rw
* cell instance $10902 m0 *1 75.435,60.06
X$10902 279 43 280 644 645 cell_1rw
* cell instance $10903 m0 *1 76.14,60.06
X$10903 281 43 282 644 645 cell_1rw
* cell instance $10904 m0 *1 76.845,60.06
X$10904 283 43 284 644 645 cell_1rw
* cell instance $10905 m0 *1 77.55,60.06
X$10905 285 43 286 644 645 cell_1rw
* cell instance $10906 m0 *1 78.255,60.06
X$10906 287 43 288 644 645 cell_1rw
* cell instance $10907 m0 *1 78.96,60.06
X$10907 289 43 290 644 645 cell_1rw
* cell instance $10908 m0 *1 79.665,60.06
X$10908 291 43 292 644 645 cell_1rw
* cell instance $10909 m0 *1 80.37,60.06
X$10909 293 43 294 644 645 cell_1rw
* cell instance $10910 m0 *1 81.075,60.06
X$10910 295 43 296 644 645 cell_1rw
* cell instance $10911 m0 *1 81.78,60.06
X$10911 297 43 298 644 645 cell_1rw
* cell instance $10912 m0 *1 82.485,60.06
X$10912 299 43 300 644 645 cell_1rw
* cell instance $10913 m0 *1 83.19,60.06
X$10913 301 43 302 644 645 cell_1rw
* cell instance $10914 m0 *1 83.895,60.06
X$10914 303 43 304 644 645 cell_1rw
* cell instance $10915 m0 *1 84.6,60.06
X$10915 305 43 306 644 645 cell_1rw
* cell instance $10916 m0 *1 85.305,60.06
X$10916 307 43 308 644 645 cell_1rw
* cell instance $10917 m0 *1 86.01,60.06
X$10917 309 43 310 644 645 cell_1rw
* cell instance $10918 m0 *1 86.715,60.06
X$10918 311 43 312 644 645 cell_1rw
* cell instance $10919 m0 *1 87.42,60.06
X$10919 313 43 314 644 645 cell_1rw
* cell instance $10920 m0 *1 88.125,60.06
X$10920 315 43 316 644 645 cell_1rw
* cell instance $10921 m0 *1 88.83,60.06
X$10921 317 43 318 644 645 cell_1rw
* cell instance $10922 m0 *1 89.535,60.06
X$10922 319 43 320 644 645 cell_1rw
* cell instance $10923 m0 *1 90.24,60.06
X$10923 321 43 323 644 645 cell_1rw
* cell instance $10924 m0 *1 90.945,60.06
X$10924 324 43 325 644 645 cell_1rw
* cell instance $10925 m0 *1 91.65,60.06
X$10925 326 43 327 644 645 cell_1rw
* cell instance $10926 m0 *1 92.355,60.06
X$10926 328 43 329 644 645 cell_1rw
* cell instance $10927 m0 *1 93.06,60.06
X$10927 330 43 331 644 645 cell_1rw
* cell instance $10928 m0 *1 93.765,60.06
X$10928 332 43 333 644 645 cell_1rw
* cell instance $10929 m0 *1 94.47,60.06
X$10929 334 43 335 644 645 cell_1rw
* cell instance $10930 m0 *1 95.175,60.06
X$10930 336 43 337 644 645 cell_1rw
* cell instance $10931 m0 *1 95.88,60.06
X$10931 338 43 339 644 645 cell_1rw
* cell instance $10932 m0 *1 96.585,60.06
X$10932 340 43 341 644 645 cell_1rw
* cell instance $10933 m0 *1 97.29,60.06
X$10933 342 43 343 644 645 cell_1rw
* cell instance $10934 m0 *1 97.995,60.06
X$10934 344 43 345 644 645 cell_1rw
* cell instance $10935 m0 *1 98.7,60.06
X$10935 346 43 347 644 645 cell_1rw
* cell instance $10936 m0 *1 99.405,60.06
X$10936 348 43 349 644 645 cell_1rw
* cell instance $10937 m0 *1 100.11,60.06
X$10937 350 43 351 644 645 cell_1rw
* cell instance $10938 m0 *1 100.815,60.06
X$10938 352 43 353 644 645 cell_1rw
* cell instance $10939 m0 *1 101.52,60.06
X$10939 354 43 355 644 645 cell_1rw
* cell instance $10940 m0 *1 102.225,60.06
X$10940 356 43 357 644 645 cell_1rw
* cell instance $10941 m0 *1 102.93,60.06
X$10941 358 43 359 644 645 cell_1rw
* cell instance $10942 m0 *1 103.635,60.06
X$10942 360 43 361 644 645 cell_1rw
* cell instance $10943 m0 *1 104.34,60.06
X$10943 362 43 363 644 645 cell_1rw
* cell instance $10944 m0 *1 105.045,60.06
X$10944 364 43 365 644 645 cell_1rw
* cell instance $10945 m0 *1 105.75,60.06
X$10945 366 43 367 644 645 cell_1rw
* cell instance $10946 m0 *1 106.455,60.06
X$10946 368 43 369 644 645 cell_1rw
* cell instance $10947 m0 *1 107.16,60.06
X$10947 370 43 371 644 645 cell_1rw
* cell instance $10948 m0 *1 107.865,60.06
X$10948 372 43 373 644 645 cell_1rw
* cell instance $10949 m0 *1 108.57,60.06
X$10949 374 43 375 644 645 cell_1rw
* cell instance $10950 m0 *1 109.275,60.06
X$10950 376 43 377 644 645 cell_1rw
* cell instance $10951 m0 *1 109.98,60.06
X$10951 378 43 379 644 645 cell_1rw
* cell instance $10952 m0 *1 110.685,60.06
X$10952 380 43 381 644 645 cell_1rw
* cell instance $10953 m0 *1 111.39,60.06
X$10953 382 43 383 644 645 cell_1rw
* cell instance $10954 m0 *1 112.095,60.06
X$10954 384 43 385 644 645 cell_1rw
* cell instance $10955 m0 *1 112.8,60.06
X$10955 386 43 387 644 645 cell_1rw
* cell instance $10956 m0 *1 113.505,60.06
X$10956 388 43 389 644 645 cell_1rw
* cell instance $10957 m0 *1 114.21,60.06
X$10957 390 43 391 644 645 cell_1rw
* cell instance $10958 m0 *1 114.915,60.06
X$10958 392 43 393 644 645 cell_1rw
* cell instance $10959 m0 *1 115.62,60.06
X$10959 394 43 395 644 645 cell_1rw
* cell instance $10960 m0 *1 116.325,60.06
X$10960 396 43 397 644 645 cell_1rw
* cell instance $10961 m0 *1 117.03,60.06
X$10961 398 43 399 644 645 cell_1rw
* cell instance $10962 m0 *1 117.735,60.06
X$10962 400 43 401 644 645 cell_1rw
* cell instance $10963 m0 *1 118.44,60.06
X$10963 402 43 403 644 645 cell_1rw
* cell instance $10964 m0 *1 119.145,60.06
X$10964 404 43 405 644 645 cell_1rw
* cell instance $10965 m0 *1 119.85,60.06
X$10965 406 43 407 644 645 cell_1rw
* cell instance $10966 m0 *1 120.555,60.06
X$10966 408 43 409 644 645 cell_1rw
* cell instance $10967 m0 *1 121.26,60.06
X$10967 410 43 411 644 645 cell_1rw
* cell instance $10968 m0 *1 121.965,60.06
X$10968 412 43 413 644 645 cell_1rw
* cell instance $10969 m0 *1 122.67,60.06
X$10969 414 43 415 644 645 cell_1rw
* cell instance $10970 m0 *1 123.375,60.06
X$10970 416 43 417 644 645 cell_1rw
* cell instance $10971 m0 *1 124.08,60.06
X$10971 418 43 419 644 645 cell_1rw
* cell instance $10972 m0 *1 124.785,60.06
X$10972 420 43 421 644 645 cell_1rw
* cell instance $10973 m0 *1 125.49,60.06
X$10973 422 43 423 644 645 cell_1rw
* cell instance $10974 m0 *1 126.195,60.06
X$10974 424 43 425 644 645 cell_1rw
* cell instance $10975 m0 *1 126.9,60.06
X$10975 426 43 427 644 645 cell_1rw
* cell instance $10976 m0 *1 127.605,60.06
X$10976 428 43 429 644 645 cell_1rw
* cell instance $10977 m0 *1 128.31,60.06
X$10977 430 43 431 644 645 cell_1rw
* cell instance $10978 m0 *1 129.015,60.06
X$10978 432 43 433 644 645 cell_1rw
* cell instance $10979 m0 *1 129.72,60.06
X$10979 434 43 435 644 645 cell_1rw
* cell instance $10980 m0 *1 130.425,60.06
X$10980 436 43 437 644 645 cell_1rw
* cell instance $10981 m0 *1 131.13,60.06
X$10981 438 43 439 644 645 cell_1rw
* cell instance $10982 m0 *1 131.835,60.06
X$10982 440 43 441 644 645 cell_1rw
* cell instance $10983 m0 *1 132.54,60.06
X$10983 442 43 443 644 645 cell_1rw
* cell instance $10984 m0 *1 133.245,60.06
X$10984 444 43 445 644 645 cell_1rw
* cell instance $10985 m0 *1 133.95,60.06
X$10985 446 43 447 644 645 cell_1rw
* cell instance $10986 m0 *1 134.655,60.06
X$10986 448 43 449 644 645 cell_1rw
* cell instance $10987 m0 *1 135.36,60.06
X$10987 450 43 451 644 645 cell_1rw
* cell instance $10988 m0 *1 136.065,60.06
X$10988 452 43 453 644 645 cell_1rw
* cell instance $10989 m0 *1 136.77,60.06
X$10989 454 43 455 644 645 cell_1rw
* cell instance $10990 m0 *1 137.475,60.06
X$10990 456 43 457 644 645 cell_1rw
* cell instance $10991 m0 *1 138.18,60.06
X$10991 458 43 459 644 645 cell_1rw
* cell instance $10992 m0 *1 138.885,60.06
X$10992 460 43 461 644 645 cell_1rw
* cell instance $10993 m0 *1 139.59,60.06
X$10993 462 43 463 644 645 cell_1rw
* cell instance $10994 m0 *1 140.295,60.06
X$10994 464 43 465 644 645 cell_1rw
* cell instance $10995 m0 *1 141,60.06
X$10995 466 43 467 644 645 cell_1rw
* cell instance $10996 m0 *1 141.705,60.06
X$10996 468 43 469 644 645 cell_1rw
* cell instance $10997 m0 *1 142.41,60.06
X$10997 470 43 471 644 645 cell_1rw
* cell instance $10998 m0 *1 143.115,60.06
X$10998 472 43 473 644 645 cell_1rw
* cell instance $10999 m0 *1 143.82,60.06
X$10999 474 43 475 644 645 cell_1rw
* cell instance $11000 m0 *1 144.525,60.06
X$11000 476 43 477 644 645 cell_1rw
* cell instance $11001 m0 *1 145.23,60.06
X$11001 478 43 479 644 645 cell_1rw
* cell instance $11002 m0 *1 145.935,60.06
X$11002 480 43 481 644 645 cell_1rw
* cell instance $11003 m0 *1 146.64,60.06
X$11003 482 43 483 644 645 cell_1rw
* cell instance $11004 m0 *1 147.345,60.06
X$11004 484 43 485 644 645 cell_1rw
* cell instance $11005 m0 *1 148.05,60.06
X$11005 486 43 487 644 645 cell_1rw
* cell instance $11006 m0 *1 148.755,60.06
X$11006 488 43 489 644 645 cell_1rw
* cell instance $11007 m0 *1 149.46,60.06
X$11007 490 43 491 644 645 cell_1rw
* cell instance $11008 m0 *1 150.165,60.06
X$11008 492 43 493 644 645 cell_1rw
* cell instance $11009 m0 *1 150.87,60.06
X$11009 494 43 495 644 645 cell_1rw
* cell instance $11010 m0 *1 151.575,60.06
X$11010 496 43 497 644 645 cell_1rw
* cell instance $11011 m0 *1 152.28,60.06
X$11011 498 43 499 644 645 cell_1rw
* cell instance $11012 m0 *1 152.985,60.06
X$11012 500 43 501 644 645 cell_1rw
* cell instance $11013 m0 *1 153.69,60.06
X$11013 502 43 503 644 645 cell_1rw
* cell instance $11014 m0 *1 154.395,60.06
X$11014 504 43 505 644 645 cell_1rw
* cell instance $11015 m0 *1 155.1,60.06
X$11015 506 43 507 644 645 cell_1rw
* cell instance $11016 m0 *1 155.805,60.06
X$11016 508 43 509 644 645 cell_1rw
* cell instance $11017 m0 *1 156.51,60.06
X$11017 510 43 511 644 645 cell_1rw
* cell instance $11018 m0 *1 157.215,60.06
X$11018 512 43 513 644 645 cell_1rw
* cell instance $11019 m0 *1 157.92,60.06
X$11019 514 43 515 644 645 cell_1rw
* cell instance $11020 m0 *1 158.625,60.06
X$11020 516 43 517 644 645 cell_1rw
* cell instance $11021 m0 *1 159.33,60.06
X$11021 518 43 519 644 645 cell_1rw
* cell instance $11022 m0 *1 160.035,60.06
X$11022 520 43 521 644 645 cell_1rw
* cell instance $11023 m0 *1 160.74,60.06
X$11023 522 43 523 644 645 cell_1rw
* cell instance $11024 m0 *1 161.445,60.06
X$11024 524 43 525 644 645 cell_1rw
* cell instance $11025 m0 *1 162.15,60.06
X$11025 526 43 527 644 645 cell_1rw
* cell instance $11026 m0 *1 162.855,60.06
X$11026 528 43 529 644 645 cell_1rw
* cell instance $11027 m0 *1 163.56,60.06
X$11027 530 43 531 644 645 cell_1rw
* cell instance $11028 m0 *1 164.265,60.06
X$11028 532 43 533 644 645 cell_1rw
* cell instance $11029 m0 *1 164.97,60.06
X$11029 534 43 535 644 645 cell_1rw
* cell instance $11030 m0 *1 165.675,60.06
X$11030 536 43 537 644 645 cell_1rw
* cell instance $11031 m0 *1 166.38,60.06
X$11031 538 43 539 644 645 cell_1rw
* cell instance $11032 m0 *1 167.085,60.06
X$11032 540 43 541 644 645 cell_1rw
* cell instance $11033 m0 *1 167.79,60.06
X$11033 542 43 543 644 645 cell_1rw
* cell instance $11034 m0 *1 168.495,60.06
X$11034 544 43 545 644 645 cell_1rw
* cell instance $11035 m0 *1 169.2,60.06
X$11035 546 43 547 644 645 cell_1rw
* cell instance $11036 m0 *1 169.905,60.06
X$11036 548 43 549 644 645 cell_1rw
* cell instance $11037 m0 *1 170.61,60.06
X$11037 550 43 551 644 645 cell_1rw
* cell instance $11038 m0 *1 171.315,60.06
X$11038 552 43 553 644 645 cell_1rw
* cell instance $11039 m0 *1 172.02,60.06
X$11039 554 43 555 644 645 cell_1rw
* cell instance $11040 m0 *1 172.725,60.06
X$11040 556 43 557 644 645 cell_1rw
* cell instance $11041 m0 *1 173.43,60.06
X$11041 558 43 559 644 645 cell_1rw
* cell instance $11042 m0 *1 174.135,60.06
X$11042 560 43 561 644 645 cell_1rw
* cell instance $11043 m0 *1 174.84,60.06
X$11043 562 43 563 644 645 cell_1rw
* cell instance $11044 m0 *1 175.545,60.06
X$11044 564 43 565 644 645 cell_1rw
* cell instance $11045 m0 *1 176.25,60.06
X$11045 566 43 567 644 645 cell_1rw
* cell instance $11046 m0 *1 176.955,60.06
X$11046 568 43 569 644 645 cell_1rw
* cell instance $11047 m0 *1 177.66,60.06
X$11047 570 43 571 644 645 cell_1rw
* cell instance $11048 m0 *1 178.365,60.06
X$11048 572 43 573 644 645 cell_1rw
* cell instance $11049 m0 *1 179.07,60.06
X$11049 574 43 575 644 645 cell_1rw
* cell instance $11050 m0 *1 179.775,60.06
X$11050 576 43 577 644 645 cell_1rw
* cell instance $11051 m0 *1 180.48,60.06
X$11051 578 43 579 644 645 cell_1rw
* cell instance $11052 r0 *1 0.705,57.33
X$11052 67 44 68 644 645 cell_1rw
* cell instance $11053 r0 *1 0,57.33
X$11053 65 44 66 644 645 cell_1rw
* cell instance $11054 r0 *1 1.41,57.33
X$11054 69 44 70 644 645 cell_1rw
* cell instance $11055 r0 *1 2.115,57.33
X$11055 71 44 72 644 645 cell_1rw
* cell instance $11056 r0 *1 2.82,57.33
X$11056 73 44 74 644 645 cell_1rw
* cell instance $11057 r0 *1 3.525,57.33
X$11057 75 44 76 644 645 cell_1rw
* cell instance $11058 r0 *1 4.23,57.33
X$11058 77 44 78 644 645 cell_1rw
* cell instance $11059 r0 *1 4.935,57.33
X$11059 79 44 80 644 645 cell_1rw
* cell instance $11060 r0 *1 5.64,57.33
X$11060 81 44 82 644 645 cell_1rw
* cell instance $11061 r0 *1 6.345,57.33
X$11061 83 44 84 644 645 cell_1rw
* cell instance $11062 r0 *1 7.05,57.33
X$11062 85 44 86 644 645 cell_1rw
* cell instance $11063 r0 *1 7.755,57.33
X$11063 87 44 88 644 645 cell_1rw
* cell instance $11064 r0 *1 8.46,57.33
X$11064 89 44 90 644 645 cell_1rw
* cell instance $11065 r0 *1 9.165,57.33
X$11065 91 44 92 644 645 cell_1rw
* cell instance $11066 r0 *1 9.87,57.33
X$11066 93 44 94 644 645 cell_1rw
* cell instance $11067 r0 *1 10.575,57.33
X$11067 95 44 96 644 645 cell_1rw
* cell instance $11068 r0 *1 11.28,57.33
X$11068 97 44 98 644 645 cell_1rw
* cell instance $11069 r0 *1 11.985,57.33
X$11069 99 44 100 644 645 cell_1rw
* cell instance $11070 r0 *1 12.69,57.33
X$11070 101 44 102 644 645 cell_1rw
* cell instance $11071 r0 *1 13.395,57.33
X$11071 103 44 104 644 645 cell_1rw
* cell instance $11072 r0 *1 14.1,57.33
X$11072 105 44 106 644 645 cell_1rw
* cell instance $11073 r0 *1 14.805,57.33
X$11073 107 44 108 644 645 cell_1rw
* cell instance $11074 r0 *1 15.51,57.33
X$11074 109 44 110 644 645 cell_1rw
* cell instance $11075 r0 *1 16.215,57.33
X$11075 111 44 112 644 645 cell_1rw
* cell instance $11076 r0 *1 16.92,57.33
X$11076 113 44 114 644 645 cell_1rw
* cell instance $11077 r0 *1 17.625,57.33
X$11077 115 44 116 644 645 cell_1rw
* cell instance $11078 r0 *1 18.33,57.33
X$11078 117 44 118 644 645 cell_1rw
* cell instance $11079 r0 *1 19.035,57.33
X$11079 119 44 120 644 645 cell_1rw
* cell instance $11080 r0 *1 19.74,57.33
X$11080 121 44 122 644 645 cell_1rw
* cell instance $11081 r0 *1 20.445,57.33
X$11081 123 44 124 644 645 cell_1rw
* cell instance $11082 r0 *1 21.15,57.33
X$11082 125 44 126 644 645 cell_1rw
* cell instance $11083 r0 *1 21.855,57.33
X$11083 127 44 128 644 645 cell_1rw
* cell instance $11084 r0 *1 22.56,57.33
X$11084 129 44 130 644 645 cell_1rw
* cell instance $11085 r0 *1 23.265,57.33
X$11085 131 44 132 644 645 cell_1rw
* cell instance $11086 r0 *1 23.97,57.33
X$11086 133 44 134 644 645 cell_1rw
* cell instance $11087 r0 *1 24.675,57.33
X$11087 135 44 136 644 645 cell_1rw
* cell instance $11088 r0 *1 25.38,57.33
X$11088 137 44 138 644 645 cell_1rw
* cell instance $11089 r0 *1 26.085,57.33
X$11089 139 44 140 644 645 cell_1rw
* cell instance $11090 r0 *1 26.79,57.33
X$11090 141 44 142 644 645 cell_1rw
* cell instance $11091 r0 *1 27.495,57.33
X$11091 143 44 144 644 645 cell_1rw
* cell instance $11092 r0 *1 28.2,57.33
X$11092 145 44 146 644 645 cell_1rw
* cell instance $11093 r0 *1 28.905,57.33
X$11093 147 44 148 644 645 cell_1rw
* cell instance $11094 r0 *1 29.61,57.33
X$11094 149 44 150 644 645 cell_1rw
* cell instance $11095 r0 *1 30.315,57.33
X$11095 151 44 152 644 645 cell_1rw
* cell instance $11096 r0 *1 31.02,57.33
X$11096 153 44 154 644 645 cell_1rw
* cell instance $11097 r0 *1 31.725,57.33
X$11097 155 44 156 644 645 cell_1rw
* cell instance $11098 r0 *1 32.43,57.33
X$11098 157 44 158 644 645 cell_1rw
* cell instance $11099 r0 *1 33.135,57.33
X$11099 159 44 160 644 645 cell_1rw
* cell instance $11100 r0 *1 33.84,57.33
X$11100 161 44 162 644 645 cell_1rw
* cell instance $11101 r0 *1 34.545,57.33
X$11101 163 44 164 644 645 cell_1rw
* cell instance $11102 r0 *1 35.25,57.33
X$11102 165 44 166 644 645 cell_1rw
* cell instance $11103 r0 *1 35.955,57.33
X$11103 167 44 168 644 645 cell_1rw
* cell instance $11104 r0 *1 36.66,57.33
X$11104 169 44 170 644 645 cell_1rw
* cell instance $11105 r0 *1 37.365,57.33
X$11105 171 44 172 644 645 cell_1rw
* cell instance $11106 r0 *1 38.07,57.33
X$11106 173 44 174 644 645 cell_1rw
* cell instance $11107 r0 *1 38.775,57.33
X$11107 175 44 176 644 645 cell_1rw
* cell instance $11108 r0 *1 39.48,57.33
X$11108 177 44 178 644 645 cell_1rw
* cell instance $11109 r0 *1 40.185,57.33
X$11109 179 44 180 644 645 cell_1rw
* cell instance $11110 r0 *1 40.89,57.33
X$11110 181 44 182 644 645 cell_1rw
* cell instance $11111 r0 *1 41.595,57.33
X$11111 183 44 184 644 645 cell_1rw
* cell instance $11112 r0 *1 42.3,57.33
X$11112 185 44 186 644 645 cell_1rw
* cell instance $11113 r0 *1 43.005,57.33
X$11113 187 44 188 644 645 cell_1rw
* cell instance $11114 r0 *1 43.71,57.33
X$11114 189 44 190 644 645 cell_1rw
* cell instance $11115 r0 *1 44.415,57.33
X$11115 191 44 192 644 645 cell_1rw
* cell instance $11116 r0 *1 45.12,57.33
X$11116 193 44 194 644 645 cell_1rw
* cell instance $11117 r0 *1 45.825,57.33
X$11117 195 44 196 644 645 cell_1rw
* cell instance $11118 r0 *1 46.53,57.33
X$11118 197 44 198 644 645 cell_1rw
* cell instance $11119 r0 *1 47.235,57.33
X$11119 199 44 200 644 645 cell_1rw
* cell instance $11120 r0 *1 47.94,57.33
X$11120 201 44 202 644 645 cell_1rw
* cell instance $11121 r0 *1 48.645,57.33
X$11121 203 44 204 644 645 cell_1rw
* cell instance $11122 r0 *1 49.35,57.33
X$11122 205 44 206 644 645 cell_1rw
* cell instance $11123 r0 *1 50.055,57.33
X$11123 207 44 208 644 645 cell_1rw
* cell instance $11124 r0 *1 50.76,57.33
X$11124 209 44 210 644 645 cell_1rw
* cell instance $11125 r0 *1 51.465,57.33
X$11125 211 44 212 644 645 cell_1rw
* cell instance $11126 r0 *1 52.17,57.33
X$11126 213 44 214 644 645 cell_1rw
* cell instance $11127 r0 *1 52.875,57.33
X$11127 215 44 216 644 645 cell_1rw
* cell instance $11128 r0 *1 53.58,57.33
X$11128 217 44 218 644 645 cell_1rw
* cell instance $11129 r0 *1 54.285,57.33
X$11129 219 44 220 644 645 cell_1rw
* cell instance $11130 r0 *1 54.99,57.33
X$11130 221 44 222 644 645 cell_1rw
* cell instance $11131 r0 *1 55.695,57.33
X$11131 223 44 224 644 645 cell_1rw
* cell instance $11132 r0 *1 56.4,57.33
X$11132 225 44 226 644 645 cell_1rw
* cell instance $11133 r0 *1 57.105,57.33
X$11133 227 44 228 644 645 cell_1rw
* cell instance $11134 r0 *1 57.81,57.33
X$11134 229 44 230 644 645 cell_1rw
* cell instance $11135 r0 *1 58.515,57.33
X$11135 231 44 232 644 645 cell_1rw
* cell instance $11136 r0 *1 59.22,57.33
X$11136 233 44 234 644 645 cell_1rw
* cell instance $11137 r0 *1 59.925,57.33
X$11137 235 44 236 644 645 cell_1rw
* cell instance $11138 r0 *1 60.63,57.33
X$11138 237 44 238 644 645 cell_1rw
* cell instance $11139 r0 *1 61.335,57.33
X$11139 239 44 240 644 645 cell_1rw
* cell instance $11140 r0 *1 62.04,57.33
X$11140 241 44 242 644 645 cell_1rw
* cell instance $11141 r0 *1 62.745,57.33
X$11141 243 44 244 644 645 cell_1rw
* cell instance $11142 r0 *1 63.45,57.33
X$11142 245 44 246 644 645 cell_1rw
* cell instance $11143 r0 *1 64.155,57.33
X$11143 247 44 248 644 645 cell_1rw
* cell instance $11144 r0 *1 64.86,57.33
X$11144 249 44 250 644 645 cell_1rw
* cell instance $11145 r0 *1 65.565,57.33
X$11145 251 44 252 644 645 cell_1rw
* cell instance $11146 r0 *1 66.27,57.33
X$11146 253 44 254 644 645 cell_1rw
* cell instance $11147 r0 *1 66.975,57.33
X$11147 255 44 256 644 645 cell_1rw
* cell instance $11148 r0 *1 67.68,57.33
X$11148 257 44 258 644 645 cell_1rw
* cell instance $11149 r0 *1 68.385,57.33
X$11149 259 44 260 644 645 cell_1rw
* cell instance $11150 r0 *1 69.09,57.33
X$11150 261 44 262 644 645 cell_1rw
* cell instance $11151 r0 *1 69.795,57.33
X$11151 263 44 264 644 645 cell_1rw
* cell instance $11152 r0 *1 70.5,57.33
X$11152 265 44 266 644 645 cell_1rw
* cell instance $11153 r0 *1 71.205,57.33
X$11153 267 44 268 644 645 cell_1rw
* cell instance $11154 r0 *1 71.91,57.33
X$11154 269 44 270 644 645 cell_1rw
* cell instance $11155 r0 *1 72.615,57.33
X$11155 271 44 272 644 645 cell_1rw
* cell instance $11156 r0 *1 73.32,57.33
X$11156 273 44 274 644 645 cell_1rw
* cell instance $11157 r0 *1 74.025,57.33
X$11157 275 44 276 644 645 cell_1rw
* cell instance $11158 r0 *1 74.73,57.33
X$11158 277 44 278 644 645 cell_1rw
* cell instance $11159 r0 *1 75.435,57.33
X$11159 279 44 280 644 645 cell_1rw
* cell instance $11160 r0 *1 76.14,57.33
X$11160 281 44 282 644 645 cell_1rw
* cell instance $11161 r0 *1 76.845,57.33
X$11161 283 44 284 644 645 cell_1rw
* cell instance $11162 r0 *1 77.55,57.33
X$11162 285 44 286 644 645 cell_1rw
* cell instance $11163 r0 *1 78.255,57.33
X$11163 287 44 288 644 645 cell_1rw
* cell instance $11164 r0 *1 78.96,57.33
X$11164 289 44 290 644 645 cell_1rw
* cell instance $11165 r0 *1 79.665,57.33
X$11165 291 44 292 644 645 cell_1rw
* cell instance $11166 r0 *1 80.37,57.33
X$11166 293 44 294 644 645 cell_1rw
* cell instance $11167 r0 *1 81.075,57.33
X$11167 295 44 296 644 645 cell_1rw
* cell instance $11168 r0 *1 81.78,57.33
X$11168 297 44 298 644 645 cell_1rw
* cell instance $11169 r0 *1 82.485,57.33
X$11169 299 44 300 644 645 cell_1rw
* cell instance $11170 r0 *1 83.19,57.33
X$11170 301 44 302 644 645 cell_1rw
* cell instance $11171 r0 *1 83.895,57.33
X$11171 303 44 304 644 645 cell_1rw
* cell instance $11172 r0 *1 84.6,57.33
X$11172 305 44 306 644 645 cell_1rw
* cell instance $11173 r0 *1 85.305,57.33
X$11173 307 44 308 644 645 cell_1rw
* cell instance $11174 r0 *1 86.01,57.33
X$11174 309 44 310 644 645 cell_1rw
* cell instance $11175 r0 *1 86.715,57.33
X$11175 311 44 312 644 645 cell_1rw
* cell instance $11176 r0 *1 87.42,57.33
X$11176 313 44 314 644 645 cell_1rw
* cell instance $11177 r0 *1 88.125,57.33
X$11177 315 44 316 644 645 cell_1rw
* cell instance $11178 r0 *1 88.83,57.33
X$11178 317 44 318 644 645 cell_1rw
* cell instance $11179 r0 *1 89.535,57.33
X$11179 319 44 320 644 645 cell_1rw
* cell instance $11180 r0 *1 90.24,57.33
X$11180 321 44 323 644 645 cell_1rw
* cell instance $11181 r0 *1 90.945,57.33
X$11181 324 44 325 644 645 cell_1rw
* cell instance $11182 r0 *1 91.65,57.33
X$11182 326 44 327 644 645 cell_1rw
* cell instance $11183 r0 *1 92.355,57.33
X$11183 328 44 329 644 645 cell_1rw
* cell instance $11184 r0 *1 93.06,57.33
X$11184 330 44 331 644 645 cell_1rw
* cell instance $11185 r0 *1 93.765,57.33
X$11185 332 44 333 644 645 cell_1rw
* cell instance $11186 r0 *1 94.47,57.33
X$11186 334 44 335 644 645 cell_1rw
* cell instance $11187 r0 *1 95.175,57.33
X$11187 336 44 337 644 645 cell_1rw
* cell instance $11188 r0 *1 95.88,57.33
X$11188 338 44 339 644 645 cell_1rw
* cell instance $11189 r0 *1 96.585,57.33
X$11189 340 44 341 644 645 cell_1rw
* cell instance $11190 r0 *1 97.29,57.33
X$11190 342 44 343 644 645 cell_1rw
* cell instance $11191 r0 *1 97.995,57.33
X$11191 344 44 345 644 645 cell_1rw
* cell instance $11192 r0 *1 98.7,57.33
X$11192 346 44 347 644 645 cell_1rw
* cell instance $11193 r0 *1 99.405,57.33
X$11193 348 44 349 644 645 cell_1rw
* cell instance $11194 r0 *1 100.11,57.33
X$11194 350 44 351 644 645 cell_1rw
* cell instance $11195 r0 *1 100.815,57.33
X$11195 352 44 353 644 645 cell_1rw
* cell instance $11196 r0 *1 101.52,57.33
X$11196 354 44 355 644 645 cell_1rw
* cell instance $11197 r0 *1 102.225,57.33
X$11197 356 44 357 644 645 cell_1rw
* cell instance $11198 r0 *1 102.93,57.33
X$11198 358 44 359 644 645 cell_1rw
* cell instance $11199 r0 *1 103.635,57.33
X$11199 360 44 361 644 645 cell_1rw
* cell instance $11200 r0 *1 104.34,57.33
X$11200 362 44 363 644 645 cell_1rw
* cell instance $11201 r0 *1 105.045,57.33
X$11201 364 44 365 644 645 cell_1rw
* cell instance $11202 r0 *1 105.75,57.33
X$11202 366 44 367 644 645 cell_1rw
* cell instance $11203 r0 *1 106.455,57.33
X$11203 368 44 369 644 645 cell_1rw
* cell instance $11204 r0 *1 107.16,57.33
X$11204 370 44 371 644 645 cell_1rw
* cell instance $11205 r0 *1 107.865,57.33
X$11205 372 44 373 644 645 cell_1rw
* cell instance $11206 r0 *1 108.57,57.33
X$11206 374 44 375 644 645 cell_1rw
* cell instance $11207 r0 *1 109.275,57.33
X$11207 376 44 377 644 645 cell_1rw
* cell instance $11208 r0 *1 109.98,57.33
X$11208 378 44 379 644 645 cell_1rw
* cell instance $11209 r0 *1 110.685,57.33
X$11209 380 44 381 644 645 cell_1rw
* cell instance $11210 r0 *1 111.39,57.33
X$11210 382 44 383 644 645 cell_1rw
* cell instance $11211 r0 *1 112.095,57.33
X$11211 384 44 385 644 645 cell_1rw
* cell instance $11212 r0 *1 112.8,57.33
X$11212 386 44 387 644 645 cell_1rw
* cell instance $11213 r0 *1 113.505,57.33
X$11213 388 44 389 644 645 cell_1rw
* cell instance $11214 r0 *1 114.21,57.33
X$11214 390 44 391 644 645 cell_1rw
* cell instance $11215 r0 *1 114.915,57.33
X$11215 392 44 393 644 645 cell_1rw
* cell instance $11216 r0 *1 115.62,57.33
X$11216 394 44 395 644 645 cell_1rw
* cell instance $11217 r0 *1 116.325,57.33
X$11217 396 44 397 644 645 cell_1rw
* cell instance $11218 r0 *1 117.03,57.33
X$11218 398 44 399 644 645 cell_1rw
* cell instance $11219 r0 *1 117.735,57.33
X$11219 400 44 401 644 645 cell_1rw
* cell instance $11220 r0 *1 118.44,57.33
X$11220 402 44 403 644 645 cell_1rw
* cell instance $11221 r0 *1 119.145,57.33
X$11221 404 44 405 644 645 cell_1rw
* cell instance $11222 r0 *1 119.85,57.33
X$11222 406 44 407 644 645 cell_1rw
* cell instance $11223 r0 *1 120.555,57.33
X$11223 408 44 409 644 645 cell_1rw
* cell instance $11224 r0 *1 121.26,57.33
X$11224 410 44 411 644 645 cell_1rw
* cell instance $11225 r0 *1 121.965,57.33
X$11225 412 44 413 644 645 cell_1rw
* cell instance $11226 r0 *1 122.67,57.33
X$11226 414 44 415 644 645 cell_1rw
* cell instance $11227 r0 *1 123.375,57.33
X$11227 416 44 417 644 645 cell_1rw
* cell instance $11228 r0 *1 124.08,57.33
X$11228 418 44 419 644 645 cell_1rw
* cell instance $11229 r0 *1 124.785,57.33
X$11229 420 44 421 644 645 cell_1rw
* cell instance $11230 r0 *1 125.49,57.33
X$11230 422 44 423 644 645 cell_1rw
* cell instance $11231 r0 *1 126.195,57.33
X$11231 424 44 425 644 645 cell_1rw
* cell instance $11232 r0 *1 126.9,57.33
X$11232 426 44 427 644 645 cell_1rw
* cell instance $11233 r0 *1 127.605,57.33
X$11233 428 44 429 644 645 cell_1rw
* cell instance $11234 r0 *1 128.31,57.33
X$11234 430 44 431 644 645 cell_1rw
* cell instance $11235 r0 *1 129.015,57.33
X$11235 432 44 433 644 645 cell_1rw
* cell instance $11236 r0 *1 129.72,57.33
X$11236 434 44 435 644 645 cell_1rw
* cell instance $11237 r0 *1 130.425,57.33
X$11237 436 44 437 644 645 cell_1rw
* cell instance $11238 r0 *1 131.13,57.33
X$11238 438 44 439 644 645 cell_1rw
* cell instance $11239 r0 *1 131.835,57.33
X$11239 440 44 441 644 645 cell_1rw
* cell instance $11240 r0 *1 132.54,57.33
X$11240 442 44 443 644 645 cell_1rw
* cell instance $11241 r0 *1 133.245,57.33
X$11241 444 44 445 644 645 cell_1rw
* cell instance $11242 r0 *1 133.95,57.33
X$11242 446 44 447 644 645 cell_1rw
* cell instance $11243 r0 *1 134.655,57.33
X$11243 448 44 449 644 645 cell_1rw
* cell instance $11244 r0 *1 135.36,57.33
X$11244 450 44 451 644 645 cell_1rw
* cell instance $11245 r0 *1 136.065,57.33
X$11245 452 44 453 644 645 cell_1rw
* cell instance $11246 r0 *1 136.77,57.33
X$11246 454 44 455 644 645 cell_1rw
* cell instance $11247 r0 *1 137.475,57.33
X$11247 456 44 457 644 645 cell_1rw
* cell instance $11248 r0 *1 138.18,57.33
X$11248 458 44 459 644 645 cell_1rw
* cell instance $11249 r0 *1 138.885,57.33
X$11249 460 44 461 644 645 cell_1rw
* cell instance $11250 r0 *1 139.59,57.33
X$11250 462 44 463 644 645 cell_1rw
* cell instance $11251 r0 *1 140.295,57.33
X$11251 464 44 465 644 645 cell_1rw
* cell instance $11252 r0 *1 141,57.33
X$11252 466 44 467 644 645 cell_1rw
* cell instance $11253 r0 *1 141.705,57.33
X$11253 468 44 469 644 645 cell_1rw
* cell instance $11254 r0 *1 142.41,57.33
X$11254 470 44 471 644 645 cell_1rw
* cell instance $11255 r0 *1 143.115,57.33
X$11255 472 44 473 644 645 cell_1rw
* cell instance $11256 r0 *1 143.82,57.33
X$11256 474 44 475 644 645 cell_1rw
* cell instance $11257 r0 *1 144.525,57.33
X$11257 476 44 477 644 645 cell_1rw
* cell instance $11258 r0 *1 145.23,57.33
X$11258 478 44 479 644 645 cell_1rw
* cell instance $11259 r0 *1 145.935,57.33
X$11259 480 44 481 644 645 cell_1rw
* cell instance $11260 r0 *1 146.64,57.33
X$11260 482 44 483 644 645 cell_1rw
* cell instance $11261 r0 *1 147.345,57.33
X$11261 484 44 485 644 645 cell_1rw
* cell instance $11262 r0 *1 148.05,57.33
X$11262 486 44 487 644 645 cell_1rw
* cell instance $11263 r0 *1 148.755,57.33
X$11263 488 44 489 644 645 cell_1rw
* cell instance $11264 r0 *1 149.46,57.33
X$11264 490 44 491 644 645 cell_1rw
* cell instance $11265 r0 *1 150.165,57.33
X$11265 492 44 493 644 645 cell_1rw
* cell instance $11266 r0 *1 150.87,57.33
X$11266 494 44 495 644 645 cell_1rw
* cell instance $11267 r0 *1 151.575,57.33
X$11267 496 44 497 644 645 cell_1rw
* cell instance $11268 r0 *1 152.28,57.33
X$11268 498 44 499 644 645 cell_1rw
* cell instance $11269 r0 *1 152.985,57.33
X$11269 500 44 501 644 645 cell_1rw
* cell instance $11270 r0 *1 153.69,57.33
X$11270 502 44 503 644 645 cell_1rw
* cell instance $11271 r0 *1 154.395,57.33
X$11271 504 44 505 644 645 cell_1rw
* cell instance $11272 r0 *1 155.1,57.33
X$11272 506 44 507 644 645 cell_1rw
* cell instance $11273 r0 *1 155.805,57.33
X$11273 508 44 509 644 645 cell_1rw
* cell instance $11274 r0 *1 156.51,57.33
X$11274 510 44 511 644 645 cell_1rw
* cell instance $11275 r0 *1 157.215,57.33
X$11275 512 44 513 644 645 cell_1rw
* cell instance $11276 r0 *1 157.92,57.33
X$11276 514 44 515 644 645 cell_1rw
* cell instance $11277 r0 *1 158.625,57.33
X$11277 516 44 517 644 645 cell_1rw
* cell instance $11278 r0 *1 159.33,57.33
X$11278 518 44 519 644 645 cell_1rw
* cell instance $11279 r0 *1 160.035,57.33
X$11279 520 44 521 644 645 cell_1rw
* cell instance $11280 r0 *1 160.74,57.33
X$11280 522 44 523 644 645 cell_1rw
* cell instance $11281 r0 *1 161.445,57.33
X$11281 524 44 525 644 645 cell_1rw
* cell instance $11282 r0 *1 162.15,57.33
X$11282 526 44 527 644 645 cell_1rw
* cell instance $11283 r0 *1 162.855,57.33
X$11283 528 44 529 644 645 cell_1rw
* cell instance $11284 r0 *1 163.56,57.33
X$11284 530 44 531 644 645 cell_1rw
* cell instance $11285 r0 *1 164.265,57.33
X$11285 532 44 533 644 645 cell_1rw
* cell instance $11286 r0 *1 164.97,57.33
X$11286 534 44 535 644 645 cell_1rw
* cell instance $11287 r0 *1 165.675,57.33
X$11287 536 44 537 644 645 cell_1rw
* cell instance $11288 r0 *1 166.38,57.33
X$11288 538 44 539 644 645 cell_1rw
* cell instance $11289 r0 *1 167.085,57.33
X$11289 540 44 541 644 645 cell_1rw
* cell instance $11290 r0 *1 167.79,57.33
X$11290 542 44 543 644 645 cell_1rw
* cell instance $11291 r0 *1 168.495,57.33
X$11291 544 44 545 644 645 cell_1rw
* cell instance $11292 r0 *1 169.2,57.33
X$11292 546 44 547 644 645 cell_1rw
* cell instance $11293 r0 *1 169.905,57.33
X$11293 548 44 549 644 645 cell_1rw
* cell instance $11294 r0 *1 170.61,57.33
X$11294 550 44 551 644 645 cell_1rw
* cell instance $11295 r0 *1 171.315,57.33
X$11295 552 44 553 644 645 cell_1rw
* cell instance $11296 r0 *1 172.02,57.33
X$11296 554 44 555 644 645 cell_1rw
* cell instance $11297 r0 *1 172.725,57.33
X$11297 556 44 557 644 645 cell_1rw
* cell instance $11298 r0 *1 173.43,57.33
X$11298 558 44 559 644 645 cell_1rw
* cell instance $11299 r0 *1 174.135,57.33
X$11299 560 44 561 644 645 cell_1rw
* cell instance $11300 r0 *1 174.84,57.33
X$11300 562 44 563 644 645 cell_1rw
* cell instance $11301 r0 *1 175.545,57.33
X$11301 564 44 565 644 645 cell_1rw
* cell instance $11302 r0 *1 176.25,57.33
X$11302 566 44 567 644 645 cell_1rw
* cell instance $11303 r0 *1 176.955,57.33
X$11303 568 44 569 644 645 cell_1rw
* cell instance $11304 r0 *1 177.66,57.33
X$11304 570 44 571 644 645 cell_1rw
* cell instance $11305 r0 *1 178.365,57.33
X$11305 572 44 573 644 645 cell_1rw
* cell instance $11306 r0 *1 179.07,57.33
X$11306 574 44 575 644 645 cell_1rw
* cell instance $11307 r0 *1 179.775,57.33
X$11307 576 44 577 644 645 cell_1rw
* cell instance $11308 r0 *1 180.48,57.33
X$11308 578 44 579 644 645 cell_1rw
* cell instance $11309 r0 *1 0.705,60.06
X$11309 67 45 68 644 645 cell_1rw
* cell instance $11310 r0 *1 0,60.06
X$11310 65 45 66 644 645 cell_1rw
* cell instance $11311 r0 *1 1.41,60.06
X$11311 69 45 70 644 645 cell_1rw
* cell instance $11312 r0 *1 2.115,60.06
X$11312 71 45 72 644 645 cell_1rw
* cell instance $11313 r0 *1 2.82,60.06
X$11313 73 45 74 644 645 cell_1rw
* cell instance $11314 r0 *1 3.525,60.06
X$11314 75 45 76 644 645 cell_1rw
* cell instance $11315 r0 *1 4.23,60.06
X$11315 77 45 78 644 645 cell_1rw
* cell instance $11316 r0 *1 4.935,60.06
X$11316 79 45 80 644 645 cell_1rw
* cell instance $11317 r0 *1 5.64,60.06
X$11317 81 45 82 644 645 cell_1rw
* cell instance $11318 r0 *1 6.345,60.06
X$11318 83 45 84 644 645 cell_1rw
* cell instance $11319 r0 *1 7.05,60.06
X$11319 85 45 86 644 645 cell_1rw
* cell instance $11320 r0 *1 7.755,60.06
X$11320 87 45 88 644 645 cell_1rw
* cell instance $11321 r0 *1 8.46,60.06
X$11321 89 45 90 644 645 cell_1rw
* cell instance $11322 r0 *1 9.165,60.06
X$11322 91 45 92 644 645 cell_1rw
* cell instance $11323 r0 *1 9.87,60.06
X$11323 93 45 94 644 645 cell_1rw
* cell instance $11324 r0 *1 10.575,60.06
X$11324 95 45 96 644 645 cell_1rw
* cell instance $11325 r0 *1 11.28,60.06
X$11325 97 45 98 644 645 cell_1rw
* cell instance $11326 r0 *1 11.985,60.06
X$11326 99 45 100 644 645 cell_1rw
* cell instance $11327 r0 *1 12.69,60.06
X$11327 101 45 102 644 645 cell_1rw
* cell instance $11328 r0 *1 13.395,60.06
X$11328 103 45 104 644 645 cell_1rw
* cell instance $11329 r0 *1 14.1,60.06
X$11329 105 45 106 644 645 cell_1rw
* cell instance $11330 r0 *1 14.805,60.06
X$11330 107 45 108 644 645 cell_1rw
* cell instance $11331 r0 *1 15.51,60.06
X$11331 109 45 110 644 645 cell_1rw
* cell instance $11332 r0 *1 16.215,60.06
X$11332 111 45 112 644 645 cell_1rw
* cell instance $11333 r0 *1 16.92,60.06
X$11333 113 45 114 644 645 cell_1rw
* cell instance $11334 r0 *1 17.625,60.06
X$11334 115 45 116 644 645 cell_1rw
* cell instance $11335 r0 *1 18.33,60.06
X$11335 117 45 118 644 645 cell_1rw
* cell instance $11336 r0 *1 19.035,60.06
X$11336 119 45 120 644 645 cell_1rw
* cell instance $11337 r0 *1 19.74,60.06
X$11337 121 45 122 644 645 cell_1rw
* cell instance $11338 r0 *1 20.445,60.06
X$11338 123 45 124 644 645 cell_1rw
* cell instance $11339 r0 *1 21.15,60.06
X$11339 125 45 126 644 645 cell_1rw
* cell instance $11340 r0 *1 21.855,60.06
X$11340 127 45 128 644 645 cell_1rw
* cell instance $11341 r0 *1 22.56,60.06
X$11341 129 45 130 644 645 cell_1rw
* cell instance $11342 r0 *1 23.265,60.06
X$11342 131 45 132 644 645 cell_1rw
* cell instance $11343 r0 *1 23.97,60.06
X$11343 133 45 134 644 645 cell_1rw
* cell instance $11344 r0 *1 24.675,60.06
X$11344 135 45 136 644 645 cell_1rw
* cell instance $11345 r0 *1 25.38,60.06
X$11345 137 45 138 644 645 cell_1rw
* cell instance $11346 r0 *1 26.085,60.06
X$11346 139 45 140 644 645 cell_1rw
* cell instance $11347 r0 *1 26.79,60.06
X$11347 141 45 142 644 645 cell_1rw
* cell instance $11348 r0 *1 27.495,60.06
X$11348 143 45 144 644 645 cell_1rw
* cell instance $11349 r0 *1 28.2,60.06
X$11349 145 45 146 644 645 cell_1rw
* cell instance $11350 r0 *1 28.905,60.06
X$11350 147 45 148 644 645 cell_1rw
* cell instance $11351 r0 *1 29.61,60.06
X$11351 149 45 150 644 645 cell_1rw
* cell instance $11352 r0 *1 30.315,60.06
X$11352 151 45 152 644 645 cell_1rw
* cell instance $11353 r0 *1 31.02,60.06
X$11353 153 45 154 644 645 cell_1rw
* cell instance $11354 r0 *1 31.725,60.06
X$11354 155 45 156 644 645 cell_1rw
* cell instance $11355 r0 *1 32.43,60.06
X$11355 157 45 158 644 645 cell_1rw
* cell instance $11356 r0 *1 33.135,60.06
X$11356 159 45 160 644 645 cell_1rw
* cell instance $11357 r0 *1 33.84,60.06
X$11357 161 45 162 644 645 cell_1rw
* cell instance $11358 r0 *1 34.545,60.06
X$11358 163 45 164 644 645 cell_1rw
* cell instance $11359 r0 *1 35.25,60.06
X$11359 165 45 166 644 645 cell_1rw
* cell instance $11360 r0 *1 35.955,60.06
X$11360 167 45 168 644 645 cell_1rw
* cell instance $11361 r0 *1 36.66,60.06
X$11361 169 45 170 644 645 cell_1rw
* cell instance $11362 r0 *1 37.365,60.06
X$11362 171 45 172 644 645 cell_1rw
* cell instance $11363 r0 *1 38.07,60.06
X$11363 173 45 174 644 645 cell_1rw
* cell instance $11364 r0 *1 38.775,60.06
X$11364 175 45 176 644 645 cell_1rw
* cell instance $11365 r0 *1 39.48,60.06
X$11365 177 45 178 644 645 cell_1rw
* cell instance $11366 r0 *1 40.185,60.06
X$11366 179 45 180 644 645 cell_1rw
* cell instance $11367 r0 *1 40.89,60.06
X$11367 181 45 182 644 645 cell_1rw
* cell instance $11368 r0 *1 41.595,60.06
X$11368 183 45 184 644 645 cell_1rw
* cell instance $11369 r0 *1 42.3,60.06
X$11369 185 45 186 644 645 cell_1rw
* cell instance $11370 r0 *1 43.005,60.06
X$11370 187 45 188 644 645 cell_1rw
* cell instance $11371 r0 *1 43.71,60.06
X$11371 189 45 190 644 645 cell_1rw
* cell instance $11372 r0 *1 44.415,60.06
X$11372 191 45 192 644 645 cell_1rw
* cell instance $11373 r0 *1 45.12,60.06
X$11373 193 45 194 644 645 cell_1rw
* cell instance $11374 r0 *1 45.825,60.06
X$11374 195 45 196 644 645 cell_1rw
* cell instance $11375 r0 *1 46.53,60.06
X$11375 197 45 198 644 645 cell_1rw
* cell instance $11376 r0 *1 47.235,60.06
X$11376 199 45 200 644 645 cell_1rw
* cell instance $11377 r0 *1 47.94,60.06
X$11377 201 45 202 644 645 cell_1rw
* cell instance $11378 r0 *1 48.645,60.06
X$11378 203 45 204 644 645 cell_1rw
* cell instance $11379 r0 *1 49.35,60.06
X$11379 205 45 206 644 645 cell_1rw
* cell instance $11380 r0 *1 50.055,60.06
X$11380 207 45 208 644 645 cell_1rw
* cell instance $11381 r0 *1 50.76,60.06
X$11381 209 45 210 644 645 cell_1rw
* cell instance $11382 r0 *1 51.465,60.06
X$11382 211 45 212 644 645 cell_1rw
* cell instance $11383 r0 *1 52.17,60.06
X$11383 213 45 214 644 645 cell_1rw
* cell instance $11384 r0 *1 52.875,60.06
X$11384 215 45 216 644 645 cell_1rw
* cell instance $11385 r0 *1 53.58,60.06
X$11385 217 45 218 644 645 cell_1rw
* cell instance $11386 r0 *1 54.285,60.06
X$11386 219 45 220 644 645 cell_1rw
* cell instance $11387 r0 *1 54.99,60.06
X$11387 221 45 222 644 645 cell_1rw
* cell instance $11388 r0 *1 55.695,60.06
X$11388 223 45 224 644 645 cell_1rw
* cell instance $11389 r0 *1 56.4,60.06
X$11389 225 45 226 644 645 cell_1rw
* cell instance $11390 r0 *1 57.105,60.06
X$11390 227 45 228 644 645 cell_1rw
* cell instance $11391 r0 *1 57.81,60.06
X$11391 229 45 230 644 645 cell_1rw
* cell instance $11392 r0 *1 58.515,60.06
X$11392 231 45 232 644 645 cell_1rw
* cell instance $11393 r0 *1 59.22,60.06
X$11393 233 45 234 644 645 cell_1rw
* cell instance $11394 r0 *1 59.925,60.06
X$11394 235 45 236 644 645 cell_1rw
* cell instance $11395 r0 *1 60.63,60.06
X$11395 237 45 238 644 645 cell_1rw
* cell instance $11396 r0 *1 61.335,60.06
X$11396 239 45 240 644 645 cell_1rw
* cell instance $11397 r0 *1 62.04,60.06
X$11397 241 45 242 644 645 cell_1rw
* cell instance $11398 r0 *1 62.745,60.06
X$11398 243 45 244 644 645 cell_1rw
* cell instance $11399 r0 *1 63.45,60.06
X$11399 245 45 246 644 645 cell_1rw
* cell instance $11400 r0 *1 64.155,60.06
X$11400 247 45 248 644 645 cell_1rw
* cell instance $11401 r0 *1 64.86,60.06
X$11401 249 45 250 644 645 cell_1rw
* cell instance $11402 r0 *1 65.565,60.06
X$11402 251 45 252 644 645 cell_1rw
* cell instance $11403 r0 *1 66.27,60.06
X$11403 253 45 254 644 645 cell_1rw
* cell instance $11404 r0 *1 66.975,60.06
X$11404 255 45 256 644 645 cell_1rw
* cell instance $11405 r0 *1 67.68,60.06
X$11405 257 45 258 644 645 cell_1rw
* cell instance $11406 r0 *1 68.385,60.06
X$11406 259 45 260 644 645 cell_1rw
* cell instance $11407 r0 *1 69.09,60.06
X$11407 261 45 262 644 645 cell_1rw
* cell instance $11408 r0 *1 69.795,60.06
X$11408 263 45 264 644 645 cell_1rw
* cell instance $11409 r0 *1 70.5,60.06
X$11409 265 45 266 644 645 cell_1rw
* cell instance $11410 r0 *1 71.205,60.06
X$11410 267 45 268 644 645 cell_1rw
* cell instance $11411 r0 *1 71.91,60.06
X$11411 269 45 270 644 645 cell_1rw
* cell instance $11412 r0 *1 72.615,60.06
X$11412 271 45 272 644 645 cell_1rw
* cell instance $11413 r0 *1 73.32,60.06
X$11413 273 45 274 644 645 cell_1rw
* cell instance $11414 r0 *1 74.025,60.06
X$11414 275 45 276 644 645 cell_1rw
* cell instance $11415 r0 *1 74.73,60.06
X$11415 277 45 278 644 645 cell_1rw
* cell instance $11416 r0 *1 75.435,60.06
X$11416 279 45 280 644 645 cell_1rw
* cell instance $11417 r0 *1 76.14,60.06
X$11417 281 45 282 644 645 cell_1rw
* cell instance $11418 r0 *1 76.845,60.06
X$11418 283 45 284 644 645 cell_1rw
* cell instance $11419 r0 *1 77.55,60.06
X$11419 285 45 286 644 645 cell_1rw
* cell instance $11420 r0 *1 78.255,60.06
X$11420 287 45 288 644 645 cell_1rw
* cell instance $11421 r0 *1 78.96,60.06
X$11421 289 45 290 644 645 cell_1rw
* cell instance $11422 r0 *1 79.665,60.06
X$11422 291 45 292 644 645 cell_1rw
* cell instance $11423 r0 *1 80.37,60.06
X$11423 293 45 294 644 645 cell_1rw
* cell instance $11424 r0 *1 81.075,60.06
X$11424 295 45 296 644 645 cell_1rw
* cell instance $11425 r0 *1 81.78,60.06
X$11425 297 45 298 644 645 cell_1rw
* cell instance $11426 r0 *1 82.485,60.06
X$11426 299 45 300 644 645 cell_1rw
* cell instance $11427 r0 *1 83.19,60.06
X$11427 301 45 302 644 645 cell_1rw
* cell instance $11428 r0 *1 83.895,60.06
X$11428 303 45 304 644 645 cell_1rw
* cell instance $11429 r0 *1 84.6,60.06
X$11429 305 45 306 644 645 cell_1rw
* cell instance $11430 r0 *1 85.305,60.06
X$11430 307 45 308 644 645 cell_1rw
* cell instance $11431 r0 *1 86.01,60.06
X$11431 309 45 310 644 645 cell_1rw
* cell instance $11432 r0 *1 86.715,60.06
X$11432 311 45 312 644 645 cell_1rw
* cell instance $11433 r0 *1 87.42,60.06
X$11433 313 45 314 644 645 cell_1rw
* cell instance $11434 r0 *1 88.125,60.06
X$11434 315 45 316 644 645 cell_1rw
* cell instance $11435 r0 *1 88.83,60.06
X$11435 317 45 318 644 645 cell_1rw
* cell instance $11436 r0 *1 89.535,60.06
X$11436 319 45 320 644 645 cell_1rw
* cell instance $11437 r0 *1 90.24,60.06
X$11437 321 45 323 644 645 cell_1rw
* cell instance $11438 r0 *1 90.945,60.06
X$11438 324 45 325 644 645 cell_1rw
* cell instance $11439 r0 *1 91.65,60.06
X$11439 326 45 327 644 645 cell_1rw
* cell instance $11440 r0 *1 92.355,60.06
X$11440 328 45 329 644 645 cell_1rw
* cell instance $11441 r0 *1 93.06,60.06
X$11441 330 45 331 644 645 cell_1rw
* cell instance $11442 r0 *1 93.765,60.06
X$11442 332 45 333 644 645 cell_1rw
* cell instance $11443 r0 *1 94.47,60.06
X$11443 334 45 335 644 645 cell_1rw
* cell instance $11444 r0 *1 95.175,60.06
X$11444 336 45 337 644 645 cell_1rw
* cell instance $11445 r0 *1 95.88,60.06
X$11445 338 45 339 644 645 cell_1rw
* cell instance $11446 r0 *1 96.585,60.06
X$11446 340 45 341 644 645 cell_1rw
* cell instance $11447 r0 *1 97.29,60.06
X$11447 342 45 343 644 645 cell_1rw
* cell instance $11448 r0 *1 97.995,60.06
X$11448 344 45 345 644 645 cell_1rw
* cell instance $11449 r0 *1 98.7,60.06
X$11449 346 45 347 644 645 cell_1rw
* cell instance $11450 r0 *1 99.405,60.06
X$11450 348 45 349 644 645 cell_1rw
* cell instance $11451 r0 *1 100.11,60.06
X$11451 350 45 351 644 645 cell_1rw
* cell instance $11452 r0 *1 100.815,60.06
X$11452 352 45 353 644 645 cell_1rw
* cell instance $11453 r0 *1 101.52,60.06
X$11453 354 45 355 644 645 cell_1rw
* cell instance $11454 r0 *1 102.225,60.06
X$11454 356 45 357 644 645 cell_1rw
* cell instance $11455 r0 *1 102.93,60.06
X$11455 358 45 359 644 645 cell_1rw
* cell instance $11456 r0 *1 103.635,60.06
X$11456 360 45 361 644 645 cell_1rw
* cell instance $11457 r0 *1 104.34,60.06
X$11457 362 45 363 644 645 cell_1rw
* cell instance $11458 r0 *1 105.045,60.06
X$11458 364 45 365 644 645 cell_1rw
* cell instance $11459 r0 *1 105.75,60.06
X$11459 366 45 367 644 645 cell_1rw
* cell instance $11460 r0 *1 106.455,60.06
X$11460 368 45 369 644 645 cell_1rw
* cell instance $11461 r0 *1 107.16,60.06
X$11461 370 45 371 644 645 cell_1rw
* cell instance $11462 r0 *1 107.865,60.06
X$11462 372 45 373 644 645 cell_1rw
* cell instance $11463 r0 *1 108.57,60.06
X$11463 374 45 375 644 645 cell_1rw
* cell instance $11464 r0 *1 109.275,60.06
X$11464 376 45 377 644 645 cell_1rw
* cell instance $11465 r0 *1 109.98,60.06
X$11465 378 45 379 644 645 cell_1rw
* cell instance $11466 r0 *1 110.685,60.06
X$11466 380 45 381 644 645 cell_1rw
* cell instance $11467 r0 *1 111.39,60.06
X$11467 382 45 383 644 645 cell_1rw
* cell instance $11468 r0 *1 112.095,60.06
X$11468 384 45 385 644 645 cell_1rw
* cell instance $11469 r0 *1 112.8,60.06
X$11469 386 45 387 644 645 cell_1rw
* cell instance $11470 r0 *1 113.505,60.06
X$11470 388 45 389 644 645 cell_1rw
* cell instance $11471 r0 *1 114.21,60.06
X$11471 390 45 391 644 645 cell_1rw
* cell instance $11472 r0 *1 114.915,60.06
X$11472 392 45 393 644 645 cell_1rw
* cell instance $11473 r0 *1 115.62,60.06
X$11473 394 45 395 644 645 cell_1rw
* cell instance $11474 r0 *1 116.325,60.06
X$11474 396 45 397 644 645 cell_1rw
* cell instance $11475 r0 *1 117.03,60.06
X$11475 398 45 399 644 645 cell_1rw
* cell instance $11476 r0 *1 117.735,60.06
X$11476 400 45 401 644 645 cell_1rw
* cell instance $11477 r0 *1 118.44,60.06
X$11477 402 45 403 644 645 cell_1rw
* cell instance $11478 r0 *1 119.145,60.06
X$11478 404 45 405 644 645 cell_1rw
* cell instance $11479 r0 *1 119.85,60.06
X$11479 406 45 407 644 645 cell_1rw
* cell instance $11480 r0 *1 120.555,60.06
X$11480 408 45 409 644 645 cell_1rw
* cell instance $11481 r0 *1 121.26,60.06
X$11481 410 45 411 644 645 cell_1rw
* cell instance $11482 r0 *1 121.965,60.06
X$11482 412 45 413 644 645 cell_1rw
* cell instance $11483 r0 *1 122.67,60.06
X$11483 414 45 415 644 645 cell_1rw
* cell instance $11484 r0 *1 123.375,60.06
X$11484 416 45 417 644 645 cell_1rw
* cell instance $11485 r0 *1 124.08,60.06
X$11485 418 45 419 644 645 cell_1rw
* cell instance $11486 r0 *1 124.785,60.06
X$11486 420 45 421 644 645 cell_1rw
* cell instance $11487 r0 *1 125.49,60.06
X$11487 422 45 423 644 645 cell_1rw
* cell instance $11488 r0 *1 126.195,60.06
X$11488 424 45 425 644 645 cell_1rw
* cell instance $11489 r0 *1 126.9,60.06
X$11489 426 45 427 644 645 cell_1rw
* cell instance $11490 r0 *1 127.605,60.06
X$11490 428 45 429 644 645 cell_1rw
* cell instance $11491 r0 *1 128.31,60.06
X$11491 430 45 431 644 645 cell_1rw
* cell instance $11492 r0 *1 129.015,60.06
X$11492 432 45 433 644 645 cell_1rw
* cell instance $11493 r0 *1 129.72,60.06
X$11493 434 45 435 644 645 cell_1rw
* cell instance $11494 r0 *1 130.425,60.06
X$11494 436 45 437 644 645 cell_1rw
* cell instance $11495 r0 *1 131.13,60.06
X$11495 438 45 439 644 645 cell_1rw
* cell instance $11496 r0 *1 131.835,60.06
X$11496 440 45 441 644 645 cell_1rw
* cell instance $11497 r0 *1 132.54,60.06
X$11497 442 45 443 644 645 cell_1rw
* cell instance $11498 r0 *1 133.245,60.06
X$11498 444 45 445 644 645 cell_1rw
* cell instance $11499 r0 *1 133.95,60.06
X$11499 446 45 447 644 645 cell_1rw
* cell instance $11500 r0 *1 134.655,60.06
X$11500 448 45 449 644 645 cell_1rw
* cell instance $11501 r0 *1 135.36,60.06
X$11501 450 45 451 644 645 cell_1rw
* cell instance $11502 r0 *1 136.065,60.06
X$11502 452 45 453 644 645 cell_1rw
* cell instance $11503 r0 *1 136.77,60.06
X$11503 454 45 455 644 645 cell_1rw
* cell instance $11504 r0 *1 137.475,60.06
X$11504 456 45 457 644 645 cell_1rw
* cell instance $11505 r0 *1 138.18,60.06
X$11505 458 45 459 644 645 cell_1rw
* cell instance $11506 r0 *1 138.885,60.06
X$11506 460 45 461 644 645 cell_1rw
* cell instance $11507 r0 *1 139.59,60.06
X$11507 462 45 463 644 645 cell_1rw
* cell instance $11508 r0 *1 140.295,60.06
X$11508 464 45 465 644 645 cell_1rw
* cell instance $11509 r0 *1 141,60.06
X$11509 466 45 467 644 645 cell_1rw
* cell instance $11510 r0 *1 141.705,60.06
X$11510 468 45 469 644 645 cell_1rw
* cell instance $11511 r0 *1 142.41,60.06
X$11511 470 45 471 644 645 cell_1rw
* cell instance $11512 r0 *1 143.115,60.06
X$11512 472 45 473 644 645 cell_1rw
* cell instance $11513 r0 *1 143.82,60.06
X$11513 474 45 475 644 645 cell_1rw
* cell instance $11514 r0 *1 144.525,60.06
X$11514 476 45 477 644 645 cell_1rw
* cell instance $11515 r0 *1 145.23,60.06
X$11515 478 45 479 644 645 cell_1rw
* cell instance $11516 r0 *1 145.935,60.06
X$11516 480 45 481 644 645 cell_1rw
* cell instance $11517 r0 *1 146.64,60.06
X$11517 482 45 483 644 645 cell_1rw
* cell instance $11518 r0 *1 147.345,60.06
X$11518 484 45 485 644 645 cell_1rw
* cell instance $11519 r0 *1 148.05,60.06
X$11519 486 45 487 644 645 cell_1rw
* cell instance $11520 r0 *1 148.755,60.06
X$11520 488 45 489 644 645 cell_1rw
* cell instance $11521 r0 *1 149.46,60.06
X$11521 490 45 491 644 645 cell_1rw
* cell instance $11522 r0 *1 150.165,60.06
X$11522 492 45 493 644 645 cell_1rw
* cell instance $11523 r0 *1 150.87,60.06
X$11523 494 45 495 644 645 cell_1rw
* cell instance $11524 r0 *1 151.575,60.06
X$11524 496 45 497 644 645 cell_1rw
* cell instance $11525 r0 *1 152.28,60.06
X$11525 498 45 499 644 645 cell_1rw
* cell instance $11526 r0 *1 152.985,60.06
X$11526 500 45 501 644 645 cell_1rw
* cell instance $11527 r0 *1 153.69,60.06
X$11527 502 45 503 644 645 cell_1rw
* cell instance $11528 r0 *1 154.395,60.06
X$11528 504 45 505 644 645 cell_1rw
* cell instance $11529 r0 *1 155.1,60.06
X$11529 506 45 507 644 645 cell_1rw
* cell instance $11530 r0 *1 155.805,60.06
X$11530 508 45 509 644 645 cell_1rw
* cell instance $11531 r0 *1 156.51,60.06
X$11531 510 45 511 644 645 cell_1rw
* cell instance $11532 r0 *1 157.215,60.06
X$11532 512 45 513 644 645 cell_1rw
* cell instance $11533 r0 *1 157.92,60.06
X$11533 514 45 515 644 645 cell_1rw
* cell instance $11534 r0 *1 158.625,60.06
X$11534 516 45 517 644 645 cell_1rw
* cell instance $11535 r0 *1 159.33,60.06
X$11535 518 45 519 644 645 cell_1rw
* cell instance $11536 r0 *1 160.035,60.06
X$11536 520 45 521 644 645 cell_1rw
* cell instance $11537 r0 *1 160.74,60.06
X$11537 522 45 523 644 645 cell_1rw
* cell instance $11538 r0 *1 161.445,60.06
X$11538 524 45 525 644 645 cell_1rw
* cell instance $11539 r0 *1 162.15,60.06
X$11539 526 45 527 644 645 cell_1rw
* cell instance $11540 r0 *1 162.855,60.06
X$11540 528 45 529 644 645 cell_1rw
* cell instance $11541 r0 *1 163.56,60.06
X$11541 530 45 531 644 645 cell_1rw
* cell instance $11542 r0 *1 164.265,60.06
X$11542 532 45 533 644 645 cell_1rw
* cell instance $11543 r0 *1 164.97,60.06
X$11543 534 45 535 644 645 cell_1rw
* cell instance $11544 r0 *1 165.675,60.06
X$11544 536 45 537 644 645 cell_1rw
* cell instance $11545 r0 *1 166.38,60.06
X$11545 538 45 539 644 645 cell_1rw
* cell instance $11546 r0 *1 167.085,60.06
X$11546 540 45 541 644 645 cell_1rw
* cell instance $11547 r0 *1 167.79,60.06
X$11547 542 45 543 644 645 cell_1rw
* cell instance $11548 r0 *1 168.495,60.06
X$11548 544 45 545 644 645 cell_1rw
* cell instance $11549 r0 *1 169.2,60.06
X$11549 546 45 547 644 645 cell_1rw
* cell instance $11550 r0 *1 169.905,60.06
X$11550 548 45 549 644 645 cell_1rw
* cell instance $11551 r0 *1 170.61,60.06
X$11551 550 45 551 644 645 cell_1rw
* cell instance $11552 r0 *1 171.315,60.06
X$11552 552 45 553 644 645 cell_1rw
* cell instance $11553 r0 *1 172.02,60.06
X$11553 554 45 555 644 645 cell_1rw
* cell instance $11554 r0 *1 172.725,60.06
X$11554 556 45 557 644 645 cell_1rw
* cell instance $11555 r0 *1 173.43,60.06
X$11555 558 45 559 644 645 cell_1rw
* cell instance $11556 r0 *1 174.135,60.06
X$11556 560 45 561 644 645 cell_1rw
* cell instance $11557 r0 *1 174.84,60.06
X$11557 562 45 563 644 645 cell_1rw
* cell instance $11558 r0 *1 175.545,60.06
X$11558 564 45 565 644 645 cell_1rw
* cell instance $11559 r0 *1 176.25,60.06
X$11559 566 45 567 644 645 cell_1rw
* cell instance $11560 r0 *1 176.955,60.06
X$11560 568 45 569 644 645 cell_1rw
* cell instance $11561 r0 *1 177.66,60.06
X$11561 570 45 571 644 645 cell_1rw
* cell instance $11562 r0 *1 178.365,60.06
X$11562 572 45 573 644 645 cell_1rw
* cell instance $11563 r0 *1 179.07,60.06
X$11563 574 45 575 644 645 cell_1rw
* cell instance $11564 r0 *1 179.775,60.06
X$11564 576 45 577 644 645 cell_1rw
* cell instance $11565 r0 *1 180.48,60.06
X$11565 578 45 579 644 645 cell_1rw
* cell instance $11566 m0 *1 0.705,62.79
X$11566 67 46 68 644 645 cell_1rw
* cell instance $11567 m0 *1 0,62.79
X$11567 65 46 66 644 645 cell_1rw
* cell instance $11568 m0 *1 1.41,62.79
X$11568 69 46 70 644 645 cell_1rw
* cell instance $11569 m0 *1 2.115,62.79
X$11569 71 46 72 644 645 cell_1rw
* cell instance $11570 m0 *1 2.82,62.79
X$11570 73 46 74 644 645 cell_1rw
* cell instance $11571 m0 *1 3.525,62.79
X$11571 75 46 76 644 645 cell_1rw
* cell instance $11572 m0 *1 4.23,62.79
X$11572 77 46 78 644 645 cell_1rw
* cell instance $11573 m0 *1 4.935,62.79
X$11573 79 46 80 644 645 cell_1rw
* cell instance $11574 m0 *1 5.64,62.79
X$11574 81 46 82 644 645 cell_1rw
* cell instance $11575 m0 *1 6.345,62.79
X$11575 83 46 84 644 645 cell_1rw
* cell instance $11576 m0 *1 7.05,62.79
X$11576 85 46 86 644 645 cell_1rw
* cell instance $11577 m0 *1 7.755,62.79
X$11577 87 46 88 644 645 cell_1rw
* cell instance $11578 m0 *1 8.46,62.79
X$11578 89 46 90 644 645 cell_1rw
* cell instance $11579 m0 *1 9.165,62.79
X$11579 91 46 92 644 645 cell_1rw
* cell instance $11580 m0 *1 9.87,62.79
X$11580 93 46 94 644 645 cell_1rw
* cell instance $11581 m0 *1 10.575,62.79
X$11581 95 46 96 644 645 cell_1rw
* cell instance $11582 m0 *1 11.28,62.79
X$11582 97 46 98 644 645 cell_1rw
* cell instance $11583 m0 *1 11.985,62.79
X$11583 99 46 100 644 645 cell_1rw
* cell instance $11584 m0 *1 12.69,62.79
X$11584 101 46 102 644 645 cell_1rw
* cell instance $11585 m0 *1 13.395,62.79
X$11585 103 46 104 644 645 cell_1rw
* cell instance $11586 m0 *1 14.1,62.79
X$11586 105 46 106 644 645 cell_1rw
* cell instance $11587 m0 *1 14.805,62.79
X$11587 107 46 108 644 645 cell_1rw
* cell instance $11588 m0 *1 15.51,62.79
X$11588 109 46 110 644 645 cell_1rw
* cell instance $11589 m0 *1 16.215,62.79
X$11589 111 46 112 644 645 cell_1rw
* cell instance $11590 m0 *1 16.92,62.79
X$11590 113 46 114 644 645 cell_1rw
* cell instance $11591 m0 *1 17.625,62.79
X$11591 115 46 116 644 645 cell_1rw
* cell instance $11592 m0 *1 18.33,62.79
X$11592 117 46 118 644 645 cell_1rw
* cell instance $11593 m0 *1 19.035,62.79
X$11593 119 46 120 644 645 cell_1rw
* cell instance $11594 m0 *1 19.74,62.79
X$11594 121 46 122 644 645 cell_1rw
* cell instance $11595 m0 *1 20.445,62.79
X$11595 123 46 124 644 645 cell_1rw
* cell instance $11596 m0 *1 21.15,62.79
X$11596 125 46 126 644 645 cell_1rw
* cell instance $11597 m0 *1 21.855,62.79
X$11597 127 46 128 644 645 cell_1rw
* cell instance $11598 m0 *1 22.56,62.79
X$11598 129 46 130 644 645 cell_1rw
* cell instance $11599 m0 *1 23.265,62.79
X$11599 131 46 132 644 645 cell_1rw
* cell instance $11600 m0 *1 23.97,62.79
X$11600 133 46 134 644 645 cell_1rw
* cell instance $11601 m0 *1 24.675,62.79
X$11601 135 46 136 644 645 cell_1rw
* cell instance $11602 m0 *1 25.38,62.79
X$11602 137 46 138 644 645 cell_1rw
* cell instance $11603 m0 *1 26.085,62.79
X$11603 139 46 140 644 645 cell_1rw
* cell instance $11604 m0 *1 26.79,62.79
X$11604 141 46 142 644 645 cell_1rw
* cell instance $11605 m0 *1 27.495,62.79
X$11605 143 46 144 644 645 cell_1rw
* cell instance $11606 m0 *1 28.2,62.79
X$11606 145 46 146 644 645 cell_1rw
* cell instance $11607 m0 *1 28.905,62.79
X$11607 147 46 148 644 645 cell_1rw
* cell instance $11608 m0 *1 29.61,62.79
X$11608 149 46 150 644 645 cell_1rw
* cell instance $11609 m0 *1 30.315,62.79
X$11609 151 46 152 644 645 cell_1rw
* cell instance $11610 m0 *1 31.02,62.79
X$11610 153 46 154 644 645 cell_1rw
* cell instance $11611 m0 *1 31.725,62.79
X$11611 155 46 156 644 645 cell_1rw
* cell instance $11612 m0 *1 32.43,62.79
X$11612 157 46 158 644 645 cell_1rw
* cell instance $11613 m0 *1 33.135,62.79
X$11613 159 46 160 644 645 cell_1rw
* cell instance $11614 m0 *1 33.84,62.79
X$11614 161 46 162 644 645 cell_1rw
* cell instance $11615 m0 *1 34.545,62.79
X$11615 163 46 164 644 645 cell_1rw
* cell instance $11616 m0 *1 35.25,62.79
X$11616 165 46 166 644 645 cell_1rw
* cell instance $11617 m0 *1 35.955,62.79
X$11617 167 46 168 644 645 cell_1rw
* cell instance $11618 m0 *1 36.66,62.79
X$11618 169 46 170 644 645 cell_1rw
* cell instance $11619 m0 *1 37.365,62.79
X$11619 171 46 172 644 645 cell_1rw
* cell instance $11620 m0 *1 38.07,62.79
X$11620 173 46 174 644 645 cell_1rw
* cell instance $11621 m0 *1 38.775,62.79
X$11621 175 46 176 644 645 cell_1rw
* cell instance $11622 m0 *1 39.48,62.79
X$11622 177 46 178 644 645 cell_1rw
* cell instance $11623 m0 *1 40.185,62.79
X$11623 179 46 180 644 645 cell_1rw
* cell instance $11624 m0 *1 40.89,62.79
X$11624 181 46 182 644 645 cell_1rw
* cell instance $11625 m0 *1 41.595,62.79
X$11625 183 46 184 644 645 cell_1rw
* cell instance $11626 m0 *1 42.3,62.79
X$11626 185 46 186 644 645 cell_1rw
* cell instance $11627 m0 *1 43.005,62.79
X$11627 187 46 188 644 645 cell_1rw
* cell instance $11628 m0 *1 43.71,62.79
X$11628 189 46 190 644 645 cell_1rw
* cell instance $11629 m0 *1 44.415,62.79
X$11629 191 46 192 644 645 cell_1rw
* cell instance $11630 m0 *1 45.12,62.79
X$11630 193 46 194 644 645 cell_1rw
* cell instance $11631 m0 *1 45.825,62.79
X$11631 195 46 196 644 645 cell_1rw
* cell instance $11632 m0 *1 46.53,62.79
X$11632 197 46 198 644 645 cell_1rw
* cell instance $11633 m0 *1 47.235,62.79
X$11633 199 46 200 644 645 cell_1rw
* cell instance $11634 m0 *1 47.94,62.79
X$11634 201 46 202 644 645 cell_1rw
* cell instance $11635 m0 *1 48.645,62.79
X$11635 203 46 204 644 645 cell_1rw
* cell instance $11636 m0 *1 49.35,62.79
X$11636 205 46 206 644 645 cell_1rw
* cell instance $11637 m0 *1 50.055,62.79
X$11637 207 46 208 644 645 cell_1rw
* cell instance $11638 m0 *1 50.76,62.79
X$11638 209 46 210 644 645 cell_1rw
* cell instance $11639 m0 *1 51.465,62.79
X$11639 211 46 212 644 645 cell_1rw
* cell instance $11640 m0 *1 52.17,62.79
X$11640 213 46 214 644 645 cell_1rw
* cell instance $11641 m0 *1 52.875,62.79
X$11641 215 46 216 644 645 cell_1rw
* cell instance $11642 m0 *1 53.58,62.79
X$11642 217 46 218 644 645 cell_1rw
* cell instance $11643 m0 *1 54.285,62.79
X$11643 219 46 220 644 645 cell_1rw
* cell instance $11644 m0 *1 54.99,62.79
X$11644 221 46 222 644 645 cell_1rw
* cell instance $11645 m0 *1 55.695,62.79
X$11645 223 46 224 644 645 cell_1rw
* cell instance $11646 m0 *1 56.4,62.79
X$11646 225 46 226 644 645 cell_1rw
* cell instance $11647 m0 *1 57.105,62.79
X$11647 227 46 228 644 645 cell_1rw
* cell instance $11648 m0 *1 57.81,62.79
X$11648 229 46 230 644 645 cell_1rw
* cell instance $11649 m0 *1 58.515,62.79
X$11649 231 46 232 644 645 cell_1rw
* cell instance $11650 m0 *1 59.22,62.79
X$11650 233 46 234 644 645 cell_1rw
* cell instance $11651 m0 *1 59.925,62.79
X$11651 235 46 236 644 645 cell_1rw
* cell instance $11652 m0 *1 60.63,62.79
X$11652 237 46 238 644 645 cell_1rw
* cell instance $11653 m0 *1 61.335,62.79
X$11653 239 46 240 644 645 cell_1rw
* cell instance $11654 m0 *1 62.04,62.79
X$11654 241 46 242 644 645 cell_1rw
* cell instance $11655 m0 *1 62.745,62.79
X$11655 243 46 244 644 645 cell_1rw
* cell instance $11656 m0 *1 63.45,62.79
X$11656 245 46 246 644 645 cell_1rw
* cell instance $11657 m0 *1 64.155,62.79
X$11657 247 46 248 644 645 cell_1rw
* cell instance $11658 m0 *1 64.86,62.79
X$11658 249 46 250 644 645 cell_1rw
* cell instance $11659 m0 *1 65.565,62.79
X$11659 251 46 252 644 645 cell_1rw
* cell instance $11660 m0 *1 66.27,62.79
X$11660 253 46 254 644 645 cell_1rw
* cell instance $11661 m0 *1 66.975,62.79
X$11661 255 46 256 644 645 cell_1rw
* cell instance $11662 m0 *1 67.68,62.79
X$11662 257 46 258 644 645 cell_1rw
* cell instance $11663 m0 *1 68.385,62.79
X$11663 259 46 260 644 645 cell_1rw
* cell instance $11664 m0 *1 69.09,62.79
X$11664 261 46 262 644 645 cell_1rw
* cell instance $11665 m0 *1 69.795,62.79
X$11665 263 46 264 644 645 cell_1rw
* cell instance $11666 m0 *1 70.5,62.79
X$11666 265 46 266 644 645 cell_1rw
* cell instance $11667 m0 *1 71.205,62.79
X$11667 267 46 268 644 645 cell_1rw
* cell instance $11668 m0 *1 71.91,62.79
X$11668 269 46 270 644 645 cell_1rw
* cell instance $11669 m0 *1 72.615,62.79
X$11669 271 46 272 644 645 cell_1rw
* cell instance $11670 m0 *1 73.32,62.79
X$11670 273 46 274 644 645 cell_1rw
* cell instance $11671 m0 *1 74.025,62.79
X$11671 275 46 276 644 645 cell_1rw
* cell instance $11672 m0 *1 74.73,62.79
X$11672 277 46 278 644 645 cell_1rw
* cell instance $11673 m0 *1 75.435,62.79
X$11673 279 46 280 644 645 cell_1rw
* cell instance $11674 m0 *1 76.14,62.79
X$11674 281 46 282 644 645 cell_1rw
* cell instance $11675 m0 *1 76.845,62.79
X$11675 283 46 284 644 645 cell_1rw
* cell instance $11676 m0 *1 77.55,62.79
X$11676 285 46 286 644 645 cell_1rw
* cell instance $11677 m0 *1 78.255,62.79
X$11677 287 46 288 644 645 cell_1rw
* cell instance $11678 m0 *1 78.96,62.79
X$11678 289 46 290 644 645 cell_1rw
* cell instance $11679 m0 *1 79.665,62.79
X$11679 291 46 292 644 645 cell_1rw
* cell instance $11680 m0 *1 80.37,62.79
X$11680 293 46 294 644 645 cell_1rw
* cell instance $11681 m0 *1 81.075,62.79
X$11681 295 46 296 644 645 cell_1rw
* cell instance $11682 m0 *1 81.78,62.79
X$11682 297 46 298 644 645 cell_1rw
* cell instance $11683 m0 *1 82.485,62.79
X$11683 299 46 300 644 645 cell_1rw
* cell instance $11684 m0 *1 83.19,62.79
X$11684 301 46 302 644 645 cell_1rw
* cell instance $11685 m0 *1 83.895,62.79
X$11685 303 46 304 644 645 cell_1rw
* cell instance $11686 m0 *1 84.6,62.79
X$11686 305 46 306 644 645 cell_1rw
* cell instance $11687 m0 *1 85.305,62.79
X$11687 307 46 308 644 645 cell_1rw
* cell instance $11688 m0 *1 86.01,62.79
X$11688 309 46 310 644 645 cell_1rw
* cell instance $11689 m0 *1 86.715,62.79
X$11689 311 46 312 644 645 cell_1rw
* cell instance $11690 m0 *1 87.42,62.79
X$11690 313 46 314 644 645 cell_1rw
* cell instance $11691 m0 *1 88.125,62.79
X$11691 315 46 316 644 645 cell_1rw
* cell instance $11692 m0 *1 88.83,62.79
X$11692 317 46 318 644 645 cell_1rw
* cell instance $11693 m0 *1 89.535,62.79
X$11693 319 46 320 644 645 cell_1rw
* cell instance $11694 m0 *1 90.24,62.79
X$11694 321 46 323 644 645 cell_1rw
* cell instance $11695 m0 *1 90.945,62.79
X$11695 324 46 325 644 645 cell_1rw
* cell instance $11696 m0 *1 91.65,62.79
X$11696 326 46 327 644 645 cell_1rw
* cell instance $11697 m0 *1 92.355,62.79
X$11697 328 46 329 644 645 cell_1rw
* cell instance $11698 m0 *1 93.06,62.79
X$11698 330 46 331 644 645 cell_1rw
* cell instance $11699 m0 *1 93.765,62.79
X$11699 332 46 333 644 645 cell_1rw
* cell instance $11700 m0 *1 94.47,62.79
X$11700 334 46 335 644 645 cell_1rw
* cell instance $11701 m0 *1 95.175,62.79
X$11701 336 46 337 644 645 cell_1rw
* cell instance $11702 m0 *1 95.88,62.79
X$11702 338 46 339 644 645 cell_1rw
* cell instance $11703 m0 *1 96.585,62.79
X$11703 340 46 341 644 645 cell_1rw
* cell instance $11704 m0 *1 97.29,62.79
X$11704 342 46 343 644 645 cell_1rw
* cell instance $11705 m0 *1 97.995,62.79
X$11705 344 46 345 644 645 cell_1rw
* cell instance $11706 m0 *1 98.7,62.79
X$11706 346 46 347 644 645 cell_1rw
* cell instance $11707 m0 *1 99.405,62.79
X$11707 348 46 349 644 645 cell_1rw
* cell instance $11708 m0 *1 100.11,62.79
X$11708 350 46 351 644 645 cell_1rw
* cell instance $11709 m0 *1 100.815,62.79
X$11709 352 46 353 644 645 cell_1rw
* cell instance $11710 m0 *1 101.52,62.79
X$11710 354 46 355 644 645 cell_1rw
* cell instance $11711 m0 *1 102.225,62.79
X$11711 356 46 357 644 645 cell_1rw
* cell instance $11712 m0 *1 102.93,62.79
X$11712 358 46 359 644 645 cell_1rw
* cell instance $11713 m0 *1 103.635,62.79
X$11713 360 46 361 644 645 cell_1rw
* cell instance $11714 m0 *1 104.34,62.79
X$11714 362 46 363 644 645 cell_1rw
* cell instance $11715 m0 *1 105.045,62.79
X$11715 364 46 365 644 645 cell_1rw
* cell instance $11716 m0 *1 105.75,62.79
X$11716 366 46 367 644 645 cell_1rw
* cell instance $11717 m0 *1 106.455,62.79
X$11717 368 46 369 644 645 cell_1rw
* cell instance $11718 m0 *1 107.16,62.79
X$11718 370 46 371 644 645 cell_1rw
* cell instance $11719 m0 *1 107.865,62.79
X$11719 372 46 373 644 645 cell_1rw
* cell instance $11720 m0 *1 108.57,62.79
X$11720 374 46 375 644 645 cell_1rw
* cell instance $11721 m0 *1 109.275,62.79
X$11721 376 46 377 644 645 cell_1rw
* cell instance $11722 m0 *1 109.98,62.79
X$11722 378 46 379 644 645 cell_1rw
* cell instance $11723 m0 *1 110.685,62.79
X$11723 380 46 381 644 645 cell_1rw
* cell instance $11724 m0 *1 111.39,62.79
X$11724 382 46 383 644 645 cell_1rw
* cell instance $11725 m0 *1 112.095,62.79
X$11725 384 46 385 644 645 cell_1rw
* cell instance $11726 m0 *1 112.8,62.79
X$11726 386 46 387 644 645 cell_1rw
* cell instance $11727 m0 *1 113.505,62.79
X$11727 388 46 389 644 645 cell_1rw
* cell instance $11728 m0 *1 114.21,62.79
X$11728 390 46 391 644 645 cell_1rw
* cell instance $11729 m0 *1 114.915,62.79
X$11729 392 46 393 644 645 cell_1rw
* cell instance $11730 m0 *1 115.62,62.79
X$11730 394 46 395 644 645 cell_1rw
* cell instance $11731 m0 *1 116.325,62.79
X$11731 396 46 397 644 645 cell_1rw
* cell instance $11732 m0 *1 117.03,62.79
X$11732 398 46 399 644 645 cell_1rw
* cell instance $11733 m0 *1 117.735,62.79
X$11733 400 46 401 644 645 cell_1rw
* cell instance $11734 m0 *1 118.44,62.79
X$11734 402 46 403 644 645 cell_1rw
* cell instance $11735 m0 *1 119.145,62.79
X$11735 404 46 405 644 645 cell_1rw
* cell instance $11736 m0 *1 119.85,62.79
X$11736 406 46 407 644 645 cell_1rw
* cell instance $11737 m0 *1 120.555,62.79
X$11737 408 46 409 644 645 cell_1rw
* cell instance $11738 m0 *1 121.26,62.79
X$11738 410 46 411 644 645 cell_1rw
* cell instance $11739 m0 *1 121.965,62.79
X$11739 412 46 413 644 645 cell_1rw
* cell instance $11740 m0 *1 122.67,62.79
X$11740 414 46 415 644 645 cell_1rw
* cell instance $11741 m0 *1 123.375,62.79
X$11741 416 46 417 644 645 cell_1rw
* cell instance $11742 m0 *1 124.08,62.79
X$11742 418 46 419 644 645 cell_1rw
* cell instance $11743 m0 *1 124.785,62.79
X$11743 420 46 421 644 645 cell_1rw
* cell instance $11744 m0 *1 125.49,62.79
X$11744 422 46 423 644 645 cell_1rw
* cell instance $11745 m0 *1 126.195,62.79
X$11745 424 46 425 644 645 cell_1rw
* cell instance $11746 m0 *1 126.9,62.79
X$11746 426 46 427 644 645 cell_1rw
* cell instance $11747 m0 *1 127.605,62.79
X$11747 428 46 429 644 645 cell_1rw
* cell instance $11748 m0 *1 128.31,62.79
X$11748 430 46 431 644 645 cell_1rw
* cell instance $11749 m0 *1 129.015,62.79
X$11749 432 46 433 644 645 cell_1rw
* cell instance $11750 m0 *1 129.72,62.79
X$11750 434 46 435 644 645 cell_1rw
* cell instance $11751 m0 *1 130.425,62.79
X$11751 436 46 437 644 645 cell_1rw
* cell instance $11752 m0 *1 131.13,62.79
X$11752 438 46 439 644 645 cell_1rw
* cell instance $11753 m0 *1 131.835,62.79
X$11753 440 46 441 644 645 cell_1rw
* cell instance $11754 m0 *1 132.54,62.79
X$11754 442 46 443 644 645 cell_1rw
* cell instance $11755 m0 *1 133.245,62.79
X$11755 444 46 445 644 645 cell_1rw
* cell instance $11756 m0 *1 133.95,62.79
X$11756 446 46 447 644 645 cell_1rw
* cell instance $11757 m0 *1 134.655,62.79
X$11757 448 46 449 644 645 cell_1rw
* cell instance $11758 m0 *1 135.36,62.79
X$11758 450 46 451 644 645 cell_1rw
* cell instance $11759 m0 *1 136.065,62.79
X$11759 452 46 453 644 645 cell_1rw
* cell instance $11760 m0 *1 136.77,62.79
X$11760 454 46 455 644 645 cell_1rw
* cell instance $11761 m0 *1 137.475,62.79
X$11761 456 46 457 644 645 cell_1rw
* cell instance $11762 m0 *1 138.18,62.79
X$11762 458 46 459 644 645 cell_1rw
* cell instance $11763 m0 *1 138.885,62.79
X$11763 460 46 461 644 645 cell_1rw
* cell instance $11764 m0 *1 139.59,62.79
X$11764 462 46 463 644 645 cell_1rw
* cell instance $11765 m0 *1 140.295,62.79
X$11765 464 46 465 644 645 cell_1rw
* cell instance $11766 m0 *1 141,62.79
X$11766 466 46 467 644 645 cell_1rw
* cell instance $11767 m0 *1 141.705,62.79
X$11767 468 46 469 644 645 cell_1rw
* cell instance $11768 m0 *1 142.41,62.79
X$11768 470 46 471 644 645 cell_1rw
* cell instance $11769 m0 *1 143.115,62.79
X$11769 472 46 473 644 645 cell_1rw
* cell instance $11770 m0 *1 143.82,62.79
X$11770 474 46 475 644 645 cell_1rw
* cell instance $11771 m0 *1 144.525,62.79
X$11771 476 46 477 644 645 cell_1rw
* cell instance $11772 m0 *1 145.23,62.79
X$11772 478 46 479 644 645 cell_1rw
* cell instance $11773 m0 *1 145.935,62.79
X$11773 480 46 481 644 645 cell_1rw
* cell instance $11774 m0 *1 146.64,62.79
X$11774 482 46 483 644 645 cell_1rw
* cell instance $11775 m0 *1 147.345,62.79
X$11775 484 46 485 644 645 cell_1rw
* cell instance $11776 m0 *1 148.05,62.79
X$11776 486 46 487 644 645 cell_1rw
* cell instance $11777 m0 *1 148.755,62.79
X$11777 488 46 489 644 645 cell_1rw
* cell instance $11778 m0 *1 149.46,62.79
X$11778 490 46 491 644 645 cell_1rw
* cell instance $11779 m0 *1 150.165,62.79
X$11779 492 46 493 644 645 cell_1rw
* cell instance $11780 m0 *1 150.87,62.79
X$11780 494 46 495 644 645 cell_1rw
* cell instance $11781 m0 *1 151.575,62.79
X$11781 496 46 497 644 645 cell_1rw
* cell instance $11782 m0 *1 152.28,62.79
X$11782 498 46 499 644 645 cell_1rw
* cell instance $11783 m0 *1 152.985,62.79
X$11783 500 46 501 644 645 cell_1rw
* cell instance $11784 m0 *1 153.69,62.79
X$11784 502 46 503 644 645 cell_1rw
* cell instance $11785 m0 *1 154.395,62.79
X$11785 504 46 505 644 645 cell_1rw
* cell instance $11786 m0 *1 155.1,62.79
X$11786 506 46 507 644 645 cell_1rw
* cell instance $11787 m0 *1 155.805,62.79
X$11787 508 46 509 644 645 cell_1rw
* cell instance $11788 m0 *1 156.51,62.79
X$11788 510 46 511 644 645 cell_1rw
* cell instance $11789 m0 *1 157.215,62.79
X$11789 512 46 513 644 645 cell_1rw
* cell instance $11790 m0 *1 157.92,62.79
X$11790 514 46 515 644 645 cell_1rw
* cell instance $11791 m0 *1 158.625,62.79
X$11791 516 46 517 644 645 cell_1rw
* cell instance $11792 m0 *1 159.33,62.79
X$11792 518 46 519 644 645 cell_1rw
* cell instance $11793 m0 *1 160.035,62.79
X$11793 520 46 521 644 645 cell_1rw
* cell instance $11794 m0 *1 160.74,62.79
X$11794 522 46 523 644 645 cell_1rw
* cell instance $11795 m0 *1 161.445,62.79
X$11795 524 46 525 644 645 cell_1rw
* cell instance $11796 m0 *1 162.15,62.79
X$11796 526 46 527 644 645 cell_1rw
* cell instance $11797 m0 *1 162.855,62.79
X$11797 528 46 529 644 645 cell_1rw
* cell instance $11798 m0 *1 163.56,62.79
X$11798 530 46 531 644 645 cell_1rw
* cell instance $11799 m0 *1 164.265,62.79
X$11799 532 46 533 644 645 cell_1rw
* cell instance $11800 m0 *1 164.97,62.79
X$11800 534 46 535 644 645 cell_1rw
* cell instance $11801 m0 *1 165.675,62.79
X$11801 536 46 537 644 645 cell_1rw
* cell instance $11802 m0 *1 166.38,62.79
X$11802 538 46 539 644 645 cell_1rw
* cell instance $11803 m0 *1 167.085,62.79
X$11803 540 46 541 644 645 cell_1rw
* cell instance $11804 m0 *1 167.79,62.79
X$11804 542 46 543 644 645 cell_1rw
* cell instance $11805 m0 *1 168.495,62.79
X$11805 544 46 545 644 645 cell_1rw
* cell instance $11806 m0 *1 169.2,62.79
X$11806 546 46 547 644 645 cell_1rw
* cell instance $11807 m0 *1 169.905,62.79
X$11807 548 46 549 644 645 cell_1rw
* cell instance $11808 m0 *1 170.61,62.79
X$11808 550 46 551 644 645 cell_1rw
* cell instance $11809 m0 *1 171.315,62.79
X$11809 552 46 553 644 645 cell_1rw
* cell instance $11810 m0 *1 172.02,62.79
X$11810 554 46 555 644 645 cell_1rw
* cell instance $11811 m0 *1 172.725,62.79
X$11811 556 46 557 644 645 cell_1rw
* cell instance $11812 m0 *1 173.43,62.79
X$11812 558 46 559 644 645 cell_1rw
* cell instance $11813 m0 *1 174.135,62.79
X$11813 560 46 561 644 645 cell_1rw
* cell instance $11814 m0 *1 174.84,62.79
X$11814 562 46 563 644 645 cell_1rw
* cell instance $11815 m0 *1 175.545,62.79
X$11815 564 46 565 644 645 cell_1rw
* cell instance $11816 m0 *1 176.25,62.79
X$11816 566 46 567 644 645 cell_1rw
* cell instance $11817 m0 *1 176.955,62.79
X$11817 568 46 569 644 645 cell_1rw
* cell instance $11818 m0 *1 177.66,62.79
X$11818 570 46 571 644 645 cell_1rw
* cell instance $11819 m0 *1 178.365,62.79
X$11819 572 46 573 644 645 cell_1rw
* cell instance $11820 m0 *1 179.07,62.79
X$11820 574 46 575 644 645 cell_1rw
* cell instance $11821 m0 *1 179.775,62.79
X$11821 576 46 577 644 645 cell_1rw
* cell instance $11822 m0 *1 180.48,62.79
X$11822 578 46 579 644 645 cell_1rw
* cell instance $11823 r0 *1 0.705,62.79
X$11823 67 47 68 644 645 cell_1rw
* cell instance $11824 r0 *1 0,62.79
X$11824 65 47 66 644 645 cell_1rw
* cell instance $11825 r0 *1 1.41,62.79
X$11825 69 47 70 644 645 cell_1rw
* cell instance $11826 r0 *1 2.115,62.79
X$11826 71 47 72 644 645 cell_1rw
* cell instance $11827 r0 *1 2.82,62.79
X$11827 73 47 74 644 645 cell_1rw
* cell instance $11828 r0 *1 3.525,62.79
X$11828 75 47 76 644 645 cell_1rw
* cell instance $11829 r0 *1 4.23,62.79
X$11829 77 47 78 644 645 cell_1rw
* cell instance $11830 r0 *1 4.935,62.79
X$11830 79 47 80 644 645 cell_1rw
* cell instance $11831 r0 *1 5.64,62.79
X$11831 81 47 82 644 645 cell_1rw
* cell instance $11832 r0 *1 6.345,62.79
X$11832 83 47 84 644 645 cell_1rw
* cell instance $11833 r0 *1 7.05,62.79
X$11833 85 47 86 644 645 cell_1rw
* cell instance $11834 r0 *1 7.755,62.79
X$11834 87 47 88 644 645 cell_1rw
* cell instance $11835 r0 *1 8.46,62.79
X$11835 89 47 90 644 645 cell_1rw
* cell instance $11836 r0 *1 9.165,62.79
X$11836 91 47 92 644 645 cell_1rw
* cell instance $11837 r0 *1 9.87,62.79
X$11837 93 47 94 644 645 cell_1rw
* cell instance $11838 r0 *1 10.575,62.79
X$11838 95 47 96 644 645 cell_1rw
* cell instance $11839 r0 *1 11.28,62.79
X$11839 97 47 98 644 645 cell_1rw
* cell instance $11840 r0 *1 11.985,62.79
X$11840 99 47 100 644 645 cell_1rw
* cell instance $11841 r0 *1 12.69,62.79
X$11841 101 47 102 644 645 cell_1rw
* cell instance $11842 r0 *1 13.395,62.79
X$11842 103 47 104 644 645 cell_1rw
* cell instance $11843 r0 *1 14.1,62.79
X$11843 105 47 106 644 645 cell_1rw
* cell instance $11844 r0 *1 14.805,62.79
X$11844 107 47 108 644 645 cell_1rw
* cell instance $11845 r0 *1 15.51,62.79
X$11845 109 47 110 644 645 cell_1rw
* cell instance $11846 r0 *1 16.215,62.79
X$11846 111 47 112 644 645 cell_1rw
* cell instance $11847 r0 *1 16.92,62.79
X$11847 113 47 114 644 645 cell_1rw
* cell instance $11848 r0 *1 17.625,62.79
X$11848 115 47 116 644 645 cell_1rw
* cell instance $11849 r0 *1 18.33,62.79
X$11849 117 47 118 644 645 cell_1rw
* cell instance $11850 r0 *1 19.035,62.79
X$11850 119 47 120 644 645 cell_1rw
* cell instance $11851 r0 *1 19.74,62.79
X$11851 121 47 122 644 645 cell_1rw
* cell instance $11852 r0 *1 20.445,62.79
X$11852 123 47 124 644 645 cell_1rw
* cell instance $11853 r0 *1 21.15,62.79
X$11853 125 47 126 644 645 cell_1rw
* cell instance $11854 r0 *1 21.855,62.79
X$11854 127 47 128 644 645 cell_1rw
* cell instance $11855 r0 *1 22.56,62.79
X$11855 129 47 130 644 645 cell_1rw
* cell instance $11856 r0 *1 23.265,62.79
X$11856 131 47 132 644 645 cell_1rw
* cell instance $11857 r0 *1 23.97,62.79
X$11857 133 47 134 644 645 cell_1rw
* cell instance $11858 r0 *1 24.675,62.79
X$11858 135 47 136 644 645 cell_1rw
* cell instance $11859 r0 *1 25.38,62.79
X$11859 137 47 138 644 645 cell_1rw
* cell instance $11860 r0 *1 26.085,62.79
X$11860 139 47 140 644 645 cell_1rw
* cell instance $11861 r0 *1 26.79,62.79
X$11861 141 47 142 644 645 cell_1rw
* cell instance $11862 r0 *1 27.495,62.79
X$11862 143 47 144 644 645 cell_1rw
* cell instance $11863 r0 *1 28.2,62.79
X$11863 145 47 146 644 645 cell_1rw
* cell instance $11864 r0 *1 28.905,62.79
X$11864 147 47 148 644 645 cell_1rw
* cell instance $11865 r0 *1 29.61,62.79
X$11865 149 47 150 644 645 cell_1rw
* cell instance $11866 r0 *1 30.315,62.79
X$11866 151 47 152 644 645 cell_1rw
* cell instance $11867 r0 *1 31.02,62.79
X$11867 153 47 154 644 645 cell_1rw
* cell instance $11868 r0 *1 31.725,62.79
X$11868 155 47 156 644 645 cell_1rw
* cell instance $11869 r0 *1 32.43,62.79
X$11869 157 47 158 644 645 cell_1rw
* cell instance $11870 r0 *1 33.135,62.79
X$11870 159 47 160 644 645 cell_1rw
* cell instance $11871 r0 *1 33.84,62.79
X$11871 161 47 162 644 645 cell_1rw
* cell instance $11872 r0 *1 34.545,62.79
X$11872 163 47 164 644 645 cell_1rw
* cell instance $11873 r0 *1 35.25,62.79
X$11873 165 47 166 644 645 cell_1rw
* cell instance $11874 r0 *1 35.955,62.79
X$11874 167 47 168 644 645 cell_1rw
* cell instance $11875 r0 *1 36.66,62.79
X$11875 169 47 170 644 645 cell_1rw
* cell instance $11876 r0 *1 37.365,62.79
X$11876 171 47 172 644 645 cell_1rw
* cell instance $11877 r0 *1 38.07,62.79
X$11877 173 47 174 644 645 cell_1rw
* cell instance $11878 r0 *1 38.775,62.79
X$11878 175 47 176 644 645 cell_1rw
* cell instance $11879 r0 *1 39.48,62.79
X$11879 177 47 178 644 645 cell_1rw
* cell instance $11880 r0 *1 40.185,62.79
X$11880 179 47 180 644 645 cell_1rw
* cell instance $11881 r0 *1 40.89,62.79
X$11881 181 47 182 644 645 cell_1rw
* cell instance $11882 r0 *1 41.595,62.79
X$11882 183 47 184 644 645 cell_1rw
* cell instance $11883 r0 *1 42.3,62.79
X$11883 185 47 186 644 645 cell_1rw
* cell instance $11884 r0 *1 43.005,62.79
X$11884 187 47 188 644 645 cell_1rw
* cell instance $11885 r0 *1 43.71,62.79
X$11885 189 47 190 644 645 cell_1rw
* cell instance $11886 r0 *1 44.415,62.79
X$11886 191 47 192 644 645 cell_1rw
* cell instance $11887 r0 *1 45.12,62.79
X$11887 193 47 194 644 645 cell_1rw
* cell instance $11888 r0 *1 45.825,62.79
X$11888 195 47 196 644 645 cell_1rw
* cell instance $11889 r0 *1 46.53,62.79
X$11889 197 47 198 644 645 cell_1rw
* cell instance $11890 r0 *1 47.235,62.79
X$11890 199 47 200 644 645 cell_1rw
* cell instance $11891 r0 *1 47.94,62.79
X$11891 201 47 202 644 645 cell_1rw
* cell instance $11892 r0 *1 48.645,62.79
X$11892 203 47 204 644 645 cell_1rw
* cell instance $11893 r0 *1 49.35,62.79
X$11893 205 47 206 644 645 cell_1rw
* cell instance $11894 r0 *1 50.055,62.79
X$11894 207 47 208 644 645 cell_1rw
* cell instance $11895 r0 *1 50.76,62.79
X$11895 209 47 210 644 645 cell_1rw
* cell instance $11896 r0 *1 51.465,62.79
X$11896 211 47 212 644 645 cell_1rw
* cell instance $11897 r0 *1 52.17,62.79
X$11897 213 47 214 644 645 cell_1rw
* cell instance $11898 r0 *1 52.875,62.79
X$11898 215 47 216 644 645 cell_1rw
* cell instance $11899 r0 *1 53.58,62.79
X$11899 217 47 218 644 645 cell_1rw
* cell instance $11900 r0 *1 54.285,62.79
X$11900 219 47 220 644 645 cell_1rw
* cell instance $11901 r0 *1 54.99,62.79
X$11901 221 47 222 644 645 cell_1rw
* cell instance $11902 r0 *1 55.695,62.79
X$11902 223 47 224 644 645 cell_1rw
* cell instance $11903 r0 *1 56.4,62.79
X$11903 225 47 226 644 645 cell_1rw
* cell instance $11904 r0 *1 57.105,62.79
X$11904 227 47 228 644 645 cell_1rw
* cell instance $11905 r0 *1 57.81,62.79
X$11905 229 47 230 644 645 cell_1rw
* cell instance $11906 r0 *1 58.515,62.79
X$11906 231 47 232 644 645 cell_1rw
* cell instance $11907 r0 *1 59.22,62.79
X$11907 233 47 234 644 645 cell_1rw
* cell instance $11908 r0 *1 59.925,62.79
X$11908 235 47 236 644 645 cell_1rw
* cell instance $11909 r0 *1 60.63,62.79
X$11909 237 47 238 644 645 cell_1rw
* cell instance $11910 r0 *1 61.335,62.79
X$11910 239 47 240 644 645 cell_1rw
* cell instance $11911 r0 *1 62.04,62.79
X$11911 241 47 242 644 645 cell_1rw
* cell instance $11912 r0 *1 62.745,62.79
X$11912 243 47 244 644 645 cell_1rw
* cell instance $11913 r0 *1 63.45,62.79
X$11913 245 47 246 644 645 cell_1rw
* cell instance $11914 r0 *1 64.155,62.79
X$11914 247 47 248 644 645 cell_1rw
* cell instance $11915 r0 *1 64.86,62.79
X$11915 249 47 250 644 645 cell_1rw
* cell instance $11916 r0 *1 65.565,62.79
X$11916 251 47 252 644 645 cell_1rw
* cell instance $11917 r0 *1 66.27,62.79
X$11917 253 47 254 644 645 cell_1rw
* cell instance $11918 r0 *1 66.975,62.79
X$11918 255 47 256 644 645 cell_1rw
* cell instance $11919 r0 *1 67.68,62.79
X$11919 257 47 258 644 645 cell_1rw
* cell instance $11920 r0 *1 68.385,62.79
X$11920 259 47 260 644 645 cell_1rw
* cell instance $11921 r0 *1 69.09,62.79
X$11921 261 47 262 644 645 cell_1rw
* cell instance $11922 r0 *1 69.795,62.79
X$11922 263 47 264 644 645 cell_1rw
* cell instance $11923 r0 *1 70.5,62.79
X$11923 265 47 266 644 645 cell_1rw
* cell instance $11924 r0 *1 71.205,62.79
X$11924 267 47 268 644 645 cell_1rw
* cell instance $11925 r0 *1 71.91,62.79
X$11925 269 47 270 644 645 cell_1rw
* cell instance $11926 r0 *1 72.615,62.79
X$11926 271 47 272 644 645 cell_1rw
* cell instance $11927 r0 *1 73.32,62.79
X$11927 273 47 274 644 645 cell_1rw
* cell instance $11928 r0 *1 74.025,62.79
X$11928 275 47 276 644 645 cell_1rw
* cell instance $11929 r0 *1 74.73,62.79
X$11929 277 47 278 644 645 cell_1rw
* cell instance $11930 r0 *1 75.435,62.79
X$11930 279 47 280 644 645 cell_1rw
* cell instance $11931 r0 *1 76.14,62.79
X$11931 281 47 282 644 645 cell_1rw
* cell instance $11932 r0 *1 76.845,62.79
X$11932 283 47 284 644 645 cell_1rw
* cell instance $11933 r0 *1 77.55,62.79
X$11933 285 47 286 644 645 cell_1rw
* cell instance $11934 r0 *1 78.255,62.79
X$11934 287 47 288 644 645 cell_1rw
* cell instance $11935 r0 *1 78.96,62.79
X$11935 289 47 290 644 645 cell_1rw
* cell instance $11936 r0 *1 79.665,62.79
X$11936 291 47 292 644 645 cell_1rw
* cell instance $11937 r0 *1 80.37,62.79
X$11937 293 47 294 644 645 cell_1rw
* cell instance $11938 r0 *1 81.075,62.79
X$11938 295 47 296 644 645 cell_1rw
* cell instance $11939 r0 *1 81.78,62.79
X$11939 297 47 298 644 645 cell_1rw
* cell instance $11940 r0 *1 82.485,62.79
X$11940 299 47 300 644 645 cell_1rw
* cell instance $11941 r0 *1 83.19,62.79
X$11941 301 47 302 644 645 cell_1rw
* cell instance $11942 r0 *1 83.895,62.79
X$11942 303 47 304 644 645 cell_1rw
* cell instance $11943 r0 *1 84.6,62.79
X$11943 305 47 306 644 645 cell_1rw
* cell instance $11944 r0 *1 85.305,62.79
X$11944 307 47 308 644 645 cell_1rw
* cell instance $11945 r0 *1 86.01,62.79
X$11945 309 47 310 644 645 cell_1rw
* cell instance $11946 r0 *1 86.715,62.79
X$11946 311 47 312 644 645 cell_1rw
* cell instance $11947 r0 *1 87.42,62.79
X$11947 313 47 314 644 645 cell_1rw
* cell instance $11948 r0 *1 88.125,62.79
X$11948 315 47 316 644 645 cell_1rw
* cell instance $11949 r0 *1 88.83,62.79
X$11949 317 47 318 644 645 cell_1rw
* cell instance $11950 r0 *1 89.535,62.79
X$11950 319 47 320 644 645 cell_1rw
* cell instance $11951 r0 *1 90.24,62.79
X$11951 321 47 323 644 645 cell_1rw
* cell instance $11952 r0 *1 90.945,62.79
X$11952 324 47 325 644 645 cell_1rw
* cell instance $11953 r0 *1 91.65,62.79
X$11953 326 47 327 644 645 cell_1rw
* cell instance $11954 r0 *1 92.355,62.79
X$11954 328 47 329 644 645 cell_1rw
* cell instance $11955 r0 *1 93.06,62.79
X$11955 330 47 331 644 645 cell_1rw
* cell instance $11956 r0 *1 93.765,62.79
X$11956 332 47 333 644 645 cell_1rw
* cell instance $11957 r0 *1 94.47,62.79
X$11957 334 47 335 644 645 cell_1rw
* cell instance $11958 r0 *1 95.175,62.79
X$11958 336 47 337 644 645 cell_1rw
* cell instance $11959 r0 *1 95.88,62.79
X$11959 338 47 339 644 645 cell_1rw
* cell instance $11960 r0 *1 96.585,62.79
X$11960 340 47 341 644 645 cell_1rw
* cell instance $11961 r0 *1 97.29,62.79
X$11961 342 47 343 644 645 cell_1rw
* cell instance $11962 r0 *1 97.995,62.79
X$11962 344 47 345 644 645 cell_1rw
* cell instance $11963 r0 *1 98.7,62.79
X$11963 346 47 347 644 645 cell_1rw
* cell instance $11964 r0 *1 99.405,62.79
X$11964 348 47 349 644 645 cell_1rw
* cell instance $11965 r0 *1 100.11,62.79
X$11965 350 47 351 644 645 cell_1rw
* cell instance $11966 r0 *1 100.815,62.79
X$11966 352 47 353 644 645 cell_1rw
* cell instance $11967 r0 *1 101.52,62.79
X$11967 354 47 355 644 645 cell_1rw
* cell instance $11968 r0 *1 102.225,62.79
X$11968 356 47 357 644 645 cell_1rw
* cell instance $11969 r0 *1 102.93,62.79
X$11969 358 47 359 644 645 cell_1rw
* cell instance $11970 r0 *1 103.635,62.79
X$11970 360 47 361 644 645 cell_1rw
* cell instance $11971 r0 *1 104.34,62.79
X$11971 362 47 363 644 645 cell_1rw
* cell instance $11972 r0 *1 105.045,62.79
X$11972 364 47 365 644 645 cell_1rw
* cell instance $11973 r0 *1 105.75,62.79
X$11973 366 47 367 644 645 cell_1rw
* cell instance $11974 r0 *1 106.455,62.79
X$11974 368 47 369 644 645 cell_1rw
* cell instance $11975 r0 *1 107.16,62.79
X$11975 370 47 371 644 645 cell_1rw
* cell instance $11976 r0 *1 107.865,62.79
X$11976 372 47 373 644 645 cell_1rw
* cell instance $11977 r0 *1 108.57,62.79
X$11977 374 47 375 644 645 cell_1rw
* cell instance $11978 r0 *1 109.275,62.79
X$11978 376 47 377 644 645 cell_1rw
* cell instance $11979 r0 *1 109.98,62.79
X$11979 378 47 379 644 645 cell_1rw
* cell instance $11980 r0 *1 110.685,62.79
X$11980 380 47 381 644 645 cell_1rw
* cell instance $11981 r0 *1 111.39,62.79
X$11981 382 47 383 644 645 cell_1rw
* cell instance $11982 r0 *1 112.095,62.79
X$11982 384 47 385 644 645 cell_1rw
* cell instance $11983 r0 *1 112.8,62.79
X$11983 386 47 387 644 645 cell_1rw
* cell instance $11984 r0 *1 113.505,62.79
X$11984 388 47 389 644 645 cell_1rw
* cell instance $11985 r0 *1 114.21,62.79
X$11985 390 47 391 644 645 cell_1rw
* cell instance $11986 r0 *1 114.915,62.79
X$11986 392 47 393 644 645 cell_1rw
* cell instance $11987 r0 *1 115.62,62.79
X$11987 394 47 395 644 645 cell_1rw
* cell instance $11988 r0 *1 116.325,62.79
X$11988 396 47 397 644 645 cell_1rw
* cell instance $11989 r0 *1 117.03,62.79
X$11989 398 47 399 644 645 cell_1rw
* cell instance $11990 r0 *1 117.735,62.79
X$11990 400 47 401 644 645 cell_1rw
* cell instance $11991 r0 *1 118.44,62.79
X$11991 402 47 403 644 645 cell_1rw
* cell instance $11992 r0 *1 119.145,62.79
X$11992 404 47 405 644 645 cell_1rw
* cell instance $11993 r0 *1 119.85,62.79
X$11993 406 47 407 644 645 cell_1rw
* cell instance $11994 r0 *1 120.555,62.79
X$11994 408 47 409 644 645 cell_1rw
* cell instance $11995 r0 *1 121.26,62.79
X$11995 410 47 411 644 645 cell_1rw
* cell instance $11996 r0 *1 121.965,62.79
X$11996 412 47 413 644 645 cell_1rw
* cell instance $11997 r0 *1 122.67,62.79
X$11997 414 47 415 644 645 cell_1rw
* cell instance $11998 r0 *1 123.375,62.79
X$11998 416 47 417 644 645 cell_1rw
* cell instance $11999 r0 *1 124.08,62.79
X$11999 418 47 419 644 645 cell_1rw
* cell instance $12000 r0 *1 124.785,62.79
X$12000 420 47 421 644 645 cell_1rw
* cell instance $12001 r0 *1 125.49,62.79
X$12001 422 47 423 644 645 cell_1rw
* cell instance $12002 r0 *1 126.195,62.79
X$12002 424 47 425 644 645 cell_1rw
* cell instance $12003 r0 *1 126.9,62.79
X$12003 426 47 427 644 645 cell_1rw
* cell instance $12004 r0 *1 127.605,62.79
X$12004 428 47 429 644 645 cell_1rw
* cell instance $12005 r0 *1 128.31,62.79
X$12005 430 47 431 644 645 cell_1rw
* cell instance $12006 r0 *1 129.015,62.79
X$12006 432 47 433 644 645 cell_1rw
* cell instance $12007 r0 *1 129.72,62.79
X$12007 434 47 435 644 645 cell_1rw
* cell instance $12008 r0 *1 130.425,62.79
X$12008 436 47 437 644 645 cell_1rw
* cell instance $12009 r0 *1 131.13,62.79
X$12009 438 47 439 644 645 cell_1rw
* cell instance $12010 r0 *1 131.835,62.79
X$12010 440 47 441 644 645 cell_1rw
* cell instance $12011 r0 *1 132.54,62.79
X$12011 442 47 443 644 645 cell_1rw
* cell instance $12012 r0 *1 133.245,62.79
X$12012 444 47 445 644 645 cell_1rw
* cell instance $12013 r0 *1 133.95,62.79
X$12013 446 47 447 644 645 cell_1rw
* cell instance $12014 r0 *1 134.655,62.79
X$12014 448 47 449 644 645 cell_1rw
* cell instance $12015 r0 *1 135.36,62.79
X$12015 450 47 451 644 645 cell_1rw
* cell instance $12016 r0 *1 136.065,62.79
X$12016 452 47 453 644 645 cell_1rw
* cell instance $12017 r0 *1 136.77,62.79
X$12017 454 47 455 644 645 cell_1rw
* cell instance $12018 r0 *1 137.475,62.79
X$12018 456 47 457 644 645 cell_1rw
* cell instance $12019 r0 *1 138.18,62.79
X$12019 458 47 459 644 645 cell_1rw
* cell instance $12020 r0 *1 138.885,62.79
X$12020 460 47 461 644 645 cell_1rw
* cell instance $12021 r0 *1 139.59,62.79
X$12021 462 47 463 644 645 cell_1rw
* cell instance $12022 r0 *1 140.295,62.79
X$12022 464 47 465 644 645 cell_1rw
* cell instance $12023 r0 *1 141,62.79
X$12023 466 47 467 644 645 cell_1rw
* cell instance $12024 r0 *1 141.705,62.79
X$12024 468 47 469 644 645 cell_1rw
* cell instance $12025 r0 *1 142.41,62.79
X$12025 470 47 471 644 645 cell_1rw
* cell instance $12026 r0 *1 143.115,62.79
X$12026 472 47 473 644 645 cell_1rw
* cell instance $12027 r0 *1 143.82,62.79
X$12027 474 47 475 644 645 cell_1rw
* cell instance $12028 r0 *1 144.525,62.79
X$12028 476 47 477 644 645 cell_1rw
* cell instance $12029 r0 *1 145.23,62.79
X$12029 478 47 479 644 645 cell_1rw
* cell instance $12030 r0 *1 145.935,62.79
X$12030 480 47 481 644 645 cell_1rw
* cell instance $12031 r0 *1 146.64,62.79
X$12031 482 47 483 644 645 cell_1rw
* cell instance $12032 r0 *1 147.345,62.79
X$12032 484 47 485 644 645 cell_1rw
* cell instance $12033 r0 *1 148.05,62.79
X$12033 486 47 487 644 645 cell_1rw
* cell instance $12034 r0 *1 148.755,62.79
X$12034 488 47 489 644 645 cell_1rw
* cell instance $12035 r0 *1 149.46,62.79
X$12035 490 47 491 644 645 cell_1rw
* cell instance $12036 r0 *1 150.165,62.79
X$12036 492 47 493 644 645 cell_1rw
* cell instance $12037 r0 *1 150.87,62.79
X$12037 494 47 495 644 645 cell_1rw
* cell instance $12038 r0 *1 151.575,62.79
X$12038 496 47 497 644 645 cell_1rw
* cell instance $12039 r0 *1 152.28,62.79
X$12039 498 47 499 644 645 cell_1rw
* cell instance $12040 r0 *1 152.985,62.79
X$12040 500 47 501 644 645 cell_1rw
* cell instance $12041 r0 *1 153.69,62.79
X$12041 502 47 503 644 645 cell_1rw
* cell instance $12042 r0 *1 154.395,62.79
X$12042 504 47 505 644 645 cell_1rw
* cell instance $12043 r0 *1 155.1,62.79
X$12043 506 47 507 644 645 cell_1rw
* cell instance $12044 r0 *1 155.805,62.79
X$12044 508 47 509 644 645 cell_1rw
* cell instance $12045 r0 *1 156.51,62.79
X$12045 510 47 511 644 645 cell_1rw
* cell instance $12046 r0 *1 157.215,62.79
X$12046 512 47 513 644 645 cell_1rw
* cell instance $12047 r0 *1 157.92,62.79
X$12047 514 47 515 644 645 cell_1rw
* cell instance $12048 r0 *1 158.625,62.79
X$12048 516 47 517 644 645 cell_1rw
* cell instance $12049 r0 *1 159.33,62.79
X$12049 518 47 519 644 645 cell_1rw
* cell instance $12050 r0 *1 160.035,62.79
X$12050 520 47 521 644 645 cell_1rw
* cell instance $12051 r0 *1 160.74,62.79
X$12051 522 47 523 644 645 cell_1rw
* cell instance $12052 r0 *1 161.445,62.79
X$12052 524 47 525 644 645 cell_1rw
* cell instance $12053 r0 *1 162.15,62.79
X$12053 526 47 527 644 645 cell_1rw
* cell instance $12054 r0 *1 162.855,62.79
X$12054 528 47 529 644 645 cell_1rw
* cell instance $12055 r0 *1 163.56,62.79
X$12055 530 47 531 644 645 cell_1rw
* cell instance $12056 r0 *1 164.265,62.79
X$12056 532 47 533 644 645 cell_1rw
* cell instance $12057 r0 *1 164.97,62.79
X$12057 534 47 535 644 645 cell_1rw
* cell instance $12058 r0 *1 165.675,62.79
X$12058 536 47 537 644 645 cell_1rw
* cell instance $12059 r0 *1 166.38,62.79
X$12059 538 47 539 644 645 cell_1rw
* cell instance $12060 r0 *1 167.085,62.79
X$12060 540 47 541 644 645 cell_1rw
* cell instance $12061 r0 *1 167.79,62.79
X$12061 542 47 543 644 645 cell_1rw
* cell instance $12062 r0 *1 168.495,62.79
X$12062 544 47 545 644 645 cell_1rw
* cell instance $12063 r0 *1 169.2,62.79
X$12063 546 47 547 644 645 cell_1rw
* cell instance $12064 r0 *1 169.905,62.79
X$12064 548 47 549 644 645 cell_1rw
* cell instance $12065 r0 *1 170.61,62.79
X$12065 550 47 551 644 645 cell_1rw
* cell instance $12066 r0 *1 171.315,62.79
X$12066 552 47 553 644 645 cell_1rw
* cell instance $12067 r0 *1 172.02,62.79
X$12067 554 47 555 644 645 cell_1rw
* cell instance $12068 r0 *1 172.725,62.79
X$12068 556 47 557 644 645 cell_1rw
* cell instance $12069 r0 *1 173.43,62.79
X$12069 558 47 559 644 645 cell_1rw
* cell instance $12070 r0 *1 174.135,62.79
X$12070 560 47 561 644 645 cell_1rw
* cell instance $12071 r0 *1 174.84,62.79
X$12071 562 47 563 644 645 cell_1rw
* cell instance $12072 r0 *1 175.545,62.79
X$12072 564 47 565 644 645 cell_1rw
* cell instance $12073 r0 *1 176.25,62.79
X$12073 566 47 567 644 645 cell_1rw
* cell instance $12074 r0 *1 176.955,62.79
X$12074 568 47 569 644 645 cell_1rw
* cell instance $12075 r0 *1 177.66,62.79
X$12075 570 47 571 644 645 cell_1rw
* cell instance $12076 r0 *1 178.365,62.79
X$12076 572 47 573 644 645 cell_1rw
* cell instance $12077 r0 *1 179.07,62.79
X$12077 574 47 575 644 645 cell_1rw
* cell instance $12078 r0 *1 179.775,62.79
X$12078 576 47 577 644 645 cell_1rw
* cell instance $12079 r0 *1 180.48,62.79
X$12079 578 47 579 644 645 cell_1rw
* cell instance $12080 m0 *1 0.705,65.52
X$12080 67 48 68 644 645 cell_1rw
* cell instance $12081 m0 *1 0,65.52
X$12081 65 48 66 644 645 cell_1rw
* cell instance $12082 m0 *1 1.41,65.52
X$12082 69 48 70 644 645 cell_1rw
* cell instance $12083 m0 *1 2.115,65.52
X$12083 71 48 72 644 645 cell_1rw
* cell instance $12084 m0 *1 2.82,65.52
X$12084 73 48 74 644 645 cell_1rw
* cell instance $12085 m0 *1 3.525,65.52
X$12085 75 48 76 644 645 cell_1rw
* cell instance $12086 m0 *1 4.23,65.52
X$12086 77 48 78 644 645 cell_1rw
* cell instance $12087 m0 *1 4.935,65.52
X$12087 79 48 80 644 645 cell_1rw
* cell instance $12088 m0 *1 5.64,65.52
X$12088 81 48 82 644 645 cell_1rw
* cell instance $12089 m0 *1 6.345,65.52
X$12089 83 48 84 644 645 cell_1rw
* cell instance $12090 m0 *1 7.05,65.52
X$12090 85 48 86 644 645 cell_1rw
* cell instance $12091 m0 *1 7.755,65.52
X$12091 87 48 88 644 645 cell_1rw
* cell instance $12092 m0 *1 8.46,65.52
X$12092 89 48 90 644 645 cell_1rw
* cell instance $12093 m0 *1 9.165,65.52
X$12093 91 48 92 644 645 cell_1rw
* cell instance $12094 m0 *1 9.87,65.52
X$12094 93 48 94 644 645 cell_1rw
* cell instance $12095 m0 *1 10.575,65.52
X$12095 95 48 96 644 645 cell_1rw
* cell instance $12096 m0 *1 11.28,65.52
X$12096 97 48 98 644 645 cell_1rw
* cell instance $12097 m0 *1 11.985,65.52
X$12097 99 48 100 644 645 cell_1rw
* cell instance $12098 m0 *1 12.69,65.52
X$12098 101 48 102 644 645 cell_1rw
* cell instance $12099 m0 *1 13.395,65.52
X$12099 103 48 104 644 645 cell_1rw
* cell instance $12100 m0 *1 14.1,65.52
X$12100 105 48 106 644 645 cell_1rw
* cell instance $12101 m0 *1 14.805,65.52
X$12101 107 48 108 644 645 cell_1rw
* cell instance $12102 m0 *1 15.51,65.52
X$12102 109 48 110 644 645 cell_1rw
* cell instance $12103 m0 *1 16.215,65.52
X$12103 111 48 112 644 645 cell_1rw
* cell instance $12104 m0 *1 16.92,65.52
X$12104 113 48 114 644 645 cell_1rw
* cell instance $12105 m0 *1 17.625,65.52
X$12105 115 48 116 644 645 cell_1rw
* cell instance $12106 m0 *1 18.33,65.52
X$12106 117 48 118 644 645 cell_1rw
* cell instance $12107 m0 *1 19.035,65.52
X$12107 119 48 120 644 645 cell_1rw
* cell instance $12108 m0 *1 19.74,65.52
X$12108 121 48 122 644 645 cell_1rw
* cell instance $12109 m0 *1 20.445,65.52
X$12109 123 48 124 644 645 cell_1rw
* cell instance $12110 m0 *1 21.15,65.52
X$12110 125 48 126 644 645 cell_1rw
* cell instance $12111 m0 *1 21.855,65.52
X$12111 127 48 128 644 645 cell_1rw
* cell instance $12112 m0 *1 22.56,65.52
X$12112 129 48 130 644 645 cell_1rw
* cell instance $12113 m0 *1 23.265,65.52
X$12113 131 48 132 644 645 cell_1rw
* cell instance $12114 m0 *1 23.97,65.52
X$12114 133 48 134 644 645 cell_1rw
* cell instance $12115 m0 *1 24.675,65.52
X$12115 135 48 136 644 645 cell_1rw
* cell instance $12116 m0 *1 25.38,65.52
X$12116 137 48 138 644 645 cell_1rw
* cell instance $12117 m0 *1 26.085,65.52
X$12117 139 48 140 644 645 cell_1rw
* cell instance $12118 m0 *1 26.79,65.52
X$12118 141 48 142 644 645 cell_1rw
* cell instance $12119 m0 *1 27.495,65.52
X$12119 143 48 144 644 645 cell_1rw
* cell instance $12120 m0 *1 28.2,65.52
X$12120 145 48 146 644 645 cell_1rw
* cell instance $12121 m0 *1 28.905,65.52
X$12121 147 48 148 644 645 cell_1rw
* cell instance $12122 m0 *1 29.61,65.52
X$12122 149 48 150 644 645 cell_1rw
* cell instance $12123 m0 *1 30.315,65.52
X$12123 151 48 152 644 645 cell_1rw
* cell instance $12124 m0 *1 31.02,65.52
X$12124 153 48 154 644 645 cell_1rw
* cell instance $12125 m0 *1 31.725,65.52
X$12125 155 48 156 644 645 cell_1rw
* cell instance $12126 m0 *1 32.43,65.52
X$12126 157 48 158 644 645 cell_1rw
* cell instance $12127 m0 *1 33.135,65.52
X$12127 159 48 160 644 645 cell_1rw
* cell instance $12128 m0 *1 33.84,65.52
X$12128 161 48 162 644 645 cell_1rw
* cell instance $12129 m0 *1 34.545,65.52
X$12129 163 48 164 644 645 cell_1rw
* cell instance $12130 m0 *1 35.25,65.52
X$12130 165 48 166 644 645 cell_1rw
* cell instance $12131 m0 *1 35.955,65.52
X$12131 167 48 168 644 645 cell_1rw
* cell instance $12132 m0 *1 36.66,65.52
X$12132 169 48 170 644 645 cell_1rw
* cell instance $12133 m0 *1 37.365,65.52
X$12133 171 48 172 644 645 cell_1rw
* cell instance $12134 m0 *1 38.07,65.52
X$12134 173 48 174 644 645 cell_1rw
* cell instance $12135 m0 *1 38.775,65.52
X$12135 175 48 176 644 645 cell_1rw
* cell instance $12136 m0 *1 39.48,65.52
X$12136 177 48 178 644 645 cell_1rw
* cell instance $12137 m0 *1 40.185,65.52
X$12137 179 48 180 644 645 cell_1rw
* cell instance $12138 m0 *1 40.89,65.52
X$12138 181 48 182 644 645 cell_1rw
* cell instance $12139 m0 *1 41.595,65.52
X$12139 183 48 184 644 645 cell_1rw
* cell instance $12140 m0 *1 42.3,65.52
X$12140 185 48 186 644 645 cell_1rw
* cell instance $12141 m0 *1 43.005,65.52
X$12141 187 48 188 644 645 cell_1rw
* cell instance $12142 m0 *1 43.71,65.52
X$12142 189 48 190 644 645 cell_1rw
* cell instance $12143 m0 *1 44.415,65.52
X$12143 191 48 192 644 645 cell_1rw
* cell instance $12144 m0 *1 45.12,65.52
X$12144 193 48 194 644 645 cell_1rw
* cell instance $12145 m0 *1 45.825,65.52
X$12145 195 48 196 644 645 cell_1rw
* cell instance $12146 m0 *1 46.53,65.52
X$12146 197 48 198 644 645 cell_1rw
* cell instance $12147 m0 *1 47.235,65.52
X$12147 199 48 200 644 645 cell_1rw
* cell instance $12148 m0 *1 47.94,65.52
X$12148 201 48 202 644 645 cell_1rw
* cell instance $12149 m0 *1 48.645,65.52
X$12149 203 48 204 644 645 cell_1rw
* cell instance $12150 m0 *1 49.35,65.52
X$12150 205 48 206 644 645 cell_1rw
* cell instance $12151 m0 *1 50.055,65.52
X$12151 207 48 208 644 645 cell_1rw
* cell instance $12152 m0 *1 50.76,65.52
X$12152 209 48 210 644 645 cell_1rw
* cell instance $12153 m0 *1 51.465,65.52
X$12153 211 48 212 644 645 cell_1rw
* cell instance $12154 m0 *1 52.17,65.52
X$12154 213 48 214 644 645 cell_1rw
* cell instance $12155 m0 *1 52.875,65.52
X$12155 215 48 216 644 645 cell_1rw
* cell instance $12156 m0 *1 53.58,65.52
X$12156 217 48 218 644 645 cell_1rw
* cell instance $12157 m0 *1 54.285,65.52
X$12157 219 48 220 644 645 cell_1rw
* cell instance $12158 m0 *1 54.99,65.52
X$12158 221 48 222 644 645 cell_1rw
* cell instance $12159 m0 *1 55.695,65.52
X$12159 223 48 224 644 645 cell_1rw
* cell instance $12160 m0 *1 56.4,65.52
X$12160 225 48 226 644 645 cell_1rw
* cell instance $12161 m0 *1 57.105,65.52
X$12161 227 48 228 644 645 cell_1rw
* cell instance $12162 m0 *1 57.81,65.52
X$12162 229 48 230 644 645 cell_1rw
* cell instance $12163 m0 *1 58.515,65.52
X$12163 231 48 232 644 645 cell_1rw
* cell instance $12164 m0 *1 59.22,65.52
X$12164 233 48 234 644 645 cell_1rw
* cell instance $12165 m0 *1 59.925,65.52
X$12165 235 48 236 644 645 cell_1rw
* cell instance $12166 m0 *1 60.63,65.52
X$12166 237 48 238 644 645 cell_1rw
* cell instance $12167 m0 *1 61.335,65.52
X$12167 239 48 240 644 645 cell_1rw
* cell instance $12168 m0 *1 62.04,65.52
X$12168 241 48 242 644 645 cell_1rw
* cell instance $12169 m0 *1 62.745,65.52
X$12169 243 48 244 644 645 cell_1rw
* cell instance $12170 m0 *1 63.45,65.52
X$12170 245 48 246 644 645 cell_1rw
* cell instance $12171 m0 *1 64.155,65.52
X$12171 247 48 248 644 645 cell_1rw
* cell instance $12172 m0 *1 64.86,65.52
X$12172 249 48 250 644 645 cell_1rw
* cell instance $12173 m0 *1 65.565,65.52
X$12173 251 48 252 644 645 cell_1rw
* cell instance $12174 m0 *1 66.27,65.52
X$12174 253 48 254 644 645 cell_1rw
* cell instance $12175 m0 *1 66.975,65.52
X$12175 255 48 256 644 645 cell_1rw
* cell instance $12176 m0 *1 67.68,65.52
X$12176 257 48 258 644 645 cell_1rw
* cell instance $12177 m0 *1 68.385,65.52
X$12177 259 48 260 644 645 cell_1rw
* cell instance $12178 m0 *1 69.09,65.52
X$12178 261 48 262 644 645 cell_1rw
* cell instance $12179 m0 *1 69.795,65.52
X$12179 263 48 264 644 645 cell_1rw
* cell instance $12180 m0 *1 70.5,65.52
X$12180 265 48 266 644 645 cell_1rw
* cell instance $12181 m0 *1 71.205,65.52
X$12181 267 48 268 644 645 cell_1rw
* cell instance $12182 m0 *1 71.91,65.52
X$12182 269 48 270 644 645 cell_1rw
* cell instance $12183 m0 *1 72.615,65.52
X$12183 271 48 272 644 645 cell_1rw
* cell instance $12184 m0 *1 73.32,65.52
X$12184 273 48 274 644 645 cell_1rw
* cell instance $12185 m0 *1 74.025,65.52
X$12185 275 48 276 644 645 cell_1rw
* cell instance $12186 m0 *1 74.73,65.52
X$12186 277 48 278 644 645 cell_1rw
* cell instance $12187 m0 *1 75.435,65.52
X$12187 279 48 280 644 645 cell_1rw
* cell instance $12188 m0 *1 76.14,65.52
X$12188 281 48 282 644 645 cell_1rw
* cell instance $12189 m0 *1 76.845,65.52
X$12189 283 48 284 644 645 cell_1rw
* cell instance $12190 m0 *1 77.55,65.52
X$12190 285 48 286 644 645 cell_1rw
* cell instance $12191 m0 *1 78.255,65.52
X$12191 287 48 288 644 645 cell_1rw
* cell instance $12192 m0 *1 78.96,65.52
X$12192 289 48 290 644 645 cell_1rw
* cell instance $12193 m0 *1 79.665,65.52
X$12193 291 48 292 644 645 cell_1rw
* cell instance $12194 m0 *1 80.37,65.52
X$12194 293 48 294 644 645 cell_1rw
* cell instance $12195 m0 *1 81.075,65.52
X$12195 295 48 296 644 645 cell_1rw
* cell instance $12196 m0 *1 81.78,65.52
X$12196 297 48 298 644 645 cell_1rw
* cell instance $12197 m0 *1 82.485,65.52
X$12197 299 48 300 644 645 cell_1rw
* cell instance $12198 m0 *1 83.19,65.52
X$12198 301 48 302 644 645 cell_1rw
* cell instance $12199 m0 *1 83.895,65.52
X$12199 303 48 304 644 645 cell_1rw
* cell instance $12200 m0 *1 84.6,65.52
X$12200 305 48 306 644 645 cell_1rw
* cell instance $12201 m0 *1 85.305,65.52
X$12201 307 48 308 644 645 cell_1rw
* cell instance $12202 m0 *1 86.01,65.52
X$12202 309 48 310 644 645 cell_1rw
* cell instance $12203 m0 *1 86.715,65.52
X$12203 311 48 312 644 645 cell_1rw
* cell instance $12204 m0 *1 87.42,65.52
X$12204 313 48 314 644 645 cell_1rw
* cell instance $12205 m0 *1 88.125,65.52
X$12205 315 48 316 644 645 cell_1rw
* cell instance $12206 m0 *1 88.83,65.52
X$12206 317 48 318 644 645 cell_1rw
* cell instance $12207 m0 *1 89.535,65.52
X$12207 319 48 320 644 645 cell_1rw
* cell instance $12208 m0 *1 90.24,65.52
X$12208 321 48 323 644 645 cell_1rw
* cell instance $12209 m0 *1 90.945,65.52
X$12209 324 48 325 644 645 cell_1rw
* cell instance $12210 m0 *1 91.65,65.52
X$12210 326 48 327 644 645 cell_1rw
* cell instance $12211 m0 *1 92.355,65.52
X$12211 328 48 329 644 645 cell_1rw
* cell instance $12212 m0 *1 93.06,65.52
X$12212 330 48 331 644 645 cell_1rw
* cell instance $12213 m0 *1 93.765,65.52
X$12213 332 48 333 644 645 cell_1rw
* cell instance $12214 m0 *1 94.47,65.52
X$12214 334 48 335 644 645 cell_1rw
* cell instance $12215 m0 *1 95.175,65.52
X$12215 336 48 337 644 645 cell_1rw
* cell instance $12216 m0 *1 95.88,65.52
X$12216 338 48 339 644 645 cell_1rw
* cell instance $12217 m0 *1 96.585,65.52
X$12217 340 48 341 644 645 cell_1rw
* cell instance $12218 m0 *1 97.29,65.52
X$12218 342 48 343 644 645 cell_1rw
* cell instance $12219 m0 *1 97.995,65.52
X$12219 344 48 345 644 645 cell_1rw
* cell instance $12220 m0 *1 98.7,65.52
X$12220 346 48 347 644 645 cell_1rw
* cell instance $12221 m0 *1 99.405,65.52
X$12221 348 48 349 644 645 cell_1rw
* cell instance $12222 m0 *1 100.11,65.52
X$12222 350 48 351 644 645 cell_1rw
* cell instance $12223 m0 *1 100.815,65.52
X$12223 352 48 353 644 645 cell_1rw
* cell instance $12224 m0 *1 101.52,65.52
X$12224 354 48 355 644 645 cell_1rw
* cell instance $12225 m0 *1 102.225,65.52
X$12225 356 48 357 644 645 cell_1rw
* cell instance $12226 m0 *1 102.93,65.52
X$12226 358 48 359 644 645 cell_1rw
* cell instance $12227 m0 *1 103.635,65.52
X$12227 360 48 361 644 645 cell_1rw
* cell instance $12228 m0 *1 104.34,65.52
X$12228 362 48 363 644 645 cell_1rw
* cell instance $12229 m0 *1 105.045,65.52
X$12229 364 48 365 644 645 cell_1rw
* cell instance $12230 m0 *1 105.75,65.52
X$12230 366 48 367 644 645 cell_1rw
* cell instance $12231 m0 *1 106.455,65.52
X$12231 368 48 369 644 645 cell_1rw
* cell instance $12232 m0 *1 107.16,65.52
X$12232 370 48 371 644 645 cell_1rw
* cell instance $12233 m0 *1 107.865,65.52
X$12233 372 48 373 644 645 cell_1rw
* cell instance $12234 m0 *1 108.57,65.52
X$12234 374 48 375 644 645 cell_1rw
* cell instance $12235 m0 *1 109.275,65.52
X$12235 376 48 377 644 645 cell_1rw
* cell instance $12236 m0 *1 109.98,65.52
X$12236 378 48 379 644 645 cell_1rw
* cell instance $12237 m0 *1 110.685,65.52
X$12237 380 48 381 644 645 cell_1rw
* cell instance $12238 m0 *1 111.39,65.52
X$12238 382 48 383 644 645 cell_1rw
* cell instance $12239 m0 *1 112.095,65.52
X$12239 384 48 385 644 645 cell_1rw
* cell instance $12240 m0 *1 112.8,65.52
X$12240 386 48 387 644 645 cell_1rw
* cell instance $12241 m0 *1 113.505,65.52
X$12241 388 48 389 644 645 cell_1rw
* cell instance $12242 m0 *1 114.21,65.52
X$12242 390 48 391 644 645 cell_1rw
* cell instance $12243 m0 *1 114.915,65.52
X$12243 392 48 393 644 645 cell_1rw
* cell instance $12244 m0 *1 115.62,65.52
X$12244 394 48 395 644 645 cell_1rw
* cell instance $12245 m0 *1 116.325,65.52
X$12245 396 48 397 644 645 cell_1rw
* cell instance $12246 m0 *1 117.03,65.52
X$12246 398 48 399 644 645 cell_1rw
* cell instance $12247 m0 *1 117.735,65.52
X$12247 400 48 401 644 645 cell_1rw
* cell instance $12248 m0 *1 118.44,65.52
X$12248 402 48 403 644 645 cell_1rw
* cell instance $12249 m0 *1 119.145,65.52
X$12249 404 48 405 644 645 cell_1rw
* cell instance $12250 m0 *1 119.85,65.52
X$12250 406 48 407 644 645 cell_1rw
* cell instance $12251 m0 *1 120.555,65.52
X$12251 408 48 409 644 645 cell_1rw
* cell instance $12252 m0 *1 121.26,65.52
X$12252 410 48 411 644 645 cell_1rw
* cell instance $12253 m0 *1 121.965,65.52
X$12253 412 48 413 644 645 cell_1rw
* cell instance $12254 m0 *1 122.67,65.52
X$12254 414 48 415 644 645 cell_1rw
* cell instance $12255 m0 *1 123.375,65.52
X$12255 416 48 417 644 645 cell_1rw
* cell instance $12256 m0 *1 124.08,65.52
X$12256 418 48 419 644 645 cell_1rw
* cell instance $12257 m0 *1 124.785,65.52
X$12257 420 48 421 644 645 cell_1rw
* cell instance $12258 m0 *1 125.49,65.52
X$12258 422 48 423 644 645 cell_1rw
* cell instance $12259 m0 *1 126.195,65.52
X$12259 424 48 425 644 645 cell_1rw
* cell instance $12260 m0 *1 126.9,65.52
X$12260 426 48 427 644 645 cell_1rw
* cell instance $12261 m0 *1 127.605,65.52
X$12261 428 48 429 644 645 cell_1rw
* cell instance $12262 m0 *1 128.31,65.52
X$12262 430 48 431 644 645 cell_1rw
* cell instance $12263 m0 *1 129.015,65.52
X$12263 432 48 433 644 645 cell_1rw
* cell instance $12264 m0 *1 129.72,65.52
X$12264 434 48 435 644 645 cell_1rw
* cell instance $12265 m0 *1 130.425,65.52
X$12265 436 48 437 644 645 cell_1rw
* cell instance $12266 m0 *1 131.13,65.52
X$12266 438 48 439 644 645 cell_1rw
* cell instance $12267 m0 *1 131.835,65.52
X$12267 440 48 441 644 645 cell_1rw
* cell instance $12268 m0 *1 132.54,65.52
X$12268 442 48 443 644 645 cell_1rw
* cell instance $12269 m0 *1 133.245,65.52
X$12269 444 48 445 644 645 cell_1rw
* cell instance $12270 m0 *1 133.95,65.52
X$12270 446 48 447 644 645 cell_1rw
* cell instance $12271 m0 *1 134.655,65.52
X$12271 448 48 449 644 645 cell_1rw
* cell instance $12272 m0 *1 135.36,65.52
X$12272 450 48 451 644 645 cell_1rw
* cell instance $12273 m0 *1 136.065,65.52
X$12273 452 48 453 644 645 cell_1rw
* cell instance $12274 m0 *1 136.77,65.52
X$12274 454 48 455 644 645 cell_1rw
* cell instance $12275 m0 *1 137.475,65.52
X$12275 456 48 457 644 645 cell_1rw
* cell instance $12276 m0 *1 138.18,65.52
X$12276 458 48 459 644 645 cell_1rw
* cell instance $12277 m0 *1 138.885,65.52
X$12277 460 48 461 644 645 cell_1rw
* cell instance $12278 m0 *1 139.59,65.52
X$12278 462 48 463 644 645 cell_1rw
* cell instance $12279 m0 *1 140.295,65.52
X$12279 464 48 465 644 645 cell_1rw
* cell instance $12280 m0 *1 141,65.52
X$12280 466 48 467 644 645 cell_1rw
* cell instance $12281 m0 *1 141.705,65.52
X$12281 468 48 469 644 645 cell_1rw
* cell instance $12282 m0 *1 142.41,65.52
X$12282 470 48 471 644 645 cell_1rw
* cell instance $12283 m0 *1 143.115,65.52
X$12283 472 48 473 644 645 cell_1rw
* cell instance $12284 m0 *1 143.82,65.52
X$12284 474 48 475 644 645 cell_1rw
* cell instance $12285 m0 *1 144.525,65.52
X$12285 476 48 477 644 645 cell_1rw
* cell instance $12286 m0 *1 145.23,65.52
X$12286 478 48 479 644 645 cell_1rw
* cell instance $12287 m0 *1 145.935,65.52
X$12287 480 48 481 644 645 cell_1rw
* cell instance $12288 m0 *1 146.64,65.52
X$12288 482 48 483 644 645 cell_1rw
* cell instance $12289 m0 *1 147.345,65.52
X$12289 484 48 485 644 645 cell_1rw
* cell instance $12290 m0 *1 148.05,65.52
X$12290 486 48 487 644 645 cell_1rw
* cell instance $12291 m0 *1 148.755,65.52
X$12291 488 48 489 644 645 cell_1rw
* cell instance $12292 m0 *1 149.46,65.52
X$12292 490 48 491 644 645 cell_1rw
* cell instance $12293 m0 *1 150.165,65.52
X$12293 492 48 493 644 645 cell_1rw
* cell instance $12294 m0 *1 150.87,65.52
X$12294 494 48 495 644 645 cell_1rw
* cell instance $12295 m0 *1 151.575,65.52
X$12295 496 48 497 644 645 cell_1rw
* cell instance $12296 m0 *1 152.28,65.52
X$12296 498 48 499 644 645 cell_1rw
* cell instance $12297 m0 *1 152.985,65.52
X$12297 500 48 501 644 645 cell_1rw
* cell instance $12298 m0 *1 153.69,65.52
X$12298 502 48 503 644 645 cell_1rw
* cell instance $12299 m0 *1 154.395,65.52
X$12299 504 48 505 644 645 cell_1rw
* cell instance $12300 m0 *1 155.1,65.52
X$12300 506 48 507 644 645 cell_1rw
* cell instance $12301 m0 *1 155.805,65.52
X$12301 508 48 509 644 645 cell_1rw
* cell instance $12302 m0 *1 156.51,65.52
X$12302 510 48 511 644 645 cell_1rw
* cell instance $12303 m0 *1 157.215,65.52
X$12303 512 48 513 644 645 cell_1rw
* cell instance $12304 m0 *1 157.92,65.52
X$12304 514 48 515 644 645 cell_1rw
* cell instance $12305 m0 *1 158.625,65.52
X$12305 516 48 517 644 645 cell_1rw
* cell instance $12306 m0 *1 159.33,65.52
X$12306 518 48 519 644 645 cell_1rw
* cell instance $12307 m0 *1 160.035,65.52
X$12307 520 48 521 644 645 cell_1rw
* cell instance $12308 m0 *1 160.74,65.52
X$12308 522 48 523 644 645 cell_1rw
* cell instance $12309 m0 *1 161.445,65.52
X$12309 524 48 525 644 645 cell_1rw
* cell instance $12310 m0 *1 162.15,65.52
X$12310 526 48 527 644 645 cell_1rw
* cell instance $12311 m0 *1 162.855,65.52
X$12311 528 48 529 644 645 cell_1rw
* cell instance $12312 m0 *1 163.56,65.52
X$12312 530 48 531 644 645 cell_1rw
* cell instance $12313 m0 *1 164.265,65.52
X$12313 532 48 533 644 645 cell_1rw
* cell instance $12314 m0 *1 164.97,65.52
X$12314 534 48 535 644 645 cell_1rw
* cell instance $12315 m0 *1 165.675,65.52
X$12315 536 48 537 644 645 cell_1rw
* cell instance $12316 m0 *1 166.38,65.52
X$12316 538 48 539 644 645 cell_1rw
* cell instance $12317 m0 *1 167.085,65.52
X$12317 540 48 541 644 645 cell_1rw
* cell instance $12318 m0 *1 167.79,65.52
X$12318 542 48 543 644 645 cell_1rw
* cell instance $12319 m0 *1 168.495,65.52
X$12319 544 48 545 644 645 cell_1rw
* cell instance $12320 m0 *1 169.2,65.52
X$12320 546 48 547 644 645 cell_1rw
* cell instance $12321 m0 *1 169.905,65.52
X$12321 548 48 549 644 645 cell_1rw
* cell instance $12322 m0 *1 170.61,65.52
X$12322 550 48 551 644 645 cell_1rw
* cell instance $12323 m0 *1 171.315,65.52
X$12323 552 48 553 644 645 cell_1rw
* cell instance $12324 m0 *1 172.02,65.52
X$12324 554 48 555 644 645 cell_1rw
* cell instance $12325 m0 *1 172.725,65.52
X$12325 556 48 557 644 645 cell_1rw
* cell instance $12326 m0 *1 173.43,65.52
X$12326 558 48 559 644 645 cell_1rw
* cell instance $12327 m0 *1 174.135,65.52
X$12327 560 48 561 644 645 cell_1rw
* cell instance $12328 m0 *1 174.84,65.52
X$12328 562 48 563 644 645 cell_1rw
* cell instance $12329 m0 *1 175.545,65.52
X$12329 564 48 565 644 645 cell_1rw
* cell instance $12330 m0 *1 176.25,65.52
X$12330 566 48 567 644 645 cell_1rw
* cell instance $12331 m0 *1 176.955,65.52
X$12331 568 48 569 644 645 cell_1rw
* cell instance $12332 m0 *1 177.66,65.52
X$12332 570 48 571 644 645 cell_1rw
* cell instance $12333 m0 *1 178.365,65.52
X$12333 572 48 573 644 645 cell_1rw
* cell instance $12334 m0 *1 179.07,65.52
X$12334 574 48 575 644 645 cell_1rw
* cell instance $12335 m0 *1 179.775,65.52
X$12335 576 48 577 644 645 cell_1rw
* cell instance $12336 m0 *1 180.48,65.52
X$12336 578 48 579 644 645 cell_1rw
* cell instance $12337 r0 *1 0.705,65.52
X$12337 67 49 68 644 645 cell_1rw
* cell instance $12338 r0 *1 0,65.52
X$12338 65 49 66 644 645 cell_1rw
* cell instance $12339 r0 *1 1.41,65.52
X$12339 69 49 70 644 645 cell_1rw
* cell instance $12340 r0 *1 2.115,65.52
X$12340 71 49 72 644 645 cell_1rw
* cell instance $12341 r0 *1 2.82,65.52
X$12341 73 49 74 644 645 cell_1rw
* cell instance $12342 r0 *1 3.525,65.52
X$12342 75 49 76 644 645 cell_1rw
* cell instance $12343 r0 *1 4.23,65.52
X$12343 77 49 78 644 645 cell_1rw
* cell instance $12344 r0 *1 4.935,65.52
X$12344 79 49 80 644 645 cell_1rw
* cell instance $12345 r0 *1 5.64,65.52
X$12345 81 49 82 644 645 cell_1rw
* cell instance $12346 r0 *1 6.345,65.52
X$12346 83 49 84 644 645 cell_1rw
* cell instance $12347 r0 *1 7.05,65.52
X$12347 85 49 86 644 645 cell_1rw
* cell instance $12348 r0 *1 7.755,65.52
X$12348 87 49 88 644 645 cell_1rw
* cell instance $12349 r0 *1 8.46,65.52
X$12349 89 49 90 644 645 cell_1rw
* cell instance $12350 r0 *1 9.165,65.52
X$12350 91 49 92 644 645 cell_1rw
* cell instance $12351 r0 *1 9.87,65.52
X$12351 93 49 94 644 645 cell_1rw
* cell instance $12352 r0 *1 10.575,65.52
X$12352 95 49 96 644 645 cell_1rw
* cell instance $12353 r0 *1 11.28,65.52
X$12353 97 49 98 644 645 cell_1rw
* cell instance $12354 r0 *1 11.985,65.52
X$12354 99 49 100 644 645 cell_1rw
* cell instance $12355 r0 *1 12.69,65.52
X$12355 101 49 102 644 645 cell_1rw
* cell instance $12356 r0 *1 13.395,65.52
X$12356 103 49 104 644 645 cell_1rw
* cell instance $12357 r0 *1 14.1,65.52
X$12357 105 49 106 644 645 cell_1rw
* cell instance $12358 r0 *1 14.805,65.52
X$12358 107 49 108 644 645 cell_1rw
* cell instance $12359 r0 *1 15.51,65.52
X$12359 109 49 110 644 645 cell_1rw
* cell instance $12360 r0 *1 16.215,65.52
X$12360 111 49 112 644 645 cell_1rw
* cell instance $12361 r0 *1 16.92,65.52
X$12361 113 49 114 644 645 cell_1rw
* cell instance $12362 r0 *1 17.625,65.52
X$12362 115 49 116 644 645 cell_1rw
* cell instance $12363 r0 *1 18.33,65.52
X$12363 117 49 118 644 645 cell_1rw
* cell instance $12364 r0 *1 19.035,65.52
X$12364 119 49 120 644 645 cell_1rw
* cell instance $12365 r0 *1 19.74,65.52
X$12365 121 49 122 644 645 cell_1rw
* cell instance $12366 r0 *1 20.445,65.52
X$12366 123 49 124 644 645 cell_1rw
* cell instance $12367 r0 *1 21.15,65.52
X$12367 125 49 126 644 645 cell_1rw
* cell instance $12368 r0 *1 21.855,65.52
X$12368 127 49 128 644 645 cell_1rw
* cell instance $12369 r0 *1 22.56,65.52
X$12369 129 49 130 644 645 cell_1rw
* cell instance $12370 r0 *1 23.265,65.52
X$12370 131 49 132 644 645 cell_1rw
* cell instance $12371 r0 *1 23.97,65.52
X$12371 133 49 134 644 645 cell_1rw
* cell instance $12372 r0 *1 24.675,65.52
X$12372 135 49 136 644 645 cell_1rw
* cell instance $12373 r0 *1 25.38,65.52
X$12373 137 49 138 644 645 cell_1rw
* cell instance $12374 r0 *1 26.085,65.52
X$12374 139 49 140 644 645 cell_1rw
* cell instance $12375 r0 *1 26.79,65.52
X$12375 141 49 142 644 645 cell_1rw
* cell instance $12376 r0 *1 27.495,65.52
X$12376 143 49 144 644 645 cell_1rw
* cell instance $12377 r0 *1 28.2,65.52
X$12377 145 49 146 644 645 cell_1rw
* cell instance $12378 r0 *1 28.905,65.52
X$12378 147 49 148 644 645 cell_1rw
* cell instance $12379 r0 *1 29.61,65.52
X$12379 149 49 150 644 645 cell_1rw
* cell instance $12380 r0 *1 30.315,65.52
X$12380 151 49 152 644 645 cell_1rw
* cell instance $12381 r0 *1 31.02,65.52
X$12381 153 49 154 644 645 cell_1rw
* cell instance $12382 r0 *1 31.725,65.52
X$12382 155 49 156 644 645 cell_1rw
* cell instance $12383 r0 *1 32.43,65.52
X$12383 157 49 158 644 645 cell_1rw
* cell instance $12384 r0 *1 33.135,65.52
X$12384 159 49 160 644 645 cell_1rw
* cell instance $12385 r0 *1 33.84,65.52
X$12385 161 49 162 644 645 cell_1rw
* cell instance $12386 r0 *1 34.545,65.52
X$12386 163 49 164 644 645 cell_1rw
* cell instance $12387 r0 *1 35.25,65.52
X$12387 165 49 166 644 645 cell_1rw
* cell instance $12388 r0 *1 35.955,65.52
X$12388 167 49 168 644 645 cell_1rw
* cell instance $12389 r0 *1 36.66,65.52
X$12389 169 49 170 644 645 cell_1rw
* cell instance $12390 r0 *1 37.365,65.52
X$12390 171 49 172 644 645 cell_1rw
* cell instance $12391 r0 *1 38.07,65.52
X$12391 173 49 174 644 645 cell_1rw
* cell instance $12392 r0 *1 38.775,65.52
X$12392 175 49 176 644 645 cell_1rw
* cell instance $12393 r0 *1 39.48,65.52
X$12393 177 49 178 644 645 cell_1rw
* cell instance $12394 r0 *1 40.185,65.52
X$12394 179 49 180 644 645 cell_1rw
* cell instance $12395 r0 *1 40.89,65.52
X$12395 181 49 182 644 645 cell_1rw
* cell instance $12396 r0 *1 41.595,65.52
X$12396 183 49 184 644 645 cell_1rw
* cell instance $12397 r0 *1 42.3,65.52
X$12397 185 49 186 644 645 cell_1rw
* cell instance $12398 r0 *1 43.005,65.52
X$12398 187 49 188 644 645 cell_1rw
* cell instance $12399 r0 *1 43.71,65.52
X$12399 189 49 190 644 645 cell_1rw
* cell instance $12400 r0 *1 44.415,65.52
X$12400 191 49 192 644 645 cell_1rw
* cell instance $12401 r0 *1 45.12,65.52
X$12401 193 49 194 644 645 cell_1rw
* cell instance $12402 r0 *1 45.825,65.52
X$12402 195 49 196 644 645 cell_1rw
* cell instance $12403 r0 *1 46.53,65.52
X$12403 197 49 198 644 645 cell_1rw
* cell instance $12404 r0 *1 47.235,65.52
X$12404 199 49 200 644 645 cell_1rw
* cell instance $12405 r0 *1 47.94,65.52
X$12405 201 49 202 644 645 cell_1rw
* cell instance $12406 r0 *1 48.645,65.52
X$12406 203 49 204 644 645 cell_1rw
* cell instance $12407 r0 *1 49.35,65.52
X$12407 205 49 206 644 645 cell_1rw
* cell instance $12408 r0 *1 50.055,65.52
X$12408 207 49 208 644 645 cell_1rw
* cell instance $12409 r0 *1 50.76,65.52
X$12409 209 49 210 644 645 cell_1rw
* cell instance $12410 r0 *1 51.465,65.52
X$12410 211 49 212 644 645 cell_1rw
* cell instance $12411 r0 *1 52.17,65.52
X$12411 213 49 214 644 645 cell_1rw
* cell instance $12412 r0 *1 52.875,65.52
X$12412 215 49 216 644 645 cell_1rw
* cell instance $12413 r0 *1 53.58,65.52
X$12413 217 49 218 644 645 cell_1rw
* cell instance $12414 r0 *1 54.285,65.52
X$12414 219 49 220 644 645 cell_1rw
* cell instance $12415 r0 *1 54.99,65.52
X$12415 221 49 222 644 645 cell_1rw
* cell instance $12416 r0 *1 55.695,65.52
X$12416 223 49 224 644 645 cell_1rw
* cell instance $12417 r0 *1 56.4,65.52
X$12417 225 49 226 644 645 cell_1rw
* cell instance $12418 r0 *1 57.105,65.52
X$12418 227 49 228 644 645 cell_1rw
* cell instance $12419 r0 *1 57.81,65.52
X$12419 229 49 230 644 645 cell_1rw
* cell instance $12420 r0 *1 58.515,65.52
X$12420 231 49 232 644 645 cell_1rw
* cell instance $12421 r0 *1 59.22,65.52
X$12421 233 49 234 644 645 cell_1rw
* cell instance $12422 r0 *1 59.925,65.52
X$12422 235 49 236 644 645 cell_1rw
* cell instance $12423 r0 *1 60.63,65.52
X$12423 237 49 238 644 645 cell_1rw
* cell instance $12424 r0 *1 61.335,65.52
X$12424 239 49 240 644 645 cell_1rw
* cell instance $12425 r0 *1 62.04,65.52
X$12425 241 49 242 644 645 cell_1rw
* cell instance $12426 r0 *1 62.745,65.52
X$12426 243 49 244 644 645 cell_1rw
* cell instance $12427 r0 *1 63.45,65.52
X$12427 245 49 246 644 645 cell_1rw
* cell instance $12428 r0 *1 64.155,65.52
X$12428 247 49 248 644 645 cell_1rw
* cell instance $12429 r0 *1 64.86,65.52
X$12429 249 49 250 644 645 cell_1rw
* cell instance $12430 r0 *1 65.565,65.52
X$12430 251 49 252 644 645 cell_1rw
* cell instance $12431 r0 *1 66.27,65.52
X$12431 253 49 254 644 645 cell_1rw
* cell instance $12432 r0 *1 66.975,65.52
X$12432 255 49 256 644 645 cell_1rw
* cell instance $12433 r0 *1 67.68,65.52
X$12433 257 49 258 644 645 cell_1rw
* cell instance $12434 r0 *1 68.385,65.52
X$12434 259 49 260 644 645 cell_1rw
* cell instance $12435 r0 *1 69.09,65.52
X$12435 261 49 262 644 645 cell_1rw
* cell instance $12436 r0 *1 69.795,65.52
X$12436 263 49 264 644 645 cell_1rw
* cell instance $12437 r0 *1 70.5,65.52
X$12437 265 49 266 644 645 cell_1rw
* cell instance $12438 r0 *1 71.205,65.52
X$12438 267 49 268 644 645 cell_1rw
* cell instance $12439 r0 *1 71.91,65.52
X$12439 269 49 270 644 645 cell_1rw
* cell instance $12440 r0 *1 72.615,65.52
X$12440 271 49 272 644 645 cell_1rw
* cell instance $12441 r0 *1 73.32,65.52
X$12441 273 49 274 644 645 cell_1rw
* cell instance $12442 r0 *1 74.025,65.52
X$12442 275 49 276 644 645 cell_1rw
* cell instance $12443 r0 *1 74.73,65.52
X$12443 277 49 278 644 645 cell_1rw
* cell instance $12444 r0 *1 75.435,65.52
X$12444 279 49 280 644 645 cell_1rw
* cell instance $12445 r0 *1 76.14,65.52
X$12445 281 49 282 644 645 cell_1rw
* cell instance $12446 r0 *1 76.845,65.52
X$12446 283 49 284 644 645 cell_1rw
* cell instance $12447 r0 *1 77.55,65.52
X$12447 285 49 286 644 645 cell_1rw
* cell instance $12448 r0 *1 78.255,65.52
X$12448 287 49 288 644 645 cell_1rw
* cell instance $12449 r0 *1 78.96,65.52
X$12449 289 49 290 644 645 cell_1rw
* cell instance $12450 r0 *1 79.665,65.52
X$12450 291 49 292 644 645 cell_1rw
* cell instance $12451 r0 *1 80.37,65.52
X$12451 293 49 294 644 645 cell_1rw
* cell instance $12452 r0 *1 81.075,65.52
X$12452 295 49 296 644 645 cell_1rw
* cell instance $12453 r0 *1 81.78,65.52
X$12453 297 49 298 644 645 cell_1rw
* cell instance $12454 r0 *1 82.485,65.52
X$12454 299 49 300 644 645 cell_1rw
* cell instance $12455 r0 *1 83.19,65.52
X$12455 301 49 302 644 645 cell_1rw
* cell instance $12456 r0 *1 83.895,65.52
X$12456 303 49 304 644 645 cell_1rw
* cell instance $12457 r0 *1 84.6,65.52
X$12457 305 49 306 644 645 cell_1rw
* cell instance $12458 r0 *1 85.305,65.52
X$12458 307 49 308 644 645 cell_1rw
* cell instance $12459 r0 *1 86.01,65.52
X$12459 309 49 310 644 645 cell_1rw
* cell instance $12460 r0 *1 86.715,65.52
X$12460 311 49 312 644 645 cell_1rw
* cell instance $12461 r0 *1 87.42,65.52
X$12461 313 49 314 644 645 cell_1rw
* cell instance $12462 r0 *1 88.125,65.52
X$12462 315 49 316 644 645 cell_1rw
* cell instance $12463 r0 *1 88.83,65.52
X$12463 317 49 318 644 645 cell_1rw
* cell instance $12464 r0 *1 89.535,65.52
X$12464 319 49 320 644 645 cell_1rw
* cell instance $12465 r0 *1 90.24,65.52
X$12465 321 49 323 644 645 cell_1rw
* cell instance $12466 r0 *1 90.945,65.52
X$12466 324 49 325 644 645 cell_1rw
* cell instance $12467 r0 *1 91.65,65.52
X$12467 326 49 327 644 645 cell_1rw
* cell instance $12468 r0 *1 92.355,65.52
X$12468 328 49 329 644 645 cell_1rw
* cell instance $12469 r0 *1 93.06,65.52
X$12469 330 49 331 644 645 cell_1rw
* cell instance $12470 r0 *1 93.765,65.52
X$12470 332 49 333 644 645 cell_1rw
* cell instance $12471 r0 *1 94.47,65.52
X$12471 334 49 335 644 645 cell_1rw
* cell instance $12472 r0 *1 95.175,65.52
X$12472 336 49 337 644 645 cell_1rw
* cell instance $12473 r0 *1 95.88,65.52
X$12473 338 49 339 644 645 cell_1rw
* cell instance $12474 r0 *1 96.585,65.52
X$12474 340 49 341 644 645 cell_1rw
* cell instance $12475 r0 *1 97.29,65.52
X$12475 342 49 343 644 645 cell_1rw
* cell instance $12476 r0 *1 97.995,65.52
X$12476 344 49 345 644 645 cell_1rw
* cell instance $12477 r0 *1 98.7,65.52
X$12477 346 49 347 644 645 cell_1rw
* cell instance $12478 r0 *1 99.405,65.52
X$12478 348 49 349 644 645 cell_1rw
* cell instance $12479 r0 *1 100.11,65.52
X$12479 350 49 351 644 645 cell_1rw
* cell instance $12480 r0 *1 100.815,65.52
X$12480 352 49 353 644 645 cell_1rw
* cell instance $12481 r0 *1 101.52,65.52
X$12481 354 49 355 644 645 cell_1rw
* cell instance $12482 r0 *1 102.225,65.52
X$12482 356 49 357 644 645 cell_1rw
* cell instance $12483 r0 *1 102.93,65.52
X$12483 358 49 359 644 645 cell_1rw
* cell instance $12484 r0 *1 103.635,65.52
X$12484 360 49 361 644 645 cell_1rw
* cell instance $12485 r0 *1 104.34,65.52
X$12485 362 49 363 644 645 cell_1rw
* cell instance $12486 r0 *1 105.045,65.52
X$12486 364 49 365 644 645 cell_1rw
* cell instance $12487 r0 *1 105.75,65.52
X$12487 366 49 367 644 645 cell_1rw
* cell instance $12488 r0 *1 106.455,65.52
X$12488 368 49 369 644 645 cell_1rw
* cell instance $12489 r0 *1 107.16,65.52
X$12489 370 49 371 644 645 cell_1rw
* cell instance $12490 r0 *1 107.865,65.52
X$12490 372 49 373 644 645 cell_1rw
* cell instance $12491 r0 *1 108.57,65.52
X$12491 374 49 375 644 645 cell_1rw
* cell instance $12492 r0 *1 109.275,65.52
X$12492 376 49 377 644 645 cell_1rw
* cell instance $12493 r0 *1 109.98,65.52
X$12493 378 49 379 644 645 cell_1rw
* cell instance $12494 r0 *1 110.685,65.52
X$12494 380 49 381 644 645 cell_1rw
* cell instance $12495 r0 *1 111.39,65.52
X$12495 382 49 383 644 645 cell_1rw
* cell instance $12496 r0 *1 112.095,65.52
X$12496 384 49 385 644 645 cell_1rw
* cell instance $12497 r0 *1 112.8,65.52
X$12497 386 49 387 644 645 cell_1rw
* cell instance $12498 r0 *1 113.505,65.52
X$12498 388 49 389 644 645 cell_1rw
* cell instance $12499 r0 *1 114.21,65.52
X$12499 390 49 391 644 645 cell_1rw
* cell instance $12500 r0 *1 114.915,65.52
X$12500 392 49 393 644 645 cell_1rw
* cell instance $12501 r0 *1 115.62,65.52
X$12501 394 49 395 644 645 cell_1rw
* cell instance $12502 r0 *1 116.325,65.52
X$12502 396 49 397 644 645 cell_1rw
* cell instance $12503 r0 *1 117.03,65.52
X$12503 398 49 399 644 645 cell_1rw
* cell instance $12504 r0 *1 117.735,65.52
X$12504 400 49 401 644 645 cell_1rw
* cell instance $12505 r0 *1 118.44,65.52
X$12505 402 49 403 644 645 cell_1rw
* cell instance $12506 r0 *1 119.145,65.52
X$12506 404 49 405 644 645 cell_1rw
* cell instance $12507 r0 *1 119.85,65.52
X$12507 406 49 407 644 645 cell_1rw
* cell instance $12508 r0 *1 120.555,65.52
X$12508 408 49 409 644 645 cell_1rw
* cell instance $12509 r0 *1 121.26,65.52
X$12509 410 49 411 644 645 cell_1rw
* cell instance $12510 r0 *1 121.965,65.52
X$12510 412 49 413 644 645 cell_1rw
* cell instance $12511 r0 *1 122.67,65.52
X$12511 414 49 415 644 645 cell_1rw
* cell instance $12512 r0 *1 123.375,65.52
X$12512 416 49 417 644 645 cell_1rw
* cell instance $12513 r0 *1 124.08,65.52
X$12513 418 49 419 644 645 cell_1rw
* cell instance $12514 r0 *1 124.785,65.52
X$12514 420 49 421 644 645 cell_1rw
* cell instance $12515 r0 *1 125.49,65.52
X$12515 422 49 423 644 645 cell_1rw
* cell instance $12516 r0 *1 126.195,65.52
X$12516 424 49 425 644 645 cell_1rw
* cell instance $12517 r0 *1 126.9,65.52
X$12517 426 49 427 644 645 cell_1rw
* cell instance $12518 r0 *1 127.605,65.52
X$12518 428 49 429 644 645 cell_1rw
* cell instance $12519 r0 *1 128.31,65.52
X$12519 430 49 431 644 645 cell_1rw
* cell instance $12520 r0 *1 129.015,65.52
X$12520 432 49 433 644 645 cell_1rw
* cell instance $12521 r0 *1 129.72,65.52
X$12521 434 49 435 644 645 cell_1rw
* cell instance $12522 r0 *1 130.425,65.52
X$12522 436 49 437 644 645 cell_1rw
* cell instance $12523 r0 *1 131.13,65.52
X$12523 438 49 439 644 645 cell_1rw
* cell instance $12524 r0 *1 131.835,65.52
X$12524 440 49 441 644 645 cell_1rw
* cell instance $12525 r0 *1 132.54,65.52
X$12525 442 49 443 644 645 cell_1rw
* cell instance $12526 r0 *1 133.245,65.52
X$12526 444 49 445 644 645 cell_1rw
* cell instance $12527 r0 *1 133.95,65.52
X$12527 446 49 447 644 645 cell_1rw
* cell instance $12528 r0 *1 134.655,65.52
X$12528 448 49 449 644 645 cell_1rw
* cell instance $12529 r0 *1 135.36,65.52
X$12529 450 49 451 644 645 cell_1rw
* cell instance $12530 r0 *1 136.065,65.52
X$12530 452 49 453 644 645 cell_1rw
* cell instance $12531 r0 *1 136.77,65.52
X$12531 454 49 455 644 645 cell_1rw
* cell instance $12532 r0 *1 137.475,65.52
X$12532 456 49 457 644 645 cell_1rw
* cell instance $12533 r0 *1 138.18,65.52
X$12533 458 49 459 644 645 cell_1rw
* cell instance $12534 r0 *1 138.885,65.52
X$12534 460 49 461 644 645 cell_1rw
* cell instance $12535 r0 *1 139.59,65.52
X$12535 462 49 463 644 645 cell_1rw
* cell instance $12536 r0 *1 140.295,65.52
X$12536 464 49 465 644 645 cell_1rw
* cell instance $12537 r0 *1 141,65.52
X$12537 466 49 467 644 645 cell_1rw
* cell instance $12538 r0 *1 141.705,65.52
X$12538 468 49 469 644 645 cell_1rw
* cell instance $12539 r0 *1 142.41,65.52
X$12539 470 49 471 644 645 cell_1rw
* cell instance $12540 r0 *1 143.115,65.52
X$12540 472 49 473 644 645 cell_1rw
* cell instance $12541 r0 *1 143.82,65.52
X$12541 474 49 475 644 645 cell_1rw
* cell instance $12542 r0 *1 144.525,65.52
X$12542 476 49 477 644 645 cell_1rw
* cell instance $12543 r0 *1 145.23,65.52
X$12543 478 49 479 644 645 cell_1rw
* cell instance $12544 r0 *1 145.935,65.52
X$12544 480 49 481 644 645 cell_1rw
* cell instance $12545 r0 *1 146.64,65.52
X$12545 482 49 483 644 645 cell_1rw
* cell instance $12546 r0 *1 147.345,65.52
X$12546 484 49 485 644 645 cell_1rw
* cell instance $12547 r0 *1 148.05,65.52
X$12547 486 49 487 644 645 cell_1rw
* cell instance $12548 r0 *1 148.755,65.52
X$12548 488 49 489 644 645 cell_1rw
* cell instance $12549 r0 *1 149.46,65.52
X$12549 490 49 491 644 645 cell_1rw
* cell instance $12550 r0 *1 150.165,65.52
X$12550 492 49 493 644 645 cell_1rw
* cell instance $12551 r0 *1 150.87,65.52
X$12551 494 49 495 644 645 cell_1rw
* cell instance $12552 r0 *1 151.575,65.52
X$12552 496 49 497 644 645 cell_1rw
* cell instance $12553 r0 *1 152.28,65.52
X$12553 498 49 499 644 645 cell_1rw
* cell instance $12554 r0 *1 152.985,65.52
X$12554 500 49 501 644 645 cell_1rw
* cell instance $12555 r0 *1 153.69,65.52
X$12555 502 49 503 644 645 cell_1rw
* cell instance $12556 r0 *1 154.395,65.52
X$12556 504 49 505 644 645 cell_1rw
* cell instance $12557 r0 *1 155.1,65.52
X$12557 506 49 507 644 645 cell_1rw
* cell instance $12558 r0 *1 155.805,65.52
X$12558 508 49 509 644 645 cell_1rw
* cell instance $12559 r0 *1 156.51,65.52
X$12559 510 49 511 644 645 cell_1rw
* cell instance $12560 r0 *1 157.215,65.52
X$12560 512 49 513 644 645 cell_1rw
* cell instance $12561 r0 *1 157.92,65.52
X$12561 514 49 515 644 645 cell_1rw
* cell instance $12562 r0 *1 158.625,65.52
X$12562 516 49 517 644 645 cell_1rw
* cell instance $12563 r0 *1 159.33,65.52
X$12563 518 49 519 644 645 cell_1rw
* cell instance $12564 r0 *1 160.035,65.52
X$12564 520 49 521 644 645 cell_1rw
* cell instance $12565 r0 *1 160.74,65.52
X$12565 522 49 523 644 645 cell_1rw
* cell instance $12566 r0 *1 161.445,65.52
X$12566 524 49 525 644 645 cell_1rw
* cell instance $12567 r0 *1 162.15,65.52
X$12567 526 49 527 644 645 cell_1rw
* cell instance $12568 r0 *1 162.855,65.52
X$12568 528 49 529 644 645 cell_1rw
* cell instance $12569 r0 *1 163.56,65.52
X$12569 530 49 531 644 645 cell_1rw
* cell instance $12570 r0 *1 164.265,65.52
X$12570 532 49 533 644 645 cell_1rw
* cell instance $12571 r0 *1 164.97,65.52
X$12571 534 49 535 644 645 cell_1rw
* cell instance $12572 r0 *1 165.675,65.52
X$12572 536 49 537 644 645 cell_1rw
* cell instance $12573 r0 *1 166.38,65.52
X$12573 538 49 539 644 645 cell_1rw
* cell instance $12574 r0 *1 167.085,65.52
X$12574 540 49 541 644 645 cell_1rw
* cell instance $12575 r0 *1 167.79,65.52
X$12575 542 49 543 644 645 cell_1rw
* cell instance $12576 r0 *1 168.495,65.52
X$12576 544 49 545 644 645 cell_1rw
* cell instance $12577 r0 *1 169.2,65.52
X$12577 546 49 547 644 645 cell_1rw
* cell instance $12578 r0 *1 169.905,65.52
X$12578 548 49 549 644 645 cell_1rw
* cell instance $12579 r0 *1 170.61,65.52
X$12579 550 49 551 644 645 cell_1rw
* cell instance $12580 r0 *1 171.315,65.52
X$12580 552 49 553 644 645 cell_1rw
* cell instance $12581 r0 *1 172.02,65.52
X$12581 554 49 555 644 645 cell_1rw
* cell instance $12582 r0 *1 172.725,65.52
X$12582 556 49 557 644 645 cell_1rw
* cell instance $12583 r0 *1 173.43,65.52
X$12583 558 49 559 644 645 cell_1rw
* cell instance $12584 r0 *1 174.135,65.52
X$12584 560 49 561 644 645 cell_1rw
* cell instance $12585 r0 *1 174.84,65.52
X$12585 562 49 563 644 645 cell_1rw
* cell instance $12586 r0 *1 175.545,65.52
X$12586 564 49 565 644 645 cell_1rw
* cell instance $12587 r0 *1 176.25,65.52
X$12587 566 49 567 644 645 cell_1rw
* cell instance $12588 r0 *1 176.955,65.52
X$12588 568 49 569 644 645 cell_1rw
* cell instance $12589 r0 *1 177.66,65.52
X$12589 570 49 571 644 645 cell_1rw
* cell instance $12590 r0 *1 178.365,65.52
X$12590 572 49 573 644 645 cell_1rw
* cell instance $12591 r0 *1 179.07,65.52
X$12591 574 49 575 644 645 cell_1rw
* cell instance $12592 r0 *1 179.775,65.52
X$12592 576 49 577 644 645 cell_1rw
* cell instance $12593 r0 *1 180.48,65.52
X$12593 578 49 579 644 645 cell_1rw
* cell instance $12594 m0 *1 0.705,68.25
X$12594 67 50 68 644 645 cell_1rw
* cell instance $12595 m0 *1 0,68.25
X$12595 65 50 66 644 645 cell_1rw
* cell instance $12596 m0 *1 1.41,68.25
X$12596 69 50 70 644 645 cell_1rw
* cell instance $12597 m0 *1 2.115,68.25
X$12597 71 50 72 644 645 cell_1rw
* cell instance $12598 m0 *1 2.82,68.25
X$12598 73 50 74 644 645 cell_1rw
* cell instance $12599 m0 *1 3.525,68.25
X$12599 75 50 76 644 645 cell_1rw
* cell instance $12600 m0 *1 4.23,68.25
X$12600 77 50 78 644 645 cell_1rw
* cell instance $12601 m0 *1 4.935,68.25
X$12601 79 50 80 644 645 cell_1rw
* cell instance $12602 m0 *1 5.64,68.25
X$12602 81 50 82 644 645 cell_1rw
* cell instance $12603 m0 *1 6.345,68.25
X$12603 83 50 84 644 645 cell_1rw
* cell instance $12604 m0 *1 7.05,68.25
X$12604 85 50 86 644 645 cell_1rw
* cell instance $12605 m0 *1 7.755,68.25
X$12605 87 50 88 644 645 cell_1rw
* cell instance $12606 m0 *1 8.46,68.25
X$12606 89 50 90 644 645 cell_1rw
* cell instance $12607 m0 *1 9.165,68.25
X$12607 91 50 92 644 645 cell_1rw
* cell instance $12608 m0 *1 9.87,68.25
X$12608 93 50 94 644 645 cell_1rw
* cell instance $12609 m0 *1 10.575,68.25
X$12609 95 50 96 644 645 cell_1rw
* cell instance $12610 m0 *1 11.28,68.25
X$12610 97 50 98 644 645 cell_1rw
* cell instance $12611 m0 *1 11.985,68.25
X$12611 99 50 100 644 645 cell_1rw
* cell instance $12612 m0 *1 12.69,68.25
X$12612 101 50 102 644 645 cell_1rw
* cell instance $12613 m0 *1 13.395,68.25
X$12613 103 50 104 644 645 cell_1rw
* cell instance $12614 m0 *1 14.1,68.25
X$12614 105 50 106 644 645 cell_1rw
* cell instance $12615 m0 *1 14.805,68.25
X$12615 107 50 108 644 645 cell_1rw
* cell instance $12616 m0 *1 15.51,68.25
X$12616 109 50 110 644 645 cell_1rw
* cell instance $12617 m0 *1 16.215,68.25
X$12617 111 50 112 644 645 cell_1rw
* cell instance $12618 m0 *1 16.92,68.25
X$12618 113 50 114 644 645 cell_1rw
* cell instance $12619 m0 *1 17.625,68.25
X$12619 115 50 116 644 645 cell_1rw
* cell instance $12620 m0 *1 18.33,68.25
X$12620 117 50 118 644 645 cell_1rw
* cell instance $12621 m0 *1 19.035,68.25
X$12621 119 50 120 644 645 cell_1rw
* cell instance $12622 m0 *1 19.74,68.25
X$12622 121 50 122 644 645 cell_1rw
* cell instance $12623 m0 *1 20.445,68.25
X$12623 123 50 124 644 645 cell_1rw
* cell instance $12624 m0 *1 21.15,68.25
X$12624 125 50 126 644 645 cell_1rw
* cell instance $12625 m0 *1 21.855,68.25
X$12625 127 50 128 644 645 cell_1rw
* cell instance $12626 m0 *1 22.56,68.25
X$12626 129 50 130 644 645 cell_1rw
* cell instance $12627 m0 *1 23.265,68.25
X$12627 131 50 132 644 645 cell_1rw
* cell instance $12628 m0 *1 23.97,68.25
X$12628 133 50 134 644 645 cell_1rw
* cell instance $12629 m0 *1 24.675,68.25
X$12629 135 50 136 644 645 cell_1rw
* cell instance $12630 m0 *1 25.38,68.25
X$12630 137 50 138 644 645 cell_1rw
* cell instance $12631 m0 *1 26.085,68.25
X$12631 139 50 140 644 645 cell_1rw
* cell instance $12632 m0 *1 26.79,68.25
X$12632 141 50 142 644 645 cell_1rw
* cell instance $12633 m0 *1 27.495,68.25
X$12633 143 50 144 644 645 cell_1rw
* cell instance $12634 m0 *1 28.2,68.25
X$12634 145 50 146 644 645 cell_1rw
* cell instance $12635 m0 *1 28.905,68.25
X$12635 147 50 148 644 645 cell_1rw
* cell instance $12636 m0 *1 29.61,68.25
X$12636 149 50 150 644 645 cell_1rw
* cell instance $12637 m0 *1 30.315,68.25
X$12637 151 50 152 644 645 cell_1rw
* cell instance $12638 m0 *1 31.02,68.25
X$12638 153 50 154 644 645 cell_1rw
* cell instance $12639 m0 *1 31.725,68.25
X$12639 155 50 156 644 645 cell_1rw
* cell instance $12640 m0 *1 32.43,68.25
X$12640 157 50 158 644 645 cell_1rw
* cell instance $12641 m0 *1 33.135,68.25
X$12641 159 50 160 644 645 cell_1rw
* cell instance $12642 m0 *1 33.84,68.25
X$12642 161 50 162 644 645 cell_1rw
* cell instance $12643 m0 *1 34.545,68.25
X$12643 163 50 164 644 645 cell_1rw
* cell instance $12644 m0 *1 35.25,68.25
X$12644 165 50 166 644 645 cell_1rw
* cell instance $12645 m0 *1 35.955,68.25
X$12645 167 50 168 644 645 cell_1rw
* cell instance $12646 m0 *1 36.66,68.25
X$12646 169 50 170 644 645 cell_1rw
* cell instance $12647 m0 *1 37.365,68.25
X$12647 171 50 172 644 645 cell_1rw
* cell instance $12648 m0 *1 38.07,68.25
X$12648 173 50 174 644 645 cell_1rw
* cell instance $12649 m0 *1 38.775,68.25
X$12649 175 50 176 644 645 cell_1rw
* cell instance $12650 m0 *1 39.48,68.25
X$12650 177 50 178 644 645 cell_1rw
* cell instance $12651 m0 *1 40.185,68.25
X$12651 179 50 180 644 645 cell_1rw
* cell instance $12652 m0 *1 40.89,68.25
X$12652 181 50 182 644 645 cell_1rw
* cell instance $12653 m0 *1 41.595,68.25
X$12653 183 50 184 644 645 cell_1rw
* cell instance $12654 m0 *1 42.3,68.25
X$12654 185 50 186 644 645 cell_1rw
* cell instance $12655 m0 *1 43.005,68.25
X$12655 187 50 188 644 645 cell_1rw
* cell instance $12656 m0 *1 43.71,68.25
X$12656 189 50 190 644 645 cell_1rw
* cell instance $12657 m0 *1 44.415,68.25
X$12657 191 50 192 644 645 cell_1rw
* cell instance $12658 m0 *1 45.12,68.25
X$12658 193 50 194 644 645 cell_1rw
* cell instance $12659 m0 *1 45.825,68.25
X$12659 195 50 196 644 645 cell_1rw
* cell instance $12660 m0 *1 46.53,68.25
X$12660 197 50 198 644 645 cell_1rw
* cell instance $12661 m0 *1 47.235,68.25
X$12661 199 50 200 644 645 cell_1rw
* cell instance $12662 m0 *1 47.94,68.25
X$12662 201 50 202 644 645 cell_1rw
* cell instance $12663 m0 *1 48.645,68.25
X$12663 203 50 204 644 645 cell_1rw
* cell instance $12664 m0 *1 49.35,68.25
X$12664 205 50 206 644 645 cell_1rw
* cell instance $12665 m0 *1 50.055,68.25
X$12665 207 50 208 644 645 cell_1rw
* cell instance $12666 m0 *1 50.76,68.25
X$12666 209 50 210 644 645 cell_1rw
* cell instance $12667 m0 *1 51.465,68.25
X$12667 211 50 212 644 645 cell_1rw
* cell instance $12668 m0 *1 52.17,68.25
X$12668 213 50 214 644 645 cell_1rw
* cell instance $12669 m0 *1 52.875,68.25
X$12669 215 50 216 644 645 cell_1rw
* cell instance $12670 m0 *1 53.58,68.25
X$12670 217 50 218 644 645 cell_1rw
* cell instance $12671 m0 *1 54.285,68.25
X$12671 219 50 220 644 645 cell_1rw
* cell instance $12672 m0 *1 54.99,68.25
X$12672 221 50 222 644 645 cell_1rw
* cell instance $12673 m0 *1 55.695,68.25
X$12673 223 50 224 644 645 cell_1rw
* cell instance $12674 m0 *1 56.4,68.25
X$12674 225 50 226 644 645 cell_1rw
* cell instance $12675 m0 *1 57.105,68.25
X$12675 227 50 228 644 645 cell_1rw
* cell instance $12676 m0 *1 57.81,68.25
X$12676 229 50 230 644 645 cell_1rw
* cell instance $12677 m0 *1 58.515,68.25
X$12677 231 50 232 644 645 cell_1rw
* cell instance $12678 m0 *1 59.22,68.25
X$12678 233 50 234 644 645 cell_1rw
* cell instance $12679 m0 *1 59.925,68.25
X$12679 235 50 236 644 645 cell_1rw
* cell instance $12680 m0 *1 60.63,68.25
X$12680 237 50 238 644 645 cell_1rw
* cell instance $12681 m0 *1 61.335,68.25
X$12681 239 50 240 644 645 cell_1rw
* cell instance $12682 m0 *1 62.04,68.25
X$12682 241 50 242 644 645 cell_1rw
* cell instance $12683 m0 *1 62.745,68.25
X$12683 243 50 244 644 645 cell_1rw
* cell instance $12684 m0 *1 63.45,68.25
X$12684 245 50 246 644 645 cell_1rw
* cell instance $12685 m0 *1 64.155,68.25
X$12685 247 50 248 644 645 cell_1rw
* cell instance $12686 m0 *1 64.86,68.25
X$12686 249 50 250 644 645 cell_1rw
* cell instance $12687 m0 *1 65.565,68.25
X$12687 251 50 252 644 645 cell_1rw
* cell instance $12688 m0 *1 66.27,68.25
X$12688 253 50 254 644 645 cell_1rw
* cell instance $12689 m0 *1 66.975,68.25
X$12689 255 50 256 644 645 cell_1rw
* cell instance $12690 m0 *1 67.68,68.25
X$12690 257 50 258 644 645 cell_1rw
* cell instance $12691 m0 *1 68.385,68.25
X$12691 259 50 260 644 645 cell_1rw
* cell instance $12692 m0 *1 69.09,68.25
X$12692 261 50 262 644 645 cell_1rw
* cell instance $12693 m0 *1 69.795,68.25
X$12693 263 50 264 644 645 cell_1rw
* cell instance $12694 m0 *1 70.5,68.25
X$12694 265 50 266 644 645 cell_1rw
* cell instance $12695 m0 *1 71.205,68.25
X$12695 267 50 268 644 645 cell_1rw
* cell instance $12696 m0 *1 71.91,68.25
X$12696 269 50 270 644 645 cell_1rw
* cell instance $12697 m0 *1 72.615,68.25
X$12697 271 50 272 644 645 cell_1rw
* cell instance $12698 m0 *1 73.32,68.25
X$12698 273 50 274 644 645 cell_1rw
* cell instance $12699 m0 *1 74.025,68.25
X$12699 275 50 276 644 645 cell_1rw
* cell instance $12700 m0 *1 74.73,68.25
X$12700 277 50 278 644 645 cell_1rw
* cell instance $12701 m0 *1 75.435,68.25
X$12701 279 50 280 644 645 cell_1rw
* cell instance $12702 m0 *1 76.14,68.25
X$12702 281 50 282 644 645 cell_1rw
* cell instance $12703 m0 *1 76.845,68.25
X$12703 283 50 284 644 645 cell_1rw
* cell instance $12704 m0 *1 77.55,68.25
X$12704 285 50 286 644 645 cell_1rw
* cell instance $12705 m0 *1 78.255,68.25
X$12705 287 50 288 644 645 cell_1rw
* cell instance $12706 m0 *1 78.96,68.25
X$12706 289 50 290 644 645 cell_1rw
* cell instance $12707 m0 *1 79.665,68.25
X$12707 291 50 292 644 645 cell_1rw
* cell instance $12708 m0 *1 80.37,68.25
X$12708 293 50 294 644 645 cell_1rw
* cell instance $12709 m0 *1 81.075,68.25
X$12709 295 50 296 644 645 cell_1rw
* cell instance $12710 m0 *1 81.78,68.25
X$12710 297 50 298 644 645 cell_1rw
* cell instance $12711 m0 *1 82.485,68.25
X$12711 299 50 300 644 645 cell_1rw
* cell instance $12712 m0 *1 83.19,68.25
X$12712 301 50 302 644 645 cell_1rw
* cell instance $12713 m0 *1 83.895,68.25
X$12713 303 50 304 644 645 cell_1rw
* cell instance $12714 m0 *1 84.6,68.25
X$12714 305 50 306 644 645 cell_1rw
* cell instance $12715 m0 *1 85.305,68.25
X$12715 307 50 308 644 645 cell_1rw
* cell instance $12716 m0 *1 86.01,68.25
X$12716 309 50 310 644 645 cell_1rw
* cell instance $12717 m0 *1 86.715,68.25
X$12717 311 50 312 644 645 cell_1rw
* cell instance $12718 m0 *1 87.42,68.25
X$12718 313 50 314 644 645 cell_1rw
* cell instance $12719 m0 *1 88.125,68.25
X$12719 315 50 316 644 645 cell_1rw
* cell instance $12720 m0 *1 88.83,68.25
X$12720 317 50 318 644 645 cell_1rw
* cell instance $12721 m0 *1 89.535,68.25
X$12721 319 50 320 644 645 cell_1rw
* cell instance $12722 m0 *1 90.24,68.25
X$12722 321 50 323 644 645 cell_1rw
* cell instance $12723 m0 *1 90.945,68.25
X$12723 324 50 325 644 645 cell_1rw
* cell instance $12724 m0 *1 91.65,68.25
X$12724 326 50 327 644 645 cell_1rw
* cell instance $12725 m0 *1 92.355,68.25
X$12725 328 50 329 644 645 cell_1rw
* cell instance $12726 m0 *1 93.06,68.25
X$12726 330 50 331 644 645 cell_1rw
* cell instance $12727 m0 *1 93.765,68.25
X$12727 332 50 333 644 645 cell_1rw
* cell instance $12728 m0 *1 94.47,68.25
X$12728 334 50 335 644 645 cell_1rw
* cell instance $12729 m0 *1 95.175,68.25
X$12729 336 50 337 644 645 cell_1rw
* cell instance $12730 m0 *1 95.88,68.25
X$12730 338 50 339 644 645 cell_1rw
* cell instance $12731 m0 *1 96.585,68.25
X$12731 340 50 341 644 645 cell_1rw
* cell instance $12732 m0 *1 97.29,68.25
X$12732 342 50 343 644 645 cell_1rw
* cell instance $12733 m0 *1 97.995,68.25
X$12733 344 50 345 644 645 cell_1rw
* cell instance $12734 m0 *1 98.7,68.25
X$12734 346 50 347 644 645 cell_1rw
* cell instance $12735 m0 *1 99.405,68.25
X$12735 348 50 349 644 645 cell_1rw
* cell instance $12736 m0 *1 100.11,68.25
X$12736 350 50 351 644 645 cell_1rw
* cell instance $12737 m0 *1 100.815,68.25
X$12737 352 50 353 644 645 cell_1rw
* cell instance $12738 m0 *1 101.52,68.25
X$12738 354 50 355 644 645 cell_1rw
* cell instance $12739 m0 *1 102.225,68.25
X$12739 356 50 357 644 645 cell_1rw
* cell instance $12740 m0 *1 102.93,68.25
X$12740 358 50 359 644 645 cell_1rw
* cell instance $12741 m0 *1 103.635,68.25
X$12741 360 50 361 644 645 cell_1rw
* cell instance $12742 m0 *1 104.34,68.25
X$12742 362 50 363 644 645 cell_1rw
* cell instance $12743 m0 *1 105.045,68.25
X$12743 364 50 365 644 645 cell_1rw
* cell instance $12744 m0 *1 105.75,68.25
X$12744 366 50 367 644 645 cell_1rw
* cell instance $12745 m0 *1 106.455,68.25
X$12745 368 50 369 644 645 cell_1rw
* cell instance $12746 m0 *1 107.16,68.25
X$12746 370 50 371 644 645 cell_1rw
* cell instance $12747 m0 *1 107.865,68.25
X$12747 372 50 373 644 645 cell_1rw
* cell instance $12748 m0 *1 108.57,68.25
X$12748 374 50 375 644 645 cell_1rw
* cell instance $12749 m0 *1 109.275,68.25
X$12749 376 50 377 644 645 cell_1rw
* cell instance $12750 m0 *1 109.98,68.25
X$12750 378 50 379 644 645 cell_1rw
* cell instance $12751 m0 *1 110.685,68.25
X$12751 380 50 381 644 645 cell_1rw
* cell instance $12752 m0 *1 111.39,68.25
X$12752 382 50 383 644 645 cell_1rw
* cell instance $12753 m0 *1 112.095,68.25
X$12753 384 50 385 644 645 cell_1rw
* cell instance $12754 m0 *1 112.8,68.25
X$12754 386 50 387 644 645 cell_1rw
* cell instance $12755 m0 *1 113.505,68.25
X$12755 388 50 389 644 645 cell_1rw
* cell instance $12756 m0 *1 114.21,68.25
X$12756 390 50 391 644 645 cell_1rw
* cell instance $12757 m0 *1 114.915,68.25
X$12757 392 50 393 644 645 cell_1rw
* cell instance $12758 m0 *1 115.62,68.25
X$12758 394 50 395 644 645 cell_1rw
* cell instance $12759 m0 *1 116.325,68.25
X$12759 396 50 397 644 645 cell_1rw
* cell instance $12760 m0 *1 117.03,68.25
X$12760 398 50 399 644 645 cell_1rw
* cell instance $12761 m0 *1 117.735,68.25
X$12761 400 50 401 644 645 cell_1rw
* cell instance $12762 m0 *1 118.44,68.25
X$12762 402 50 403 644 645 cell_1rw
* cell instance $12763 m0 *1 119.145,68.25
X$12763 404 50 405 644 645 cell_1rw
* cell instance $12764 m0 *1 119.85,68.25
X$12764 406 50 407 644 645 cell_1rw
* cell instance $12765 m0 *1 120.555,68.25
X$12765 408 50 409 644 645 cell_1rw
* cell instance $12766 m0 *1 121.26,68.25
X$12766 410 50 411 644 645 cell_1rw
* cell instance $12767 m0 *1 121.965,68.25
X$12767 412 50 413 644 645 cell_1rw
* cell instance $12768 m0 *1 122.67,68.25
X$12768 414 50 415 644 645 cell_1rw
* cell instance $12769 m0 *1 123.375,68.25
X$12769 416 50 417 644 645 cell_1rw
* cell instance $12770 m0 *1 124.08,68.25
X$12770 418 50 419 644 645 cell_1rw
* cell instance $12771 m0 *1 124.785,68.25
X$12771 420 50 421 644 645 cell_1rw
* cell instance $12772 m0 *1 125.49,68.25
X$12772 422 50 423 644 645 cell_1rw
* cell instance $12773 m0 *1 126.195,68.25
X$12773 424 50 425 644 645 cell_1rw
* cell instance $12774 m0 *1 126.9,68.25
X$12774 426 50 427 644 645 cell_1rw
* cell instance $12775 m0 *1 127.605,68.25
X$12775 428 50 429 644 645 cell_1rw
* cell instance $12776 m0 *1 128.31,68.25
X$12776 430 50 431 644 645 cell_1rw
* cell instance $12777 m0 *1 129.015,68.25
X$12777 432 50 433 644 645 cell_1rw
* cell instance $12778 m0 *1 129.72,68.25
X$12778 434 50 435 644 645 cell_1rw
* cell instance $12779 m0 *1 130.425,68.25
X$12779 436 50 437 644 645 cell_1rw
* cell instance $12780 m0 *1 131.13,68.25
X$12780 438 50 439 644 645 cell_1rw
* cell instance $12781 m0 *1 131.835,68.25
X$12781 440 50 441 644 645 cell_1rw
* cell instance $12782 m0 *1 132.54,68.25
X$12782 442 50 443 644 645 cell_1rw
* cell instance $12783 m0 *1 133.245,68.25
X$12783 444 50 445 644 645 cell_1rw
* cell instance $12784 m0 *1 133.95,68.25
X$12784 446 50 447 644 645 cell_1rw
* cell instance $12785 m0 *1 134.655,68.25
X$12785 448 50 449 644 645 cell_1rw
* cell instance $12786 m0 *1 135.36,68.25
X$12786 450 50 451 644 645 cell_1rw
* cell instance $12787 m0 *1 136.065,68.25
X$12787 452 50 453 644 645 cell_1rw
* cell instance $12788 m0 *1 136.77,68.25
X$12788 454 50 455 644 645 cell_1rw
* cell instance $12789 m0 *1 137.475,68.25
X$12789 456 50 457 644 645 cell_1rw
* cell instance $12790 m0 *1 138.18,68.25
X$12790 458 50 459 644 645 cell_1rw
* cell instance $12791 m0 *1 138.885,68.25
X$12791 460 50 461 644 645 cell_1rw
* cell instance $12792 m0 *1 139.59,68.25
X$12792 462 50 463 644 645 cell_1rw
* cell instance $12793 m0 *1 140.295,68.25
X$12793 464 50 465 644 645 cell_1rw
* cell instance $12794 m0 *1 141,68.25
X$12794 466 50 467 644 645 cell_1rw
* cell instance $12795 m0 *1 141.705,68.25
X$12795 468 50 469 644 645 cell_1rw
* cell instance $12796 m0 *1 142.41,68.25
X$12796 470 50 471 644 645 cell_1rw
* cell instance $12797 m0 *1 143.115,68.25
X$12797 472 50 473 644 645 cell_1rw
* cell instance $12798 m0 *1 143.82,68.25
X$12798 474 50 475 644 645 cell_1rw
* cell instance $12799 m0 *1 144.525,68.25
X$12799 476 50 477 644 645 cell_1rw
* cell instance $12800 m0 *1 145.23,68.25
X$12800 478 50 479 644 645 cell_1rw
* cell instance $12801 m0 *1 145.935,68.25
X$12801 480 50 481 644 645 cell_1rw
* cell instance $12802 m0 *1 146.64,68.25
X$12802 482 50 483 644 645 cell_1rw
* cell instance $12803 m0 *1 147.345,68.25
X$12803 484 50 485 644 645 cell_1rw
* cell instance $12804 m0 *1 148.05,68.25
X$12804 486 50 487 644 645 cell_1rw
* cell instance $12805 m0 *1 148.755,68.25
X$12805 488 50 489 644 645 cell_1rw
* cell instance $12806 m0 *1 149.46,68.25
X$12806 490 50 491 644 645 cell_1rw
* cell instance $12807 m0 *1 150.165,68.25
X$12807 492 50 493 644 645 cell_1rw
* cell instance $12808 m0 *1 150.87,68.25
X$12808 494 50 495 644 645 cell_1rw
* cell instance $12809 m0 *1 151.575,68.25
X$12809 496 50 497 644 645 cell_1rw
* cell instance $12810 m0 *1 152.28,68.25
X$12810 498 50 499 644 645 cell_1rw
* cell instance $12811 m0 *1 152.985,68.25
X$12811 500 50 501 644 645 cell_1rw
* cell instance $12812 m0 *1 153.69,68.25
X$12812 502 50 503 644 645 cell_1rw
* cell instance $12813 m0 *1 154.395,68.25
X$12813 504 50 505 644 645 cell_1rw
* cell instance $12814 m0 *1 155.1,68.25
X$12814 506 50 507 644 645 cell_1rw
* cell instance $12815 m0 *1 155.805,68.25
X$12815 508 50 509 644 645 cell_1rw
* cell instance $12816 m0 *1 156.51,68.25
X$12816 510 50 511 644 645 cell_1rw
* cell instance $12817 m0 *1 157.215,68.25
X$12817 512 50 513 644 645 cell_1rw
* cell instance $12818 m0 *1 157.92,68.25
X$12818 514 50 515 644 645 cell_1rw
* cell instance $12819 m0 *1 158.625,68.25
X$12819 516 50 517 644 645 cell_1rw
* cell instance $12820 m0 *1 159.33,68.25
X$12820 518 50 519 644 645 cell_1rw
* cell instance $12821 m0 *1 160.035,68.25
X$12821 520 50 521 644 645 cell_1rw
* cell instance $12822 m0 *1 160.74,68.25
X$12822 522 50 523 644 645 cell_1rw
* cell instance $12823 m0 *1 161.445,68.25
X$12823 524 50 525 644 645 cell_1rw
* cell instance $12824 m0 *1 162.15,68.25
X$12824 526 50 527 644 645 cell_1rw
* cell instance $12825 m0 *1 162.855,68.25
X$12825 528 50 529 644 645 cell_1rw
* cell instance $12826 m0 *1 163.56,68.25
X$12826 530 50 531 644 645 cell_1rw
* cell instance $12827 m0 *1 164.265,68.25
X$12827 532 50 533 644 645 cell_1rw
* cell instance $12828 m0 *1 164.97,68.25
X$12828 534 50 535 644 645 cell_1rw
* cell instance $12829 m0 *1 165.675,68.25
X$12829 536 50 537 644 645 cell_1rw
* cell instance $12830 m0 *1 166.38,68.25
X$12830 538 50 539 644 645 cell_1rw
* cell instance $12831 m0 *1 167.085,68.25
X$12831 540 50 541 644 645 cell_1rw
* cell instance $12832 m0 *1 167.79,68.25
X$12832 542 50 543 644 645 cell_1rw
* cell instance $12833 m0 *1 168.495,68.25
X$12833 544 50 545 644 645 cell_1rw
* cell instance $12834 m0 *1 169.2,68.25
X$12834 546 50 547 644 645 cell_1rw
* cell instance $12835 m0 *1 169.905,68.25
X$12835 548 50 549 644 645 cell_1rw
* cell instance $12836 m0 *1 170.61,68.25
X$12836 550 50 551 644 645 cell_1rw
* cell instance $12837 m0 *1 171.315,68.25
X$12837 552 50 553 644 645 cell_1rw
* cell instance $12838 m0 *1 172.02,68.25
X$12838 554 50 555 644 645 cell_1rw
* cell instance $12839 m0 *1 172.725,68.25
X$12839 556 50 557 644 645 cell_1rw
* cell instance $12840 m0 *1 173.43,68.25
X$12840 558 50 559 644 645 cell_1rw
* cell instance $12841 m0 *1 174.135,68.25
X$12841 560 50 561 644 645 cell_1rw
* cell instance $12842 m0 *1 174.84,68.25
X$12842 562 50 563 644 645 cell_1rw
* cell instance $12843 m0 *1 175.545,68.25
X$12843 564 50 565 644 645 cell_1rw
* cell instance $12844 m0 *1 176.25,68.25
X$12844 566 50 567 644 645 cell_1rw
* cell instance $12845 m0 *1 176.955,68.25
X$12845 568 50 569 644 645 cell_1rw
* cell instance $12846 m0 *1 177.66,68.25
X$12846 570 50 571 644 645 cell_1rw
* cell instance $12847 m0 *1 178.365,68.25
X$12847 572 50 573 644 645 cell_1rw
* cell instance $12848 m0 *1 179.07,68.25
X$12848 574 50 575 644 645 cell_1rw
* cell instance $12849 m0 *1 179.775,68.25
X$12849 576 50 577 644 645 cell_1rw
* cell instance $12850 m0 *1 180.48,68.25
X$12850 578 50 579 644 645 cell_1rw
* cell instance $12851 r0 *1 0.705,68.25
X$12851 67 51 68 644 645 cell_1rw
* cell instance $12852 r0 *1 0,68.25
X$12852 65 51 66 644 645 cell_1rw
* cell instance $12853 r0 *1 1.41,68.25
X$12853 69 51 70 644 645 cell_1rw
* cell instance $12854 r0 *1 2.115,68.25
X$12854 71 51 72 644 645 cell_1rw
* cell instance $12855 r0 *1 2.82,68.25
X$12855 73 51 74 644 645 cell_1rw
* cell instance $12856 r0 *1 3.525,68.25
X$12856 75 51 76 644 645 cell_1rw
* cell instance $12857 r0 *1 4.23,68.25
X$12857 77 51 78 644 645 cell_1rw
* cell instance $12858 r0 *1 4.935,68.25
X$12858 79 51 80 644 645 cell_1rw
* cell instance $12859 r0 *1 5.64,68.25
X$12859 81 51 82 644 645 cell_1rw
* cell instance $12860 r0 *1 6.345,68.25
X$12860 83 51 84 644 645 cell_1rw
* cell instance $12861 r0 *1 7.05,68.25
X$12861 85 51 86 644 645 cell_1rw
* cell instance $12862 r0 *1 7.755,68.25
X$12862 87 51 88 644 645 cell_1rw
* cell instance $12863 r0 *1 8.46,68.25
X$12863 89 51 90 644 645 cell_1rw
* cell instance $12864 r0 *1 9.165,68.25
X$12864 91 51 92 644 645 cell_1rw
* cell instance $12865 r0 *1 9.87,68.25
X$12865 93 51 94 644 645 cell_1rw
* cell instance $12866 r0 *1 10.575,68.25
X$12866 95 51 96 644 645 cell_1rw
* cell instance $12867 r0 *1 11.28,68.25
X$12867 97 51 98 644 645 cell_1rw
* cell instance $12868 r0 *1 11.985,68.25
X$12868 99 51 100 644 645 cell_1rw
* cell instance $12869 r0 *1 12.69,68.25
X$12869 101 51 102 644 645 cell_1rw
* cell instance $12870 r0 *1 13.395,68.25
X$12870 103 51 104 644 645 cell_1rw
* cell instance $12871 r0 *1 14.1,68.25
X$12871 105 51 106 644 645 cell_1rw
* cell instance $12872 r0 *1 14.805,68.25
X$12872 107 51 108 644 645 cell_1rw
* cell instance $12873 r0 *1 15.51,68.25
X$12873 109 51 110 644 645 cell_1rw
* cell instance $12874 r0 *1 16.215,68.25
X$12874 111 51 112 644 645 cell_1rw
* cell instance $12875 r0 *1 16.92,68.25
X$12875 113 51 114 644 645 cell_1rw
* cell instance $12876 r0 *1 17.625,68.25
X$12876 115 51 116 644 645 cell_1rw
* cell instance $12877 r0 *1 18.33,68.25
X$12877 117 51 118 644 645 cell_1rw
* cell instance $12878 r0 *1 19.035,68.25
X$12878 119 51 120 644 645 cell_1rw
* cell instance $12879 r0 *1 19.74,68.25
X$12879 121 51 122 644 645 cell_1rw
* cell instance $12880 r0 *1 20.445,68.25
X$12880 123 51 124 644 645 cell_1rw
* cell instance $12881 r0 *1 21.15,68.25
X$12881 125 51 126 644 645 cell_1rw
* cell instance $12882 r0 *1 21.855,68.25
X$12882 127 51 128 644 645 cell_1rw
* cell instance $12883 r0 *1 22.56,68.25
X$12883 129 51 130 644 645 cell_1rw
* cell instance $12884 r0 *1 23.265,68.25
X$12884 131 51 132 644 645 cell_1rw
* cell instance $12885 r0 *1 23.97,68.25
X$12885 133 51 134 644 645 cell_1rw
* cell instance $12886 r0 *1 24.675,68.25
X$12886 135 51 136 644 645 cell_1rw
* cell instance $12887 r0 *1 25.38,68.25
X$12887 137 51 138 644 645 cell_1rw
* cell instance $12888 r0 *1 26.085,68.25
X$12888 139 51 140 644 645 cell_1rw
* cell instance $12889 r0 *1 26.79,68.25
X$12889 141 51 142 644 645 cell_1rw
* cell instance $12890 r0 *1 27.495,68.25
X$12890 143 51 144 644 645 cell_1rw
* cell instance $12891 r0 *1 28.2,68.25
X$12891 145 51 146 644 645 cell_1rw
* cell instance $12892 r0 *1 28.905,68.25
X$12892 147 51 148 644 645 cell_1rw
* cell instance $12893 r0 *1 29.61,68.25
X$12893 149 51 150 644 645 cell_1rw
* cell instance $12894 r0 *1 30.315,68.25
X$12894 151 51 152 644 645 cell_1rw
* cell instance $12895 r0 *1 31.02,68.25
X$12895 153 51 154 644 645 cell_1rw
* cell instance $12896 r0 *1 31.725,68.25
X$12896 155 51 156 644 645 cell_1rw
* cell instance $12897 r0 *1 32.43,68.25
X$12897 157 51 158 644 645 cell_1rw
* cell instance $12898 r0 *1 33.135,68.25
X$12898 159 51 160 644 645 cell_1rw
* cell instance $12899 r0 *1 33.84,68.25
X$12899 161 51 162 644 645 cell_1rw
* cell instance $12900 r0 *1 34.545,68.25
X$12900 163 51 164 644 645 cell_1rw
* cell instance $12901 r0 *1 35.25,68.25
X$12901 165 51 166 644 645 cell_1rw
* cell instance $12902 r0 *1 35.955,68.25
X$12902 167 51 168 644 645 cell_1rw
* cell instance $12903 r0 *1 36.66,68.25
X$12903 169 51 170 644 645 cell_1rw
* cell instance $12904 r0 *1 37.365,68.25
X$12904 171 51 172 644 645 cell_1rw
* cell instance $12905 r0 *1 38.07,68.25
X$12905 173 51 174 644 645 cell_1rw
* cell instance $12906 r0 *1 38.775,68.25
X$12906 175 51 176 644 645 cell_1rw
* cell instance $12907 r0 *1 39.48,68.25
X$12907 177 51 178 644 645 cell_1rw
* cell instance $12908 r0 *1 40.185,68.25
X$12908 179 51 180 644 645 cell_1rw
* cell instance $12909 r0 *1 40.89,68.25
X$12909 181 51 182 644 645 cell_1rw
* cell instance $12910 r0 *1 41.595,68.25
X$12910 183 51 184 644 645 cell_1rw
* cell instance $12911 r0 *1 42.3,68.25
X$12911 185 51 186 644 645 cell_1rw
* cell instance $12912 r0 *1 43.005,68.25
X$12912 187 51 188 644 645 cell_1rw
* cell instance $12913 r0 *1 43.71,68.25
X$12913 189 51 190 644 645 cell_1rw
* cell instance $12914 r0 *1 44.415,68.25
X$12914 191 51 192 644 645 cell_1rw
* cell instance $12915 r0 *1 45.12,68.25
X$12915 193 51 194 644 645 cell_1rw
* cell instance $12916 r0 *1 45.825,68.25
X$12916 195 51 196 644 645 cell_1rw
* cell instance $12917 r0 *1 46.53,68.25
X$12917 197 51 198 644 645 cell_1rw
* cell instance $12918 r0 *1 47.235,68.25
X$12918 199 51 200 644 645 cell_1rw
* cell instance $12919 r0 *1 47.94,68.25
X$12919 201 51 202 644 645 cell_1rw
* cell instance $12920 r0 *1 48.645,68.25
X$12920 203 51 204 644 645 cell_1rw
* cell instance $12921 r0 *1 49.35,68.25
X$12921 205 51 206 644 645 cell_1rw
* cell instance $12922 r0 *1 50.055,68.25
X$12922 207 51 208 644 645 cell_1rw
* cell instance $12923 r0 *1 50.76,68.25
X$12923 209 51 210 644 645 cell_1rw
* cell instance $12924 r0 *1 51.465,68.25
X$12924 211 51 212 644 645 cell_1rw
* cell instance $12925 r0 *1 52.17,68.25
X$12925 213 51 214 644 645 cell_1rw
* cell instance $12926 r0 *1 52.875,68.25
X$12926 215 51 216 644 645 cell_1rw
* cell instance $12927 r0 *1 53.58,68.25
X$12927 217 51 218 644 645 cell_1rw
* cell instance $12928 r0 *1 54.285,68.25
X$12928 219 51 220 644 645 cell_1rw
* cell instance $12929 r0 *1 54.99,68.25
X$12929 221 51 222 644 645 cell_1rw
* cell instance $12930 r0 *1 55.695,68.25
X$12930 223 51 224 644 645 cell_1rw
* cell instance $12931 r0 *1 56.4,68.25
X$12931 225 51 226 644 645 cell_1rw
* cell instance $12932 r0 *1 57.105,68.25
X$12932 227 51 228 644 645 cell_1rw
* cell instance $12933 r0 *1 57.81,68.25
X$12933 229 51 230 644 645 cell_1rw
* cell instance $12934 r0 *1 58.515,68.25
X$12934 231 51 232 644 645 cell_1rw
* cell instance $12935 r0 *1 59.22,68.25
X$12935 233 51 234 644 645 cell_1rw
* cell instance $12936 r0 *1 59.925,68.25
X$12936 235 51 236 644 645 cell_1rw
* cell instance $12937 r0 *1 60.63,68.25
X$12937 237 51 238 644 645 cell_1rw
* cell instance $12938 r0 *1 61.335,68.25
X$12938 239 51 240 644 645 cell_1rw
* cell instance $12939 r0 *1 62.04,68.25
X$12939 241 51 242 644 645 cell_1rw
* cell instance $12940 r0 *1 62.745,68.25
X$12940 243 51 244 644 645 cell_1rw
* cell instance $12941 r0 *1 63.45,68.25
X$12941 245 51 246 644 645 cell_1rw
* cell instance $12942 r0 *1 64.155,68.25
X$12942 247 51 248 644 645 cell_1rw
* cell instance $12943 r0 *1 64.86,68.25
X$12943 249 51 250 644 645 cell_1rw
* cell instance $12944 r0 *1 65.565,68.25
X$12944 251 51 252 644 645 cell_1rw
* cell instance $12945 r0 *1 66.27,68.25
X$12945 253 51 254 644 645 cell_1rw
* cell instance $12946 r0 *1 66.975,68.25
X$12946 255 51 256 644 645 cell_1rw
* cell instance $12947 r0 *1 67.68,68.25
X$12947 257 51 258 644 645 cell_1rw
* cell instance $12948 r0 *1 68.385,68.25
X$12948 259 51 260 644 645 cell_1rw
* cell instance $12949 r0 *1 69.09,68.25
X$12949 261 51 262 644 645 cell_1rw
* cell instance $12950 r0 *1 69.795,68.25
X$12950 263 51 264 644 645 cell_1rw
* cell instance $12951 r0 *1 70.5,68.25
X$12951 265 51 266 644 645 cell_1rw
* cell instance $12952 r0 *1 71.205,68.25
X$12952 267 51 268 644 645 cell_1rw
* cell instance $12953 r0 *1 71.91,68.25
X$12953 269 51 270 644 645 cell_1rw
* cell instance $12954 r0 *1 72.615,68.25
X$12954 271 51 272 644 645 cell_1rw
* cell instance $12955 r0 *1 73.32,68.25
X$12955 273 51 274 644 645 cell_1rw
* cell instance $12956 r0 *1 74.025,68.25
X$12956 275 51 276 644 645 cell_1rw
* cell instance $12957 r0 *1 74.73,68.25
X$12957 277 51 278 644 645 cell_1rw
* cell instance $12958 r0 *1 75.435,68.25
X$12958 279 51 280 644 645 cell_1rw
* cell instance $12959 r0 *1 76.14,68.25
X$12959 281 51 282 644 645 cell_1rw
* cell instance $12960 r0 *1 76.845,68.25
X$12960 283 51 284 644 645 cell_1rw
* cell instance $12961 r0 *1 77.55,68.25
X$12961 285 51 286 644 645 cell_1rw
* cell instance $12962 r0 *1 78.255,68.25
X$12962 287 51 288 644 645 cell_1rw
* cell instance $12963 r0 *1 78.96,68.25
X$12963 289 51 290 644 645 cell_1rw
* cell instance $12964 r0 *1 79.665,68.25
X$12964 291 51 292 644 645 cell_1rw
* cell instance $12965 r0 *1 80.37,68.25
X$12965 293 51 294 644 645 cell_1rw
* cell instance $12966 r0 *1 81.075,68.25
X$12966 295 51 296 644 645 cell_1rw
* cell instance $12967 r0 *1 81.78,68.25
X$12967 297 51 298 644 645 cell_1rw
* cell instance $12968 r0 *1 82.485,68.25
X$12968 299 51 300 644 645 cell_1rw
* cell instance $12969 r0 *1 83.19,68.25
X$12969 301 51 302 644 645 cell_1rw
* cell instance $12970 r0 *1 83.895,68.25
X$12970 303 51 304 644 645 cell_1rw
* cell instance $12971 r0 *1 84.6,68.25
X$12971 305 51 306 644 645 cell_1rw
* cell instance $12972 r0 *1 85.305,68.25
X$12972 307 51 308 644 645 cell_1rw
* cell instance $12973 r0 *1 86.01,68.25
X$12973 309 51 310 644 645 cell_1rw
* cell instance $12974 r0 *1 86.715,68.25
X$12974 311 51 312 644 645 cell_1rw
* cell instance $12975 r0 *1 87.42,68.25
X$12975 313 51 314 644 645 cell_1rw
* cell instance $12976 r0 *1 88.125,68.25
X$12976 315 51 316 644 645 cell_1rw
* cell instance $12977 r0 *1 88.83,68.25
X$12977 317 51 318 644 645 cell_1rw
* cell instance $12978 r0 *1 89.535,68.25
X$12978 319 51 320 644 645 cell_1rw
* cell instance $12979 r0 *1 90.24,68.25
X$12979 321 51 323 644 645 cell_1rw
* cell instance $12980 r0 *1 90.945,68.25
X$12980 324 51 325 644 645 cell_1rw
* cell instance $12981 r0 *1 91.65,68.25
X$12981 326 51 327 644 645 cell_1rw
* cell instance $12982 r0 *1 92.355,68.25
X$12982 328 51 329 644 645 cell_1rw
* cell instance $12983 r0 *1 93.06,68.25
X$12983 330 51 331 644 645 cell_1rw
* cell instance $12984 r0 *1 93.765,68.25
X$12984 332 51 333 644 645 cell_1rw
* cell instance $12985 r0 *1 94.47,68.25
X$12985 334 51 335 644 645 cell_1rw
* cell instance $12986 r0 *1 95.175,68.25
X$12986 336 51 337 644 645 cell_1rw
* cell instance $12987 r0 *1 95.88,68.25
X$12987 338 51 339 644 645 cell_1rw
* cell instance $12988 r0 *1 96.585,68.25
X$12988 340 51 341 644 645 cell_1rw
* cell instance $12989 r0 *1 97.29,68.25
X$12989 342 51 343 644 645 cell_1rw
* cell instance $12990 r0 *1 97.995,68.25
X$12990 344 51 345 644 645 cell_1rw
* cell instance $12991 r0 *1 98.7,68.25
X$12991 346 51 347 644 645 cell_1rw
* cell instance $12992 r0 *1 99.405,68.25
X$12992 348 51 349 644 645 cell_1rw
* cell instance $12993 r0 *1 100.11,68.25
X$12993 350 51 351 644 645 cell_1rw
* cell instance $12994 r0 *1 100.815,68.25
X$12994 352 51 353 644 645 cell_1rw
* cell instance $12995 r0 *1 101.52,68.25
X$12995 354 51 355 644 645 cell_1rw
* cell instance $12996 r0 *1 102.225,68.25
X$12996 356 51 357 644 645 cell_1rw
* cell instance $12997 r0 *1 102.93,68.25
X$12997 358 51 359 644 645 cell_1rw
* cell instance $12998 r0 *1 103.635,68.25
X$12998 360 51 361 644 645 cell_1rw
* cell instance $12999 r0 *1 104.34,68.25
X$12999 362 51 363 644 645 cell_1rw
* cell instance $13000 r0 *1 105.045,68.25
X$13000 364 51 365 644 645 cell_1rw
* cell instance $13001 r0 *1 105.75,68.25
X$13001 366 51 367 644 645 cell_1rw
* cell instance $13002 r0 *1 106.455,68.25
X$13002 368 51 369 644 645 cell_1rw
* cell instance $13003 r0 *1 107.16,68.25
X$13003 370 51 371 644 645 cell_1rw
* cell instance $13004 r0 *1 107.865,68.25
X$13004 372 51 373 644 645 cell_1rw
* cell instance $13005 r0 *1 108.57,68.25
X$13005 374 51 375 644 645 cell_1rw
* cell instance $13006 r0 *1 109.275,68.25
X$13006 376 51 377 644 645 cell_1rw
* cell instance $13007 r0 *1 109.98,68.25
X$13007 378 51 379 644 645 cell_1rw
* cell instance $13008 r0 *1 110.685,68.25
X$13008 380 51 381 644 645 cell_1rw
* cell instance $13009 r0 *1 111.39,68.25
X$13009 382 51 383 644 645 cell_1rw
* cell instance $13010 r0 *1 112.095,68.25
X$13010 384 51 385 644 645 cell_1rw
* cell instance $13011 r0 *1 112.8,68.25
X$13011 386 51 387 644 645 cell_1rw
* cell instance $13012 r0 *1 113.505,68.25
X$13012 388 51 389 644 645 cell_1rw
* cell instance $13013 r0 *1 114.21,68.25
X$13013 390 51 391 644 645 cell_1rw
* cell instance $13014 r0 *1 114.915,68.25
X$13014 392 51 393 644 645 cell_1rw
* cell instance $13015 r0 *1 115.62,68.25
X$13015 394 51 395 644 645 cell_1rw
* cell instance $13016 r0 *1 116.325,68.25
X$13016 396 51 397 644 645 cell_1rw
* cell instance $13017 r0 *1 117.03,68.25
X$13017 398 51 399 644 645 cell_1rw
* cell instance $13018 r0 *1 117.735,68.25
X$13018 400 51 401 644 645 cell_1rw
* cell instance $13019 r0 *1 118.44,68.25
X$13019 402 51 403 644 645 cell_1rw
* cell instance $13020 r0 *1 119.145,68.25
X$13020 404 51 405 644 645 cell_1rw
* cell instance $13021 r0 *1 119.85,68.25
X$13021 406 51 407 644 645 cell_1rw
* cell instance $13022 r0 *1 120.555,68.25
X$13022 408 51 409 644 645 cell_1rw
* cell instance $13023 r0 *1 121.26,68.25
X$13023 410 51 411 644 645 cell_1rw
* cell instance $13024 r0 *1 121.965,68.25
X$13024 412 51 413 644 645 cell_1rw
* cell instance $13025 r0 *1 122.67,68.25
X$13025 414 51 415 644 645 cell_1rw
* cell instance $13026 r0 *1 123.375,68.25
X$13026 416 51 417 644 645 cell_1rw
* cell instance $13027 r0 *1 124.08,68.25
X$13027 418 51 419 644 645 cell_1rw
* cell instance $13028 r0 *1 124.785,68.25
X$13028 420 51 421 644 645 cell_1rw
* cell instance $13029 r0 *1 125.49,68.25
X$13029 422 51 423 644 645 cell_1rw
* cell instance $13030 r0 *1 126.195,68.25
X$13030 424 51 425 644 645 cell_1rw
* cell instance $13031 r0 *1 126.9,68.25
X$13031 426 51 427 644 645 cell_1rw
* cell instance $13032 r0 *1 127.605,68.25
X$13032 428 51 429 644 645 cell_1rw
* cell instance $13033 r0 *1 128.31,68.25
X$13033 430 51 431 644 645 cell_1rw
* cell instance $13034 r0 *1 129.015,68.25
X$13034 432 51 433 644 645 cell_1rw
* cell instance $13035 r0 *1 129.72,68.25
X$13035 434 51 435 644 645 cell_1rw
* cell instance $13036 r0 *1 130.425,68.25
X$13036 436 51 437 644 645 cell_1rw
* cell instance $13037 r0 *1 131.13,68.25
X$13037 438 51 439 644 645 cell_1rw
* cell instance $13038 r0 *1 131.835,68.25
X$13038 440 51 441 644 645 cell_1rw
* cell instance $13039 r0 *1 132.54,68.25
X$13039 442 51 443 644 645 cell_1rw
* cell instance $13040 r0 *1 133.245,68.25
X$13040 444 51 445 644 645 cell_1rw
* cell instance $13041 r0 *1 133.95,68.25
X$13041 446 51 447 644 645 cell_1rw
* cell instance $13042 r0 *1 134.655,68.25
X$13042 448 51 449 644 645 cell_1rw
* cell instance $13043 r0 *1 135.36,68.25
X$13043 450 51 451 644 645 cell_1rw
* cell instance $13044 r0 *1 136.065,68.25
X$13044 452 51 453 644 645 cell_1rw
* cell instance $13045 r0 *1 136.77,68.25
X$13045 454 51 455 644 645 cell_1rw
* cell instance $13046 r0 *1 137.475,68.25
X$13046 456 51 457 644 645 cell_1rw
* cell instance $13047 r0 *1 138.18,68.25
X$13047 458 51 459 644 645 cell_1rw
* cell instance $13048 r0 *1 138.885,68.25
X$13048 460 51 461 644 645 cell_1rw
* cell instance $13049 r0 *1 139.59,68.25
X$13049 462 51 463 644 645 cell_1rw
* cell instance $13050 r0 *1 140.295,68.25
X$13050 464 51 465 644 645 cell_1rw
* cell instance $13051 r0 *1 141,68.25
X$13051 466 51 467 644 645 cell_1rw
* cell instance $13052 r0 *1 141.705,68.25
X$13052 468 51 469 644 645 cell_1rw
* cell instance $13053 r0 *1 142.41,68.25
X$13053 470 51 471 644 645 cell_1rw
* cell instance $13054 r0 *1 143.115,68.25
X$13054 472 51 473 644 645 cell_1rw
* cell instance $13055 r0 *1 143.82,68.25
X$13055 474 51 475 644 645 cell_1rw
* cell instance $13056 r0 *1 144.525,68.25
X$13056 476 51 477 644 645 cell_1rw
* cell instance $13057 r0 *1 145.23,68.25
X$13057 478 51 479 644 645 cell_1rw
* cell instance $13058 r0 *1 145.935,68.25
X$13058 480 51 481 644 645 cell_1rw
* cell instance $13059 r0 *1 146.64,68.25
X$13059 482 51 483 644 645 cell_1rw
* cell instance $13060 r0 *1 147.345,68.25
X$13060 484 51 485 644 645 cell_1rw
* cell instance $13061 r0 *1 148.05,68.25
X$13061 486 51 487 644 645 cell_1rw
* cell instance $13062 r0 *1 148.755,68.25
X$13062 488 51 489 644 645 cell_1rw
* cell instance $13063 r0 *1 149.46,68.25
X$13063 490 51 491 644 645 cell_1rw
* cell instance $13064 r0 *1 150.165,68.25
X$13064 492 51 493 644 645 cell_1rw
* cell instance $13065 r0 *1 150.87,68.25
X$13065 494 51 495 644 645 cell_1rw
* cell instance $13066 r0 *1 151.575,68.25
X$13066 496 51 497 644 645 cell_1rw
* cell instance $13067 r0 *1 152.28,68.25
X$13067 498 51 499 644 645 cell_1rw
* cell instance $13068 r0 *1 152.985,68.25
X$13068 500 51 501 644 645 cell_1rw
* cell instance $13069 r0 *1 153.69,68.25
X$13069 502 51 503 644 645 cell_1rw
* cell instance $13070 r0 *1 154.395,68.25
X$13070 504 51 505 644 645 cell_1rw
* cell instance $13071 r0 *1 155.1,68.25
X$13071 506 51 507 644 645 cell_1rw
* cell instance $13072 r0 *1 155.805,68.25
X$13072 508 51 509 644 645 cell_1rw
* cell instance $13073 r0 *1 156.51,68.25
X$13073 510 51 511 644 645 cell_1rw
* cell instance $13074 r0 *1 157.215,68.25
X$13074 512 51 513 644 645 cell_1rw
* cell instance $13075 r0 *1 157.92,68.25
X$13075 514 51 515 644 645 cell_1rw
* cell instance $13076 r0 *1 158.625,68.25
X$13076 516 51 517 644 645 cell_1rw
* cell instance $13077 r0 *1 159.33,68.25
X$13077 518 51 519 644 645 cell_1rw
* cell instance $13078 r0 *1 160.035,68.25
X$13078 520 51 521 644 645 cell_1rw
* cell instance $13079 r0 *1 160.74,68.25
X$13079 522 51 523 644 645 cell_1rw
* cell instance $13080 r0 *1 161.445,68.25
X$13080 524 51 525 644 645 cell_1rw
* cell instance $13081 r0 *1 162.15,68.25
X$13081 526 51 527 644 645 cell_1rw
* cell instance $13082 r0 *1 162.855,68.25
X$13082 528 51 529 644 645 cell_1rw
* cell instance $13083 r0 *1 163.56,68.25
X$13083 530 51 531 644 645 cell_1rw
* cell instance $13084 r0 *1 164.265,68.25
X$13084 532 51 533 644 645 cell_1rw
* cell instance $13085 r0 *1 164.97,68.25
X$13085 534 51 535 644 645 cell_1rw
* cell instance $13086 r0 *1 165.675,68.25
X$13086 536 51 537 644 645 cell_1rw
* cell instance $13087 r0 *1 166.38,68.25
X$13087 538 51 539 644 645 cell_1rw
* cell instance $13088 r0 *1 167.085,68.25
X$13088 540 51 541 644 645 cell_1rw
* cell instance $13089 r0 *1 167.79,68.25
X$13089 542 51 543 644 645 cell_1rw
* cell instance $13090 r0 *1 168.495,68.25
X$13090 544 51 545 644 645 cell_1rw
* cell instance $13091 r0 *1 169.2,68.25
X$13091 546 51 547 644 645 cell_1rw
* cell instance $13092 r0 *1 169.905,68.25
X$13092 548 51 549 644 645 cell_1rw
* cell instance $13093 r0 *1 170.61,68.25
X$13093 550 51 551 644 645 cell_1rw
* cell instance $13094 r0 *1 171.315,68.25
X$13094 552 51 553 644 645 cell_1rw
* cell instance $13095 r0 *1 172.02,68.25
X$13095 554 51 555 644 645 cell_1rw
* cell instance $13096 r0 *1 172.725,68.25
X$13096 556 51 557 644 645 cell_1rw
* cell instance $13097 r0 *1 173.43,68.25
X$13097 558 51 559 644 645 cell_1rw
* cell instance $13098 r0 *1 174.135,68.25
X$13098 560 51 561 644 645 cell_1rw
* cell instance $13099 r0 *1 174.84,68.25
X$13099 562 51 563 644 645 cell_1rw
* cell instance $13100 r0 *1 175.545,68.25
X$13100 564 51 565 644 645 cell_1rw
* cell instance $13101 r0 *1 176.25,68.25
X$13101 566 51 567 644 645 cell_1rw
* cell instance $13102 r0 *1 176.955,68.25
X$13102 568 51 569 644 645 cell_1rw
* cell instance $13103 r0 *1 177.66,68.25
X$13103 570 51 571 644 645 cell_1rw
* cell instance $13104 r0 *1 178.365,68.25
X$13104 572 51 573 644 645 cell_1rw
* cell instance $13105 r0 *1 179.07,68.25
X$13105 574 51 575 644 645 cell_1rw
* cell instance $13106 r0 *1 179.775,68.25
X$13106 576 51 577 644 645 cell_1rw
* cell instance $13107 r0 *1 180.48,68.25
X$13107 578 51 579 644 645 cell_1rw
* cell instance $13108 m0 *1 0.705,70.98
X$13108 67 52 68 644 645 cell_1rw
* cell instance $13109 m0 *1 0,70.98
X$13109 65 52 66 644 645 cell_1rw
* cell instance $13110 m0 *1 1.41,70.98
X$13110 69 52 70 644 645 cell_1rw
* cell instance $13111 m0 *1 2.115,70.98
X$13111 71 52 72 644 645 cell_1rw
* cell instance $13112 m0 *1 2.82,70.98
X$13112 73 52 74 644 645 cell_1rw
* cell instance $13113 m0 *1 3.525,70.98
X$13113 75 52 76 644 645 cell_1rw
* cell instance $13114 m0 *1 4.23,70.98
X$13114 77 52 78 644 645 cell_1rw
* cell instance $13115 m0 *1 4.935,70.98
X$13115 79 52 80 644 645 cell_1rw
* cell instance $13116 m0 *1 5.64,70.98
X$13116 81 52 82 644 645 cell_1rw
* cell instance $13117 m0 *1 6.345,70.98
X$13117 83 52 84 644 645 cell_1rw
* cell instance $13118 m0 *1 7.05,70.98
X$13118 85 52 86 644 645 cell_1rw
* cell instance $13119 m0 *1 7.755,70.98
X$13119 87 52 88 644 645 cell_1rw
* cell instance $13120 m0 *1 8.46,70.98
X$13120 89 52 90 644 645 cell_1rw
* cell instance $13121 m0 *1 9.165,70.98
X$13121 91 52 92 644 645 cell_1rw
* cell instance $13122 m0 *1 9.87,70.98
X$13122 93 52 94 644 645 cell_1rw
* cell instance $13123 m0 *1 10.575,70.98
X$13123 95 52 96 644 645 cell_1rw
* cell instance $13124 m0 *1 11.28,70.98
X$13124 97 52 98 644 645 cell_1rw
* cell instance $13125 m0 *1 11.985,70.98
X$13125 99 52 100 644 645 cell_1rw
* cell instance $13126 m0 *1 12.69,70.98
X$13126 101 52 102 644 645 cell_1rw
* cell instance $13127 m0 *1 13.395,70.98
X$13127 103 52 104 644 645 cell_1rw
* cell instance $13128 m0 *1 14.1,70.98
X$13128 105 52 106 644 645 cell_1rw
* cell instance $13129 m0 *1 14.805,70.98
X$13129 107 52 108 644 645 cell_1rw
* cell instance $13130 m0 *1 15.51,70.98
X$13130 109 52 110 644 645 cell_1rw
* cell instance $13131 m0 *1 16.215,70.98
X$13131 111 52 112 644 645 cell_1rw
* cell instance $13132 m0 *1 16.92,70.98
X$13132 113 52 114 644 645 cell_1rw
* cell instance $13133 m0 *1 17.625,70.98
X$13133 115 52 116 644 645 cell_1rw
* cell instance $13134 m0 *1 18.33,70.98
X$13134 117 52 118 644 645 cell_1rw
* cell instance $13135 m0 *1 19.035,70.98
X$13135 119 52 120 644 645 cell_1rw
* cell instance $13136 m0 *1 19.74,70.98
X$13136 121 52 122 644 645 cell_1rw
* cell instance $13137 m0 *1 20.445,70.98
X$13137 123 52 124 644 645 cell_1rw
* cell instance $13138 m0 *1 21.15,70.98
X$13138 125 52 126 644 645 cell_1rw
* cell instance $13139 m0 *1 21.855,70.98
X$13139 127 52 128 644 645 cell_1rw
* cell instance $13140 m0 *1 22.56,70.98
X$13140 129 52 130 644 645 cell_1rw
* cell instance $13141 m0 *1 23.265,70.98
X$13141 131 52 132 644 645 cell_1rw
* cell instance $13142 m0 *1 23.97,70.98
X$13142 133 52 134 644 645 cell_1rw
* cell instance $13143 m0 *1 24.675,70.98
X$13143 135 52 136 644 645 cell_1rw
* cell instance $13144 m0 *1 25.38,70.98
X$13144 137 52 138 644 645 cell_1rw
* cell instance $13145 m0 *1 26.085,70.98
X$13145 139 52 140 644 645 cell_1rw
* cell instance $13146 m0 *1 26.79,70.98
X$13146 141 52 142 644 645 cell_1rw
* cell instance $13147 m0 *1 27.495,70.98
X$13147 143 52 144 644 645 cell_1rw
* cell instance $13148 m0 *1 28.2,70.98
X$13148 145 52 146 644 645 cell_1rw
* cell instance $13149 m0 *1 28.905,70.98
X$13149 147 52 148 644 645 cell_1rw
* cell instance $13150 m0 *1 29.61,70.98
X$13150 149 52 150 644 645 cell_1rw
* cell instance $13151 m0 *1 30.315,70.98
X$13151 151 52 152 644 645 cell_1rw
* cell instance $13152 m0 *1 31.02,70.98
X$13152 153 52 154 644 645 cell_1rw
* cell instance $13153 m0 *1 31.725,70.98
X$13153 155 52 156 644 645 cell_1rw
* cell instance $13154 m0 *1 32.43,70.98
X$13154 157 52 158 644 645 cell_1rw
* cell instance $13155 m0 *1 33.135,70.98
X$13155 159 52 160 644 645 cell_1rw
* cell instance $13156 m0 *1 33.84,70.98
X$13156 161 52 162 644 645 cell_1rw
* cell instance $13157 m0 *1 34.545,70.98
X$13157 163 52 164 644 645 cell_1rw
* cell instance $13158 m0 *1 35.25,70.98
X$13158 165 52 166 644 645 cell_1rw
* cell instance $13159 m0 *1 35.955,70.98
X$13159 167 52 168 644 645 cell_1rw
* cell instance $13160 m0 *1 36.66,70.98
X$13160 169 52 170 644 645 cell_1rw
* cell instance $13161 m0 *1 37.365,70.98
X$13161 171 52 172 644 645 cell_1rw
* cell instance $13162 m0 *1 38.07,70.98
X$13162 173 52 174 644 645 cell_1rw
* cell instance $13163 m0 *1 38.775,70.98
X$13163 175 52 176 644 645 cell_1rw
* cell instance $13164 m0 *1 39.48,70.98
X$13164 177 52 178 644 645 cell_1rw
* cell instance $13165 m0 *1 40.185,70.98
X$13165 179 52 180 644 645 cell_1rw
* cell instance $13166 m0 *1 40.89,70.98
X$13166 181 52 182 644 645 cell_1rw
* cell instance $13167 m0 *1 41.595,70.98
X$13167 183 52 184 644 645 cell_1rw
* cell instance $13168 m0 *1 42.3,70.98
X$13168 185 52 186 644 645 cell_1rw
* cell instance $13169 m0 *1 43.005,70.98
X$13169 187 52 188 644 645 cell_1rw
* cell instance $13170 m0 *1 43.71,70.98
X$13170 189 52 190 644 645 cell_1rw
* cell instance $13171 m0 *1 44.415,70.98
X$13171 191 52 192 644 645 cell_1rw
* cell instance $13172 m0 *1 45.12,70.98
X$13172 193 52 194 644 645 cell_1rw
* cell instance $13173 m0 *1 45.825,70.98
X$13173 195 52 196 644 645 cell_1rw
* cell instance $13174 m0 *1 46.53,70.98
X$13174 197 52 198 644 645 cell_1rw
* cell instance $13175 m0 *1 47.235,70.98
X$13175 199 52 200 644 645 cell_1rw
* cell instance $13176 m0 *1 47.94,70.98
X$13176 201 52 202 644 645 cell_1rw
* cell instance $13177 m0 *1 48.645,70.98
X$13177 203 52 204 644 645 cell_1rw
* cell instance $13178 m0 *1 49.35,70.98
X$13178 205 52 206 644 645 cell_1rw
* cell instance $13179 m0 *1 50.055,70.98
X$13179 207 52 208 644 645 cell_1rw
* cell instance $13180 m0 *1 50.76,70.98
X$13180 209 52 210 644 645 cell_1rw
* cell instance $13181 m0 *1 51.465,70.98
X$13181 211 52 212 644 645 cell_1rw
* cell instance $13182 m0 *1 52.17,70.98
X$13182 213 52 214 644 645 cell_1rw
* cell instance $13183 m0 *1 52.875,70.98
X$13183 215 52 216 644 645 cell_1rw
* cell instance $13184 m0 *1 53.58,70.98
X$13184 217 52 218 644 645 cell_1rw
* cell instance $13185 m0 *1 54.285,70.98
X$13185 219 52 220 644 645 cell_1rw
* cell instance $13186 m0 *1 54.99,70.98
X$13186 221 52 222 644 645 cell_1rw
* cell instance $13187 m0 *1 55.695,70.98
X$13187 223 52 224 644 645 cell_1rw
* cell instance $13188 m0 *1 56.4,70.98
X$13188 225 52 226 644 645 cell_1rw
* cell instance $13189 m0 *1 57.105,70.98
X$13189 227 52 228 644 645 cell_1rw
* cell instance $13190 m0 *1 57.81,70.98
X$13190 229 52 230 644 645 cell_1rw
* cell instance $13191 m0 *1 58.515,70.98
X$13191 231 52 232 644 645 cell_1rw
* cell instance $13192 m0 *1 59.22,70.98
X$13192 233 52 234 644 645 cell_1rw
* cell instance $13193 m0 *1 59.925,70.98
X$13193 235 52 236 644 645 cell_1rw
* cell instance $13194 m0 *1 60.63,70.98
X$13194 237 52 238 644 645 cell_1rw
* cell instance $13195 m0 *1 61.335,70.98
X$13195 239 52 240 644 645 cell_1rw
* cell instance $13196 m0 *1 62.04,70.98
X$13196 241 52 242 644 645 cell_1rw
* cell instance $13197 m0 *1 62.745,70.98
X$13197 243 52 244 644 645 cell_1rw
* cell instance $13198 m0 *1 63.45,70.98
X$13198 245 52 246 644 645 cell_1rw
* cell instance $13199 m0 *1 64.155,70.98
X$13199 247 52 248 644 645 cell_1rw
* cell instance $13200 m0 *1 64.86,70.98
X$13200 249 52 250 644 645 cell_1rw
* cell instance $13201 m0 *1 65.565,70.98
X$13201 251 52 252 644 645 cell_1rw
* cell instance $13202 m0 *1 66.27,70.98
X$13202 253 52 254 644 645 cell_1rw
* cell instance $13203 m0 *1 66.975,70.98
X$13203 255 52 256 644 645 cell_1rw
* cell instance $13204 m0 *1 67.68,70.98
X$13204 257 52 258 644 645 cell_1rw
* cell instance $13205 m0 *1 68.385,70.98
X$13205 259 52 260 644 645 cell_1rw
* cell instance $13206 m0 *1 69.09,70.98
X$13206 261 52 262 644 645 cell_1rw
* cell instance $13207 m0 *1 69.795,70.98
X$13207 263 52 264 644 645 cell_1rw
* cell instance $13208 m0 *1 70.5,70.98
X$13208 265 52 266 644 645 cell_1rw
* cell instance $13209 m0 *1 71.205,70.98
X$13209 267 52 268 644 645 cell_1rw
* cell instance $13210 m0 *1 71.91,70.98
X$13210 269 52 270 644 645 cell_1rw
* cell instance $13211 m0 *1 72.615,70.98
X$13211 271 52 272 644 645 cell_1rw
* cell instance $13212 m0 *1 73.32,70.98
X$13212 273 52 274 644 645 cell_1rw
* cell instance $13213 m0 *1 74.025,70.98
X$13213 275 52 276 644 645 cell_1rw
* cell instance $13214 m0 *1 74.73,70.98
X$13214 277 52 278 644 645 cell_1rw
* cell instance $13215 m0 *1 75.435,70.98
X$13215 279 52 280 644 645 cell_1rw
* cell instance $13216 m0 *1 76.14,70.98
X$13216 281 52 282 644 645 cell_1rw
* cell instance $13217 m0 *1 76.845,70.98
X$13217 283 52 284 644 645 cell_1rw
* cell instance $13218 m0 *1 77.55,70.98
X$13218 285 52 286 644 645 cell_1rw
* cell instance $13219 m0 *1 78.255,70.98
X$13219 287 52 288 644 645 cell_1rw
* cell instance $13220 m0 *1 78.96,70.98
X$13220 289 52 290 644 645 cell_1rw
* cell instance $13221 m0 *1 79.665,70.98
X$13221 291 52 292 644 645 cell_1rw
* cell instance $13222 m0 *1 80.37,70.98
X$13222 293 52 294 644 645 cell_1rw
* cell instance $13223 m0 *1 81.075,70.98
X$13223 295 52 296 644 645 cell_1rw
* cell instance $13224 m0 *1 81.78,70.98
X$13224 297 52 298 644 645 cell_1rw
* cell instance $13225 m0 *1 82.485,70.98
X$13225 299 52 300 644 645 cell_1rw
* cell instance $13226 m0 *1 83.19,70.98
X$13226 301 52 302 644 645 cell_1rw
* cell instance $13227 m0 *1 83.895,70.98
X$13227 303 52 304 644 645 cell_1rw
* cell instance $13228 m0 *1 84.6,70.98
X$13228 305 52 306 644 645 cell_1rw
* cell instance $13229 m0 *1 85.305,70.98
X$13229 307 52 308 644 645 cell_1rw
* cell instance $13230 m0 *1 86.01,70.98
X$13230 309 52 310 644 645 cell_1rw
* cell instance $13231 m0 *1 86.715,70.98
X$13231 311 52 312 644 645 cell_1rw
* cell instance $13232 m0 *1 87.42,70.98
X$13232 313 52 314 644 645 cell_1rw
* cell instance $13233 m0 *1 88.125,70.98
X$13233 315 52 316 644 645 cell_1rw
* cell instance $13234 m0 *1 88.83,70.98
X$13234 317 52 318 644 645 cell_1rw
* cell instance $13235 m0 *1 89.535,70.98
X$13235 319 52 320 644 645 cell_1rw
* cell instance $13236 m0 *1 90.24,70.98
X$13236 321 52 323 644 645 cell_1rw
* cell instance $13237 m0 *1 90.945,70.98
X$13237 324 52 325 644 645 cell_1rw
* cell instance $13238 m0 *1 91.65,70.98
X$13238 326 52 327 644 645 cell_1rw
* cell instance $13239 m0 *1 92.355,70.98
X$13239 328 52 329 644 645 cell_1rw
* cell instance $13240 m0 *1 93.06,70.98
X$13240 330 52 331 644 645 cell_1rw
* cell instance $13241 m0 *1 93.765,70.98
X$13241 332 52 333 644 645 cell_1rw
* cell instance $13242 m0 *1 94.47,70.98
X$13242 334 52 335 644 645 cell_1rw
* cell instance $13243 m0 *1 95.175,70.98
X$13243 336 52 337 644 645 cell_1rw
* cell instance $13244 m0 *1 95.88,70.98
X$13244 338 52 339 644 645 cell_1rw
* cell instance $13245 m0 *1 96.585,70.98
X$13245 340 52 341 644 645 cell_1rw
* cell instance $13246 m0 *1 97.29,70.98
X$13246 342 52 343 644 645 cell_1rw
* cell instance $13247 m0 *1 97.995,70.98
X$13247 344 52 345 644 645 cell_1rw
* cell instance $13248 m0 *1 98.7,70.98
X$13248 346 52 347 644 645 cell_1rw
* cell instance $13249 m0 *1 99.405,70.98
X$13249 348 52 349 644 645 cell_1rw
* cell instance $13250 m0 *1 100.11,70.98
X$13250 350 52 351 644 645 cell_1rw
* cell instance $13251 m0 *1 100.815,70.98
X$13251 352 52 353 644 645 cell_1rw
* cell instance $13252 m0 *1 101.52,70.98
X$13252 354 52 355 644 645 cell_1rw
* cell instance $13253 m0 *1 102.225,70.98
X$13253 356 52 357 644 645 cell_1rw
* cell instance $13254 m0 *1 102.93,70.98
X$13254 358 52 359 644 645 cell_1rw
* cell instance $13255 m0 *1 103.635,70.98
X$13255 360 52 361 644 645 cell_1rw
* cell instance $13256 m0 *1 104.34,70.98
X$13256 362 52 363 644 645 cell_1rw
* cell instance $13257 m0 *1 105.045,70.98
X$13257 364 52 365 644 645 cell_1rw
* cell instance $13258 m0 *1 105.75,70.98
X$13258 366 52 367 644 645 cell_1rw
* cell instance $13259 m0 *1 106.455,70.98
X$13259 368 52 369 644 645 cell_1rw
* cell instance $13260 m0 *1 107.16,70.98
X$13260 370 52 371 644 645 cell_1rw
* cell instance $13261 m0 *1 107.865,70.98
X$13261 372 52 373 644 645 cell_1rw
* cell instance $13262 m0 *1 108.57,70.98
X$13262 374 52 375 644 645 cell_1rw
* cell instance $13263 m0 *1 109.275,70.98
X$13263 376 52 377 644 645 cell_1rw
* cell instance $13264 m0 *1 109.98,70.98
X$13264 378 52 379 644 645 cell_1rw
* cell instance $13265 m0 *1 110.685,70.98
X$13265 380 52 381 644 645 cell_1rw
* cell instance $13266 m0 *1 111.39,70.98
X$13266 382 52 383 644 645 cell_1rw
* cell instance $13267 m0 *1 112.095,70.98
X$13267 384 52 385 644 645 cell_1rw
* cell instance $13268 m0 *1 112.8,70.98
X$13268 386 52 387 644 645 cell_1rw
* cell instance $13269 m0 *1 113.505,70.98
X$13269 388 52 389 644 645 cell_1rw
* cell instance $13270 m0 *1 114.21,70.98
X$13270 390 52 391 644 645 cell_1rw
* cell instance $13271 m0 *1 114.915,70.98
X$13271 392 52 393 644 645 cell_1rw
* cell instance $13272 m0 *1 115.62,70.98
X$13272 394 52 395 644 645 cell_1rw
* cell instance $13273 m0 *1 116.325,70.98
X$13273 396 52 397 644 645 cell_1rw
* cell instance $13274 m0 *1 117.03,70.98
X$13274 398 52 399 644 645 cell_1rw
* cell instance $13275 m0 *1 117.735,70.98
X$13275 400 52 401 644 645 cell_1rw
* cell instance $13276 m0 *1 118.44,70.98
X$13276 402 52 403 644 645 cell_1rw
* cell instance $13277 m0 *1 119.145,70.98
X$13277 404 52 405 644 645 cell_1rw
* cell instance $13278 m0 *1 119.85,70.98
X$13278 406 52 407 644 645 cell_1rw
* cell instance $13279 m0 *1 120.555,70.98
X$13279 408 52 409 644 645 cell_1rw
* cell instance $13280 m0 *1 121.26,70.98
X$13280 410 52 411 644 645 cell_1rw
* cell instance $13281 m0 *1 121.965,70.98
X$13281 412 52 413 644 645 cell_1rw
* cell instance $13282 m0 *1 122.67,70.98
X$13282 414 52 415 644 645 cell_1rw
* cell instance $13283 m0 *1 123.375,70.98
X$13283 416 52 417 644 645 cell_1rw
* cell instance $13284 m0 *1 124.08,70.98
X$13284 418 52 419 644 645 cell_1rw
* cell instance $13285 m0 *1 124.785,70.98
X$13285 420 52 421 644 645 cell_1rw
* cell instance $13286 m0 *1 125.49,70.98
X$13286 422 52 423 644 645 cell_1rw
* cell instance $13287 m0 *1 126.195,70.98
X$13287 424 52 425 644 645 cell_1rw
* cell instance $13288 m0 *1 126.9,70.98
X$13288 426 52 427 644 645 cell_1rw
* cell instance $13289 m0 *1 127.605,70.98
X$13289 428 52 429 644 645 cell_1rw
* cell instance $13290 m0 *1 128.31,70.98
X$13290 430 52 431 644 645 cell_1rw
* cell instance $13291 m0 *1 129.015,70.98
X$13291 432 52 433 644 645 cell_1rw
* cell instance $13292 m0 *1 129.72,70.98
X$13292 434 52 435 644 645 cell_1rw
* cell instance $13293 m0 *1 130.425,70.98
X$13293 436 52 437 644 645 cell_1rw
* cell instance $13294 m0 *1 131.13,70.98
X$13294 438 52 439 644 645 cell_1rw
* cell instance $13295 m0 *1 131.835,70.98
X$13295 440 52 441 644 645 cell_1rw
* cell instance $13296 m0 *1 132.54,70.98
X$13296 442 52 443 644 645 cell_1rw
* cell instance $13297 m0 *1 133.245,70.98
X$13297 444 52 445 644 645 cell_1rw
* cell instance $13298 m0 *1 133.95,70.98
X$13298 446 52 447 644 645 cell_1rw
* cell instance $13299 m0 *1 134.655,70.98
X$13299 448 52 449 644 645 cell_1rw
* cell instance $13300 m0 *1 135.36,70.98
X$13300 450 52 451 644 645 cell_1rw
* cell instance $13301 m0 *1 136.065,70.98
X$13301 452 52 453 644 645 cell_1rw
* cell instance $13302 m0 *1 136.77,70.98
X$13302 454 52 455 644 645 cell_1rw
* cell instance $13303 m0 *1 137.475,70.98
X$13303 456 52 457 644 645 cell_1rw
* cell instance $13304 m0 *1 138.18,70.98
X$13304 458 52 459 644 645 cell_1rw
* cell instance $13305 m0 *1 138.885,70.98
X$13305 460 52 461 644 645 cell_1rw
* cell instance $13306 m0 *1 139.59,70.98
X$13306 462 52 463 644 645 cell_1rw
* cell instance $13307 m0 *1 140.295,70.98
X$13307 464 52 465 644 645 cell_1rw
* cell instance $13308 m0 *1 141,70.98
X$13308 466 52 467 644 645 cell_1rw
* cell instance $13309 m0 *1 141.705,70.98
X$13309 468 52 469 644 645 cell_1rw
* cell instance $13310 m0 *1 142.41,70.98
X$13310 470 52 471 644 645 cell_1rw
* cell instance $13311 m0 *1 143.115,70.98
X$13311 472 52 473 644 645 cell_1rw
* cell instance $13312 m0 *1 143.82,70.98
X$13312 474 52 475 644 645 cell_1rw
* cell instance $13313 m0 *1 144.525,70.98
X$13313 476 52 477 644 645 cell_1rw
* cell instance $13314 m0 *1 145.23,70.98
X$13314 478 52 479 644 645 cell_1rw
* cell instance $13315 m0 *1 145.935,70.98
X$13315 480 52 481 644 645 cell_1rw
* cell instance $13316 m0 *1 146.64,70.98
X$13316 482 52 483 644 645 cell_1rw
* cell instance $13317 m0 *1 147.345,70.98
X$13317 484 52 485 644 645 cell_1rw
* cell instance $13318 m0 *1 148.05,70.98
X$13318 486 52 487 644 645 cell_1rw
* cell instance $13319 m0 *1 148.755,70.98
X$13319 488 52 489 644 645 cell_1rw
* cell instance $13320 m0 *1 149.46,70.98
X$13320 490 52 491 644 645 cell_1rw
* cell instance $13321 m0 *1 150.165,70.98
X$13321 492 52 493 644 645 cell_1rw
* cell instance $13322 m0 *1 150.87,70.98
X$13322 494 52 495 644 645 cell_1rw
* cell instance $13323 m0 *1 151.575,70.98
X$13323 496 52 497 644 645 cell_1rw
* cell instance $13324 m0 *1 152.28,70.98
X$13324 498 52 499 644 645 cell_1rw
* cell instance $13325 m0 *1 152.985,70.98
X$13325 500 52 501 644 645 cell_1rw
* cell instance $13326 m0 *1 153.69,70.98
X$13326 502 52 503 644 645 cell_1rw
* cell instance $13327 m0 *1 154.395,70.98
X$13327 504 52 505 644 645 cell_1rw
* cell instance $13328 m0 *1 155.1,70.98
X$13328 506 52 507 644 645 cell_1rw
* cell instance $13329 m0 *1 155.805,70.98
X$13329 508 52 509 644 645 cell_1rw
* cell instance $13330 m0 *1 156.51,70.98
X$13330 510 52 511 644 645 cell_1rw
* cell instance $13331 m0 *1 157.215,70.98
X$13331 512 52 513 644 645 cell_1rw
* cell instance $13332 m0 *1 157.92,70.98
X$13332 514 52 515 644 645 cell_1rw
* cell instance $13333 m0 *1 158.625,70.98
X$13333 516 52 517 644 645 cell_1rw
* cell instance $13334 m0 *1 159.33,70.98
X$13334 518 52 519 644 645 cell_1rw
* cell instance $13335 m0 *1 160.035,70.98
X$13335 520 52 521 644 645 cell_1rw
* cell instance $13336 m0 *1 160.74,70.98
X$13336 522 52 523 644 645 cell_1rw
* cell instance $13337 m0 *1 161.445,70.98
X$13337 524 52 525 644 645 cell_1rw
* cell instance $13338 m0 *1 162.15,70.98
X$13338 526 52 527 644 645 cell_1rw
* cell instance $13339 m0 *1 162.855,70.98
X$13339 528 52 529 644 645 cell_1rw
* cell instance $13340 m0 *1 163.56,70.98
X$13340 530 52 531 644 645 cell_1rw
* cell instance $13341 m0 *1 164.265,70.98
X$13341 532 52 533 644 645 cell_1rw
* cell instance $13342 m0 *1 164.97,70.98
X$13342 534 52 535 644 645 cell_1rw
* cell instance $13343 m0 *1 165.675,70.98
X$13343 536 52 537 644 645 cell_1rw
* cell instance $13344 m0 *1 166.38,70.98
X$13344 538 52 539 644 645 cell_1rw
* cell instance $13345 m0 *1 167.085,70.98
X$13345 540 52 541 644 645 cell_1rw
* cell instance $13346 m0 *1 167.79,70.98
X$13346 542 52 543 644 645 cell_1rw
* cell instance $13347 m0 *1 168.495,70.98
X$13347 544 52 545 644 645 cell_1rw
* cell instance $13348 m0 *1 169.2,70.98
X$13348 546 52 547 644 645 cell_1rw
* cell instance $13349 m0 *1 169.905,70.98
X$13349 548 52 549 644 645 cell_1rw
* cell instance $13350 m0 *1 170.61,70.98
X$13350 550 52 551 644 645 cell_1rw
* cell instance $13351 m0 *1 171.315,70.98
X$13351 552 52 553 644 645 cell_1rw
* cell instance $13352 m0 *1 172.02,70.98
X$13352 554 52 555 644 645 cell_1rw
* cell instance $13353 m0 *1 172.725,70.98
X$13353 556 52 557 644 645 cell_1rw
* cell instance $13354 m0 *1 173.43,70.98
X$13354 558 52 559 644 645 cell_1rw
* cell instance $13355 m0 *1 174.135,70.98
X$13355 560 52 561 644 645 cell_1rw
* cell instance $13356 m0 *1 174.84,70.98
X$13356 562 52 563 644 645 cell_1rw
* cell instance $13357 m0 *1 175.545,70.98
X$13357 564 52 565 644 645 cell_1rw
* cell instance $13358 m0 *1 176.25,70.98
X$13358 566 52 567 644 645 cell_1rw
* cell instance $13359 m0 *1 176.955,70.98
X$13359 568 52 569 644 645 cell_1rw
* cell instance $13360 m0 *1 177.66,70.98
X$13360 570 52 571 644 645 cell_1rw
* cell instance $13361 m0 *1 178.365,70.98
X$13361 572 52 573 644 645 cell_1rw
* cell instance $13362 m0 *1 179.07,70.98
X$13362 574 52 575 644 645 cell_1rw
* cell instance $13363 m0 *1 179.775,70.98
X$13363 576 52 577 644 645 cell_1rw
* cell instance $13364 m0 *1 180.48,70.98
X$13364 578 52 579 644 645 cell_1rw
* cell instance $13365 r0 *1 0.705,70.98
X$13365 67 53 68 644 645 cell_1rw
* cell instance $13366 r0 *1 0,70.98
X$13366 65 53 66 644 645 cell_1rw
* cell instance $13367 r0 *1 1.41,70.98
X$13367 69 53 70 644 645 cell_1rw
* cell instance $13368 r0 *1 2.115,70.98
X$13368 71 53 72 644 645 cell_1rw
* cell instance $13369 r0 *1 2.82,70.98
X$13369 73 53 74 644 645 cell_1rw
* cell instance $13370 r0 *1 3.525,70.98
X$13370 75 53 76 644 645 cell_1rw
* cell instance $13371 r0 *1 4.23,70.98
X$13371 77 53 78 644 645 cell_1rw
* cell instance $13372 r0 *1 4.935,70.98
X$13372 79 53 80 644 645 cell_1rw
* cell instance $13373 r0 *1 5.64,70.98
X$13373 81 53 82 644 645 cell_1rw
* cell instance $13374 r0 *1 6.345,70.98
X$13374 83 53 84 644 645 cell_1rw
* cell instance $13375 r0 *1 7.05,70.98
X$13375 85 53 86 644 645 cell_1rw
* cell instance $13376 r0 *1 7.755,70.98
X$13376 87 53 88 644 645 cell_1rw
* cell instance $13377 r0 *1 8.46,70.98
X$13377 89 53 90 644 645 cell_1rw
* cell instance $13378 r0 *1 9.165,70.98
X$13378 91 53 92 644 645 cell_1rw
* cell instance $13379 r0 *1 9.87,70.98
X$13379 93 53 94 644 645 cell_1rw
* cell instance $13380 r0 *1 10.575,70.98
X$13380 95 53 96 644 645 cell_1rw
* cell instance $13381 r0 *1 11.28,70.98
X$13381 97 53 98 644 645 cell_1rw
* cell instance $13382 r0 *1 11.985,70.98
X$13382 99 53 100 644 645 cell_1rw
* cell instance $13383 r0 *1 12.69,70.98
X$13383 101 53 102 644 645 cell_1rw
* cell instance $13384 r0 *1 13.395,70.98
X$13384 103 53 104 644 645 cell_1rw
* cell instance $13385 r0 *1 14.1,70.98
X$13385 105 53 106 644 645 cell_1rw
* cell instance $13386 r0 *1 14.805,70.98
X$13386 107 53 108 644 645 cell_1rw
* cell instance $13387 r0 *1 15.51,70.98
X$13387 109 53 110 644 645 cell_1rw
* cell instance $13388 r0 *1 16.215,70.98
X$13388 111 53 112 644 645 cell_1rw
* cell instance $13389 r0 *1 16.92,70.98
X$13389 113 53 114 644 645 cell_1rw
* cell instance $13390 r0 *1 17.625,70.98
X$13390 115 53 116 644 645 cell_1rw
* cell instance $13391 r0 *1 18.33,70.98
X$13391 117 53 118 644 645 cell_1rw
* cell instance $13392 r0 *1 19.035,70.98
X$13392 119 53 120 644 645 cell_1rw
* cell instance $13393 r0 *1 19.74,70.98
X$13393 121 53 122 644 645 cell_1rw
* cell instance $13394 r0 *1 20.445,70.98
X$13394 123 53 124 644 645 cell_1rw
* cell instance $13395 r0 *1 21.15,70.98
X$13395 125 53 126 644 645 cell_1rw
* cell instance $13396 r0 *1 21.855,70.98
X$13396 127 53 128 644 645 cell_1rw
* cell instance $13397 r0 *1 22.56,70.98
X$13397 129 53 130 644 645 cell_1rw
* cell instance $13398 r0 *1 23.265,70.98
X$13398 131 53 132 644 645 cell_1rw
* cell instance $13399 r0 *1 23.97,70.98
X$13399 133 53 134 644 645 cell_1rw
* cell instance $13400 r0 *1 24.675,70.98
X$13400 135 53 136 644 645 cell_1rw
* cell instance $13401 r0 *1 25.38,70.98
X$13401 137 53 138 644 645 cell_1rw
* cell instance $13402 r0 *1 26.085,70.98
X$13402 139 53 140 644 645 cell_1rw
* cell instance $13403 r0 *1 26.79,70.98
X$13403 141 53 142 644 645 cell_1rw
* cell instance $13404 r0 *1 27.495,70.98
X$13404 143 53 144 644 645 cell_1rw
* cell instance $13405 r0 *1 28.2,70.98
X$13405 145 53 146 644 645 cell_1rw
* cell instance $13406 r0 *1 28.905,70.98
X$13406 147 53 148 644 645 cell_1rw
* cell instance $13407 r0 *1 29.61,70.98
X$13407 149 53 150 644 645 cell_1rw
* cell instance $13408 r0 *1 30.315,70.98
X$13408 151 53 152 644 645 cell_1rw
* cell instance $13409 r0 *1 31.02,70.98
X$13409 153 53 154 644 645 cell_1rw
* cell instance $13410 r0 *1 31.725,70.98
X$13410 155 53 156 644 645 cell_1rw
* cell instance $13411 r0 *1 32.43,70.98
X$13411 157 53 158 644 645 cell_1rw
* cell instance $13412 r0 *1 33.135,70.98
X$13412 159 53 160 644 645 cell_1rw
* cell instance $13413 r0 *1 33.84,70.98
X$13413 161 53 162 644 645 cell_1rw
* cell instance $13414 r0 *1 34.545,70.98
X$13414 163 53 164 644 645 cell_1rw
* cell instance $13415 r0 *1 35.25,70.98
X$13415 165 53 166 644 645 cell_1rw
* cell instance $13416 r0 *1 35.955,70.98
X$13416 167 53 168 644 645 cell_1rw
* cell instance $13417 r0 *1 36.66,70.98
X$13417 169 53 170 644 645 cell_1rw
* cell instance $13418 r0 *1 37.365,70.98
X$13418 171 53 172 644 645 cell_1rw
* cell instance $13419 r0 *1 38.07,70.98
X$13419 173 53 174 644 645 cell_1rw
* cell instance $13420 r0 *1 38.775,70.98
X$13420 175 53 176 644 645 cell_1rw
* cell instance $13421 r0 *1 39.48,70.98
X$13421 177 53 178 644 645 cell_1rw
* cell instance $13422 r0 *1 40.185,70.98
X$13422 179 53 180 644 645 cell_1rw
* cell instance $13423 r0 *1 40.89,70.98
X$13423 181 53 182 644 645 cell_1rw
* cell instance $13424 r0 *1 41.595,70.98
X$13424 183 53 184 644 645 cell_1rw
* cell instance $13425 r0 *1 42.3,70.98
X$13425 185 53 186 644 645 cell_1rw
* cell instance $13426 r0 *1 43.005,70.98
X$13426 187 53 188 644 645 cell_1rw
* cell instance $13427 r0 *1 43.71,70.98
X$13427 189 53 190 644 645 cell_1rw
* cell instance $13428 r0 *1 44.415,70.98
X$13428 191 53 192 644 645 cell_1rw
* cell instance $13429 r0 *1 45.12,70.98
X$13429 193 53 194 644 645 cell_1rw
* cell instance $13430 r0 *1 45.825,70.98
X$13430 195 53 196 644 645 cell_1rw
* cell instance $13431 r0 *1 46.53,70.98
X$13431 197 53 198 644 645 cell_1rw
* cell instance $13432 r0 *1 47.235,70.98
X$13432 199 53 200 644 645 cell_1rw
* cell instance $13433 r0 *1 47.94,70.98
X$13433 201 53 202 644 645 cell_1rw
* cell instance $13434 r0 *1 48.645,70.98
X$13434 203 53 204 644 645 cell_1rw
* cell instance $13435 r0 *1 49.35,70.98
X$13435 205 53 206 644 645 cell_1rw
* cell instance $13436 r0 *1 50.055,70.98
X$13436 207 53 208 644 645 cell_1rw
* cell instance $13437 r0 *1 50.76,70.98
X$13437 209 53 210 644 645 cell_1rw
* cell instance $13438 r0 *1 51.465,70.98
X$13438 211 53 212 644 645 cell_1rw
* cell instance $13439 r0 *1 52.17,70.98
X$13439 213 53 214 644 645 cell_1rw
* cell instance $13440 r0 *1 52.875,70.98
X$13440 215 53 216 644 645 cell_1rw
* cell instance $13441 r0 *1 53.58,70.98
X$13441 217 53 218 644 645 cell_1rw
* cell instance $13442 r0 *1 54.285,70.98
X$13442 219 53 220 644 645 cell_1rw
* cell instance $13443 r0 *1 54.99,70.98
X$13443 221 53 222 644 645 cell_1rw
* cell instance $13444 r0 *1 55.695,70.98
X$13444 223 53 224 644 645 cell_1rw
* cell instance $13445 r0 *1 56.4,70.98
X$13445 225 53 226 644 645 cell_1rw
* cell instance $13446 r0 *1 57.105,70.98
X$13446 227 53 228 644 645 cell_1rw
* cell instance $13447 r0 *1 57.81,70.98
X$13447 229 53 230 644 645 cell_1rw
* cell instance $13448 r0 *1 58.515,70.98
X$13448 231 53 232 644 645 cell_1rw
* cell instance $13449 r0 *1 59.22,70.98
X$13449 233 53 234 644 645 cell_1rw
* cell instance $13450 r0 *1 59.925,70.98
X$13450 235 53 236 644 645 cell_1rw
* cell instance $13451 r0 *1 60.63,70.98
X$13451 237 53 238 644 645 cell_1rw
* cell instance $13452 r0 *1 61.335,70.98
X$13452 239 53 240 644 645 cell_1rw
* cell instance $13453 r0 *1 62.04,70.98
X$13453 241 53 242 644 645 cell_1rw
* cell instance $13454 r0 *1 62.745,70.98
X$13454 243 53 244 644 645 cell_1rw
* cell instance $13455 r0 *1 63.45,70.98
X$13455 245 53 246 644 645 cell_1rw
* cell instance $13456 r0 *1 64.155,70.98
X$13456 247 53 248 644 645 cell_1rw
* cell instance $13457 r0 *1 64.86,70.98
X$13457 249 53 250 644 645 cell_1rw
* cell instance $13458 r0 *1 65.565,70.98
X$13458 251 53 252 644 645 cell_1rw
* cell instance $13459 r0 *1 66.27,70.98
X$13459 253 53 254 644 645 cell_1rw
* cell instance $13460 r0 *1 66.975,70.98
X$13460 255 53 256 644 645 cell_1rw
* cell instance $13461 r0 *1 67.68,70.98
X$13461 257 53 258 644 645 cell_1rw
* cell instance $13462 r0 *1 68.385,70.98
X$13462 259 53 260 644 645 cell_1rw
* cell instance $13463 r0 *1 69.09,70.98
X$13463 261 53 262 644 645 cell_1rw
* cell instance $13464 r0 *1 69.795,70.98
X$13464 263 53 264 644 645 cell_1rw
* cell instance $13465 r0 *1 70.5,70.98
X$13465 265 53 266 644 645 cell_1rw
* cell instance $13466 r0 *1 71.205,70.98
X$13466 267 53 268 644 645 cell_1rw
* cell instance $13467 r0 *1 71.91,70.98
X$13467 269 53 270 644 645 cell_1rw
* cell instance $13468 r0 *1 72.615,70.98
X$13468 271 53 272 644 645 cell_1rw
* cell instance $13469 r0 *1 73.32,70.98
X$13469 273 53 274 644 645 cell_1rw
* cell instance $13470 r0 *1 74.025,70.98
X$13470 275 53 276 644 645 cell_1rw
* cell instance $13471 r0 *1 74.73,70.98
X$13471 277 53 278 644 645 cell_1rw
* cell instance $13472 r0 *1 75.435,70.98
X$13472 279 53 280 644 645 cell_1rw
* cell instance $13473 r0 *1 76.14,70.98
X$13473 281 53 282 644 645 cell_1rw
* cell instance $13474 r0 *1 76.845,70.98
X$13474 283 53 284 644 645 cell_1rw
* cell instance $13475 r0 *1 77.55,70.98
X$13475 285 53 286 644 645 cell_1rw
* cell instance $13476 r0 *1 78.255,70.98
X$13476 287 53 288 644 645 cell_1rw
* cell instance $13477 r0 *1 78.96,70.98
X$13477 289 53 290 644 645 cell_1rw
* cell instance $13478 r0 *1 79.665,70.98
X$13478 291 53 292 644 645 cell_1rw
* cell instance $13479 r0 *1 80.37,70.98
X$13479 293 53 294 644 645 cell_1rw
* cell instance $13480 r0 *1 81.075,70.98
X$13480 295 53 296 644 645 cell_1rw
* cell instance $13481 r0 *1 81.78,70.98
X$13481 297 53 298 644 645 cell_1rw
* cell instance $13482 r0 *1 82.485,70.98
X$13482 299 53 300 644 645 cell_1rw
* cell instance $13483 r0 *1 83.19,70.98
X$13483 301 53 302 644 645 cell_1rw
* cell instance $13484 r0 *1 83.895,70.98
X$13484 303 53 304 644 645 cell_1rw
* cell instance $13485 r0 *1 84.6,70.98
X$13485 305 53 306 644 645 cell_1rw
* cell instance $13486 r0 *1 85.305,70.98
X$13486 307 53 308 644 645 cell_1rw
* cell instance $13487 r0 *1 86.01,70.98
X$13487 309 53 310 644 645 cell_1rw
* cell instance $13488 r0 *1 86.715,70.98
X$13488 311 53 312 644 645 cell_1rw
* cell instance $13489 r0 *1 87.42,70.98
X$13489 313 53 314 644 645 cell_1rw
* cell instance $13490 r0 *1 88.125,70.98
X$13490 315 53 316 644 645 cell_1rw
* cell instance $13491 r0 *1 88.83,70.98
X$13491 317 53 318 644 645 cell_1rw
* cell instance $13492 r0 *1 89.535,70.98
X$13492 319 53 320 644 645 cell_1rw
* cell instance $13493 r0 *1 90.24,70.98
X$13493 321 53 323 644 645 cell_1rw
* cell instance $13494 r0 *1 90.945,70.98
X$13494 324 53 325 644 645 cell_1rw
* cell instance $13495 r0 *1 91.65,70.98
X$13495 326 53 327 644 645 cell_1rw
* cell instance $13496 r0 *1 92.355,70.98
X$13496 328 53 329 644 645 cell_1rw
* cell instance $13497 r0 *1 93.06,70.98
X$13497 330 53 331 644 645 cell_1rw
* cell instance $13498 r0 *1 93.765,70.98
X$13498 332 53 333 644 645 cell_1rw
* cell instance $13499 r0 *1 94.47,70.98
X$13499 334 53 335 644 645 cell_1rw
* cell instance $13500 r0 *1 95.175,70.98
X$13500 336 53 337 644 645 cell_1rw
* cell instance $13501 r0 *1 95.88,70.98
X$13501 338 53 339 644 645 cell_1rw
* cell instance $13502 r0 *1 96.585,70.98
X$13502 340 53 341 644 645 cell_1rw
* cell instance $13503 r0 *1 97.29,70.98
X$13503 342 53 343 644 645 cell_1rw
* cell instance $13504 r0 *1 97.995,70.98
X$13504 344 53 345 644 645 cell_1rw
* cell instance $13505 r0 *1 98.7,70.98
X$13505 346 53 347 644 645 cell_1rw
* cell instance $13506 r0 *1 99.405,70.98
X$13506 348 53 349 644 645 cell_1rw
* cell instance $13507 r0 *1 100.11,70.98
X$13507 350 53 351 644 645 cell_1rw
* cell instance $13508 r0 *1 100.815,70.98
X$13508 352 53 353 644 645 cell_1rw
* cell instance $13509 r0 *1 101.52,70.98
X$13509 354 53 355 644 645 cell_1rw
* cell instance $13510 r0 *1 102.225,70.98
X$13510 356 53 357 644 645 cell_1rw
* cell instance $13511 r0 *1 102.93,70.98
X$13511 358 53 359 644 645 cell_1rw
* cell instance $13512 r0 *1 103.635,70.98
X$13512 360 53 361 644 645 cell_1rw
* cell instance $13513 r0 *1 104.34,70.98
X$13513 362 53 363 644 645 cell_1rw
* cell instance $13514 r0 *1 105.045,70.98
X$13514 364 53 365 644 645 cell_1rw
* cell instance $13515 r0 *1 105.75,70.98
X$13515 366 53 367 644 645 cell_1rw
* cell instance $13516 r0 *1 106.455,70.98
X$13516 368 53 369 644 645 cell_1rw
* cell instance $13517 r0 *1 107.16,70.98
X$13517 370 53 371 644 645 cell_1rw
* cell instance $13518 r0 *1 107.865,70.98
X$13518 372 53 373 644 645 cell_1rw
* cell instance $13519 r0 *1 108.57,70.98
X$13519 374 53 375 644 645 cell_1rw
* cell instance $13520 r0 *1 109.275,70.98
X$13520 376 53 377 644 645 cell_1rw
* cell instance $13521 r0 *1 109.98,70.98
X$13521 378 53 379 644 645 cell_1rw
* cell instance $13522 r0 *1 110.685,70.98
X$13522 380 53 381 644 645 cell_1rw
* cell instance $13523 r0 *1 111.39,70.98
X$13523 382 53 383 644 645 cell_1rw
* cell instance $13524 r0 *1 112.095,70.98
X$13524 384 53 385 644 645 cell_1rw
* cell instance $13525 r0 *1 112.8,70.98
X$13525 386 53 387 644 645 cell_1rw
* cell instance $13526 r0 *1 113.505,70.98
X$13526 388 53 389 644 645 cell_1rw
* cell instance $13527 r0 *1 114.21,70.98
X$13527 390 53 391 644 645 cell_1rw
* cell instance $13528 r0 *1 114.915,70.98
X$13528 392 53 393 644 645 cell_1rw
* cell instance $13529 r0 *1 115.62,70.98
X$13529 394 53 395 644 645 cell_1rw
* cell instance $13530 r0 *1 116.325,70.98
X$13530 396 53 397 644 645 cell_1rw
* cell instance $13531 r0 *1 117.03,70.98
X$13531 398 53 399 644 645 cell_1rw
* cell instance $13532 r0 *1 117.735,70.98
X$13532 400 53 401 644 645 cell_1rw
* cell instance $13533 r0 *1 118.44,70.98
X$13533 402 53 403 644 645 cell_1rw
* cell instance $13534 r0 *1 119.145,70.98
X$13534 404 53 405 644 645 cell_1rw
* cell instance $13535 r0 *1 119.85,70.98
X$13535 406 53 407 644 645 cell_1rw
* cell instance $13536 r0 *1 120.555,70.98
X$13536 408 53 409 644 645 cell_1rw
* cell instance $13537 r0 *1 121.26,70.98
X$13537 410 53 411 644 645 cell_1rw
* cell instance $13538 r0 *1 121.965,70.98
X$13538 412 53 413 644 645 cell_1rw
* cell instance $13539 r0 *1 122.67,70.98
X$13539 414 53 415 644 645 cell_1rw
* cell instance $13540 r0 *1 123.375,70.98
X$13540 416 53 417 644 645 cell_1rw
* cell instance $13541 r0 *1 124.08,70.98
X$13541 418 53 419 644 645 cell_1rw
* cell instance $13542 r0 *1 124.785,70.98
X$13542 420 53 421 644 645 cell_1rw
* cell instance $13543 r0 *1 125.49,70.98
X$13543 422 53 423 644 645 cell_1rw
* cell instance $13544 r0 *1 126.195,70.98
X$13544 424 53 425 644 645 cell_1rw
* cell instance $13545 r0 *1 126.9,70.98
X$13545 426 53 427 644 645 cell_1rw
* cell instance $13546 r0 *1 127.605,70.98
X$13546 428 53 429 644 645 cell_1rw
* cell instance $13547 r0 *1 128.31,70.98
X$13547 430 53 431 644 645 cell_1rw
* cell instance $13548 r0 *1 129.015,70.98
X$13548 432 53 433 644 645 cell_1rw
* cell instance $13549 r0 *1 129.72,70.98
X$13549 434 53 435 644 645 cell_1rw
* cell instance $13550 r0 *1 130.425,70.98
X$13550 436 53 437 644 645 cell_1rw
* cell instance $13551 r0 *1 131.13,70.98
X$13551 438 53 439 644 645 cell_1rw
* cell instance $13552 r0 *1 131.835,70.98
X$13552 440 53 441 644 645 cell_1rw
* cell instance $13553 r0 *1 132.54,70.98
X$13553 442 53 443 644 645 cell_1rw
* cell instance $13554 r0 *1 133.245,70.98
X$13554 444 53 445 644 645 cell_1rw
* cell instance $13555 r0 *1 133.95,70.98
X$13555 446 53 447 644 645 cell_1rw
* cell instance $13556 r0 *1 134.655,70.98
X$13556 448 53 449 644 645 cell_1rw
* cell instance $13557 r0 *1 135.36,70.98
X$13557 450 53 451 644 645 cell_1rw
* cell instance $13558 r0 *1 136.065,70.98
X$13558 452 53 453 644 645 cell_1rw
* cell instance $13559 r0 *1 136.77,70.98
X$13559 454 53 455 644 645 cell_1rw
* cell instance $13560 r0 *1 137.475,70.98
X$13560 456 53 457 644 645 cell_1rw
* cell instance $13561 r0 *1 138.18,70.98
X$13561 458 53 459 644 645 cell_1rw
* cell instance $13562 r0 *1 138.885,70.98
X$13562 460 53 461 644 645 cell_1rw
* cell instance $13563 r0 *1 139.59,70.98
X$13563 462 53 463 644 645 cell_1rw
* cell instance $13564 r0 *1 140.295,70.98
X$13564 464 53 465 644 645 cell_1rw
* cell instance $13565 r0 *1 141,70.98
X$13565 466 53 467 644 645 cell_1rw
* cell instance $13566 r0 *1 141.705,70.98
X$13566 468 53 469 644 645 cell_1rw
* cell instance $13567 r0 *1 142.41,70.98
X$13567 470 53 471 644 645 cell_1rw
* cell instance $13568 r0 *1 143.115,70.98
X$13568 472 53 473 644 645 cell_1rw
* cell instance $13569 r0 *1 143.82,70.98
X$13569 474 53 475 644 645 cell_1rw
* cell instance $13570 r0 *1 144.525,70.98
X$13570 476 53 477 644 645 cell_1rw
* cell instance $13571 r0 *1 145.23,70.98
X$13571 478 53 479 644 645 cell_1rw
* cell instance $13572 r0 *1 145.935,70.98
X$13572 480 53 481 644 645 cell_1rw
* cell instance $13573 r0 *1 146.64,70.98
X$13573 482 53 483 644 645 cell_1rw
* cell instance $13574 r0 *1 147.345,70.98
X$13574 484 53 485 644 645 cell_1rw
* cell instance $13575 r0 *1 148.05,70.98
X$13575 486 53 487 644 645 cell_1rw
* cell instance $13576 r0 *1 148.755,70.98
X$13576 488 53 489 644 645 cell_1rw
* cell instance $13577 r0 *1 149.46,70.98
X$13577 490 53 491 644 645 cell_1rw
* cell instance $13578 r0 *1 150.165,70.98
X$13578 492 53 493 644 645 cell_1rw
* cell instance $13579 r0 *1 150.87,70.98
X$13579 494 53 495 644 645 cell_1rw
* cell instance $13580 r0 *1 151.575,70.98
X$13580 496 53 497 644 645 cell_1rw
* cell instance $13581 r0 *1 152.28,70.98
X$13581 498 53 499 644 645 cell_1rw
* cell instance $13582 r0 *1 152.985,70.98
X$13582 500 53 501 644 645 cell_1rw
* cell instance $13583 r0 *1 153.69,70.98
X$13583 502 53 503 644 645 cell_1rw
* cell instance $13584 r0 *1 154.395,70.98
X$13584 504 53 505 644 645 cell_1rw
* cell instance $13585 r0 *1 155.1,70.98
X$13585 506 53 507 644 645 cell_1rw
* cell instance $13586 r0 *1 155.805,70.98
X$13586 508 53 509 644 645 cell_1rw
* cell instance $13587 r0 *1 156.51,70.98
X$13587 510 53 511 644 645 cell_1rw
* cell instance $13588 r0 *1 157.215,70.98
X$13588 512 53 513 644 645 cell_1rw
* cell instance $13589 r0 *1 157.92,70.98
X$13589 514 53 515 644 645 cell_1rw
* cell instance $13590 r0 *1 158.625,70.98
X$13590 516 53 517 644 645 cell_1rw
* cell instance $13591 r0 *1 159.33,70.98
X$13591 518 53 519 644 645 cell_1rw
* cell instance $13592 r0 *1 160.035,70.98
X$13592 520 53 521 644 645 cell_1rw
* cell instance $13593 r0 *1 160.74,70.98
X$13593 522 53 523 644 645 cell_1rw
* cell instance $13594 r0 *1 161.445,70.98
X$13594 524 53 525 644 645 cell_1rw
* cell instance $13595 r0 *1 162.15,70.98
X$13595 526 53 527 644 645 cell_1rw
* cell instance $13596 r0 *1 162.855,70.98
X$13596 528 53 529 644 645 cell_1rw
* cell instance $13597 r0 *1 163.56,70.98
X$13597 530 53 531 644 645 cell_1rw
* cell instance $13598 r0 *1 164.265,70.98
X$13598 532 53 533 644 645 cell_1rw
* cell instance $13599 r0 *1 164.97,70.98
X$13599 534 53 535 644 645 cell_1rw
* cell instance $13600 r0 *1 165.675,70.98
X$13600 536 53 537 644 645 cell_1rw
* cell instance $13601 r0 *1 166.38,70.98
X$13601 538 53 539 644 645 cell_1rw
* cell instance $13602 r0 *1 167.085,70.98
X$13602 540 53 541 644 645 cell_1rw
* cell instance $13603 r0 *1 167.79,70.98
X$13603 542 53 543 644 645 cell_1rw
* cell instance $13604 r0 *1 168.495,70.98
X$13604 544 53 545 644 645 cell_1rw
* cell instance $13605 r0 *1 169.2,70.98
X$13605 546 53 547 644 645 cell_1rw
* cell instance $13606 r0 *1 169.905,70.98
X$13606 548 53 549 644 645 cell_1rw
* cell instance $13607 r0 *1 170.61,70.98
X$13607 550 53 551 644 645 cell_1rw
* cell instance $13608 r0 *1 171.315,70.98
X$13608 552 53 553 644 645 cell_1rw
* cell instance $13609 r0 *1 172.02,70.98
X$13609 554 53 555 644 645 cell_1rw
* cell instance $13610 r0 *1 172.725,70.98
X$13610 556 53 557 644 645 cell_1rw
* cell instance $13611 r0 *1 173.43,70.98
X$13611 558 53 559 644 645 cell_1rw
* cell instance $13612 r0 *1 174.135,70.98
X$13612 560 53 561 644 645 cell_1rw
* cell instance $13613 r0 *1 174.84,70.98
X$13613 562 53 563 644 645 cell_1rw
* cell instance $13614 r0 *1 175.545,70.98
X$13614 564 53 565 644 645 cell_1rw
* cell instance $13615 r0 *1 176.25,70.98
X$13615 566 53 567 644 645 cell_1rw
* cell instance $13616 r0 *1 176.955,70.98
X$13616 568 53 569 644 645 cell_1rw
* cell instance $13617 r0 *1 177.66,70.98
X$13617 570 53 571 644 645 cell_1rw
* cell instance $13618 r0 *1 178.365,70.98
X$13618 572 53 573 644 645 cell_1rw
* cell instance $13619 r0 *1 179.07,70.98
X$13619 574 53 575 644 645 cell_1rw
* cell instance $13620 r0 *1 179.775,70.98
X$13620 576 53 577 644 645 cell_1rw
* cell instance $13621 r0 *1 180.48,70.98
X$13621 578 53 579 644 645 cell_1rw
* cell instance $13622 m0 *1 0.705,73.71
X$13622 67 54 68 644 645 cell_1rw
* cell instance $13623 m0 *1 0,73.71
X$13623 65 54 66 644 645 cell_1rw
* cell instance $13624 m0 *1 1.41,73.71
X$13624 69 54 70 644 645 cell_1rw
* cell instance $13625 m0 *1 2.115,73.71
X$13625 71 54 72 644 645 cell_1rw
* cell instance $13626 m0 *1 2.82,73.71
X$13626 73 54 74 644 645 cell_1rw
* cell instance $13627 m0 *1 3.525,73.71
X$13627 75 54 76 644 645 cell_1rw
* cell instance $13628 m0 *1 4.23,73.71
X$13628 77 54 78 644 645 cell_1rw
* cell instance $13629 m0 *1 4.935,73.71
X$13629 79 54 80 644 645 cell_1rw
* cell instance $13630 m0 *1 5.64,73.71
X$13630 81 54 82 644 645 cell_1rw
* cell instance $13631 m0 *1 6.345,73.71
X$13631 83 54 84 644 645 cell_1rw
* cell instance $13632 m0 *1 7.05,73.71
X$13632 85 54 86 644 645 cell_1rw
* cell instance $13633 m0 *1 7.755,73.71
X$13633 87 54 88 644 645 cell_1rw
* cell instance $13634 m0 *1 8.46,73.71
X$13634 89 54 90 644 645 cell_1rw
* cell instance $13635 m0 *1 9.165,73.71
X$13635 91 54 92 644 645 cell_1rw
* cell instance $13636 m0 *1 9.87,73.71
X$13636 93 54 94 644 645 cell_1rw
* cell instance $13637 m0 *1 10.575,73.71
X$13637 95 54 96 644 645 cell_1rw
* cell instance $13638 m0 *1 11.28,73.71
X$13638 97 54 98 644 645 cell_1rw
* cell instance $13639 m0 *1 11.985,73.71
X$13639 99 54 100 644 645 cell_1rw
* cell instance $13640 m0 *1 12.69,73.71
X$13640 101 54 102 644 645 cell_1rw
* cell instance $13641 m0 *1 13.395,73.71
X$13641 103 54 104 644 645 cell_1rw
* cell instance $13642 m0 *1 14.1,73.71
X$13642 105 54 106 644 645 cell_1rw
* cell instance $13643 m0 *1 14.805,73.71
X$13643 107 54 108 644 645 cell_1rw
* cell instance $13644 m0 *1 15.51,73.71
X$13644 109 54 110 644 645 cell_1rw
* cell instance $13645 m0 *1 16.215,73.71
X$13645 111 54 112 644 645 cell_1rw
* cell instance $13646 m0 *1 16.92,73.71
X$13646 113 54 114 644 645 cell_1rw
* cell instance $13647 m0 *1 17.625,73.71
X$13647 115 54 116 644 645 cell_1rw
* cell instance $13648 m0 *1 18.33,73.71
X$13648 117 54 118 644 645 cell_1rw
* cell instance $13649 m0 *1 19.035,73.71
X$13649 119 54 120 644 645 cell_1rw
* cell instance $13650 m0 *1 19.74,73.71
X$13650 121 54 122 644 645 cell_1rw
* cell instance $13651 m0 *1 20.445,73.71
X$13651 123 54 124 644 645 cell_1rw
* cell instance $13652 m0 *1 21.15,73.71
X$13652 125 54 126 644 645 cell_1rw
* cell instance $13653 m0 *1 21.855,73.71
X$13653 127 54 128 644 645 cell_1rw
* cell instance $13654 m0 *1 22.56,73.71
X$13654 129 54 130 644 645 cell_1rw
* cell instance $13655 m0 *1 23.265,73.71
X$13655 131 54 132 644 645 cell_1rw
* cell instance $13656 m0 *1 23.97,73.71
X$13656 133 54 134 644 645 cell_1rw
* cell instance $13657 m0 *1 24.675,73.71
X$13657 135 54 136 644 645 cell_1rw
* cell instance $13658 m0 *1 25.38,73.71
X$13658 137 54 138 644 645 cell_1rw
* cell instance $13659 m0 *1 26.085,73.71
X$13659 139 54 140 644 645 cell_1rw
* cell instance $13660 m0 *1 26.79,73.71
X$13660 141 54 142 644 645 cell_1rw
* cell instance $13661 m0 *1 27.495,73.71
X$13661 143 54 144 644 645 cell_1rw
* cell instance $13662 m0 *1 28.2,73.71
X$13662 145 54 146 644 645 cell_1rw
* cell instance $13663 m0 *1 28.905,73.71
X$13663 147 54 148 644 645 cell_1rw
* cell instance $13664 m0 *1 29.61,73.71
X$13664 149 54 150 644 645 cell_1rw
* cell instance $13665 m0 *1 30.315,73.71
X$13665 151 54 152 644 645 cell_1rw
* cell instance $13666 m0 *1 31.02,73.71
X$13666 153 54 154 644 645 cell_1rw
* cell instance $13667 m0 *1 31.725,73.71
X$13667 155 54 156 644 645 cell_1rw
* cell instance $13668 m0 *1 32.43,73.71
X$13668 157 54 158 644 645 cell_1rw
* cell instance $13669 m0 *1 33.135,73.71
X$13669 159 54 160 644 645 cell_1rw
* cell instance $13670 m0 *1 33.84,73.71
X$13670 161 54 162 644 645 cell_1rw
* cell instance $13671 m0 *1 34.545,73.71
X$13671 163 54 164 644 645 cell_1rw
* cell instance $13672 m0 *1 35.25,73.71
X$13672 165 54 166 644 645 cell_1rw
* cell instance $13673 m0 *1 35.955,73.71
X$13673 167 54 168 644 645 cell_1rw
* cell instance $13674 m0 *1 36.66,73.71
X$13674 169 54 170 644 645 cell_1rw
* cell instance $13675 m0 *1 37.365,73.71
X$13675 171 54 172 644 645 cell_1rw
* cell instance $13676 m0 *1 38.07,73.71
X$13676 173 54 174 644 645 cell_1rw
* cell instance $13677 m0 *1 38.775,73.71
X$13677 175 54 176 644 645 cell_1rw
* cell instance $13678 m0 *1 39.48,73.71
X$13678 177 54 178 644 645 cell_1rw
* cell instance $13679 m0 *1 40.185,73.71
X$13679 179 54 180 644 645 cell_1rw
* cell instance $13680 m0 *1 40.89,73.71
X$13680 181 54 182 644 645 cell_1rw
* cell instance $13681 m0 *1 41.595,73.71
X$13681 183 54 184 644 645 cell_1rw
* cell instance $13682 m0 *1 42.3,73.71
X$13682 185 54 186 644 645 cell_1rw
* cell instance $13683 m0 *1 43.005,73.71
X$13683 187 54 188 644 645 cell_1rw
* cell instance $13684 m0 *1 43.71,73.71
X$13684 189 54 190 644 645 cell_1rw
* cell instance $13685 m0 *1 44.415,73.71
X$13685 191 54 192 644 645 cell_1rw
* cell instance $13686 m0 *1 45.12,73.71
X$13686 193 54 194 644 645 cell_1rw
* cell instance $13687 m0 *1 45.825,73.71
X$13687 195 54 196 644 645 cell_1rw
* cell instance $13688 m0 *1 46.53,73.71
X$13688 197 54 198 644 645 cell_1rw
* cell instance $13689 m0 *1 47.235,73.71
X$13689 199 54 200 644 645 cell_1rw
* cell instance $13690 m0 *1 47.94,73.71
X$13690 201 54 202 644 645 cell_1rw
* cell instance $13691 m0 *1 48.645,73.71
X$13691 203 54 204 644 645 cell_1rw
* cell instance $13692 m0 *1 49.35,73.71
X$13692 205 54 206 644 645 cell_1rw
* cell instance $13693 m0 *1 50.055,73.71
X$13693 207 54 208 644 645 cell_1rw
* cell instance $13694 m0 *1 50.76,73.71
X$13694 209 54 210 644 645 cell_1rw
* cell instance $13695 m0 *1 51.465,73.71
X$13695 211 54 212 644 645 cell_1rw
* cell instance $13696 m0 *1 52.17,73.71
X$13696 213 54 214 644 645 cell_1rw
* cell instance $13697 m0 *1 52.875,73.71
X$13697 215 54 216 644 645 cell_1rw
* cell instance $13698 m0 *1 53.58,73.71
X$13698 217 54 218 644 645 cell_1rw
* cell instance $13699 m0 *1 54.285,73.71
X$13699 219 54 220 644 645 cell_1rw
* cell instance $13700 m0 *1 54.99,73.71
X$13700 221 54 222 644 645 cell_1rw
* cell instance $13701 m0 *1 55.695,73.71
X$13701 223 54 224 644 645 cell_1rw
* cell instance $13702 m0 *1 56.4,73.71
X$13702 225 54 226 644 645 cell_1rw
* cell instance $13703 m0 *1 57.105,73.71
X$13703 227 54 228 644 645 cell_1rw
* cell instance $13704 m0 *1 57.81,73.71
X$13704 229 54 230 644 645 cell_1rw
* cell instance $13705 m0 *1 58.515,73.71
X$13705 231 54 232 644 645 cell_1rw
* cell instance $13706 m0 *1 59.22,73.71
X$13706 233 54 234 644 645 cell_1rw
* cell instance $13707 m0 *1 59.925,73.71
X$13707 235 54 236 644 645 cell_1rw
* cell instance $13708 m0 *1 60.63,73.71
X$13708 237 54 238 644 645 cell_1rw
* cell instance $13709 m0 *1 61.335,73.71
X$13709 239 54 240 644 645 cell_1rw
* cell instance $13710 m0 *1 62.04,73.71
X$13710 241 54 242 644 645 cell_1rw
* cell instance $13711 m0 *1 62.745,73.71
X$13711 243 54 244 644 645 cell_1rw
* cell instance $13712 m0 *1 63.45,73.71
X$13712 245 54 246 644 645 cell_1rw
* cell instance $13713 m0 *1 64.155,73.71
X$13713 247 54 248 644 645 cell_1rw
* cell instance $13714 m0 *1 64.86,73.71
X$13714 249 54 250 644 645 cell_1rw
* cell instance $13715 m0 *1 65.565,73.71
X$13715 251 54 252 644 645 cell_1rw
* cell instance $13716 m0 *1 66.27,73.71
X$13716 253 54 254 644 645 cell_1rw
* cell instance $13717 m0 *1 66.975,73.71
X$13717 255 54 256 644 645 cell_1rw
* cell instance $13718 m0 *1 67.68,73.71
X$13718 257 54 258 644 645 cell_1rw
* cell instance $13719 m0 *1 68.385,73.71
X$13719 259 54 260 644 645 cell_1rw
* cell instance $13720 m0 *1 69.09,73.71
X$13720 261 54 262 644 645 cell_1rw
* cell instance $13721 m0 *1 69.795,73.71
X$13721 263 54 264 644 645 cell_1rw
* cell instance $13722 m0 *1 70.5,73.71
X$13722 265 54 266 644 645 cell_1rw
* cell instance $13723 m0 *1 71.205,73.71
X$13723 267 54 268 644 645 cell_1rw
* cell instance $13724 m0 *1 71.91,73.71
X$13724 269 54 270 644 645 cell_1rw
* cell instance $13725 m0 *1 72.615,73.71
X$13725 271 54 272 644 645 cell_1rw
* cell instance $13726 m0 *1 73.32,73.71
X$13726 273 54 274 644 645 cell_1rw
* cell instance $13727 m0 *1 74.025,73.71
X$13727 275 54 276 644 645 cell_1rw
* cell instance $13728 m0 *1 74.73,73.71
X$13728 277 54 278 644 645 cell_1rw
* cell instance $13729 m0 *1 75.435,73.71
X$13729 279 54 280 644 645 cell_1rw
* cell instance $13730 m0 *1 76.14,73.71
X$13730 281 54 282 644 645 cell_1rw
* cell instance $13731 m0 *1 76.845,73.71
X$13731 283 54 284 644 645 cell_1rw
* cell instance $13732 m0 *1 77.55,73.71
X$13732 285 54 286 644 645 cell_1rw
* cell instance $13733 m0 *1 78.255,73.71
X$13733 287 54 288 644 645 cell_1rw
* cell instance $13734 m0 *1 78.96,73.71
X$13734 289 54 290 644 645 cell_1rw
* cell instance $13735 m0 *1 79.665,73.71
X$13735 291 54 292 644 645 cell_1rw
* cell instance $13736 m0 *1 80.37,73.71
X$13736 293 54 294 644 645 cell_1rw
* cell instance $13737 m0 *1 81.075,73.71
X$13737 295 54 296 644 645 cell_1rw
* cell instance $13738 m0 *1 81.78,73.71
X$13738 297 54 298 644 645 cell_1rw
* cell instance $13739 m0 *1 82.485,73.71
X$13739 299 54 300 644 645 cell_1rw
* cell instance $13740 m0 *1 83.19,73.71
X$13740 301 54 302 644 645 cell_1rw
* cell instance $13741 m0 *1 83.895,73.71
X$13741 303 54 304 644 645 cell_1rw
* cell instance $13742 m0 *1 84.6,73.71
X$13742 305 54 306 644 645 cell_1rw
* cell instance $13743 m0 *1 85.305,73.71
X$13743 307 54 308 644 645 cell_1rw
* cell instance $13744 m0 *1 86.01,73.71
X$13744 309 54 310 644 645 cell_1rw
* cell instance $13745 m0 *1 86.715,73.71
X$13745 311 54 312 644 645 cell_1rw
* cell instance $13746 m0 *1 87.42,73.71
X$13746 313 54 314 644 645 cell_1rw
* cell instance $13747 m0 *1 88.125,73.71
X$13747 315 54 316 644 645 cell_1rw
* cell instance $13748 m0 *1 88.83,73.71
X$13748 317 54 318 644 645 cell_1rw
* cell instance $13749 m0 *1 89.535,73.71
X$13749 319 54 320 644 645 cell_1rw
* cell instance $13750 m0 *1 90.24,73.71
X$13750 321 54 323 644 645 cell_1rw
* cell instance $13751 m0 *1 90.945,73.71
X$13751 324 54 325 644 645 cell_1rw
* cell instance $13752 m0 *1 91.65,73.71
X$13752 326 54 327 644 645 cell_1rw
* cell instance $13753 m0 *1 92.355,73.71
X$13753 328 54 329 644 645 cell_1rw
* cell instance $13754 m0 *1 93.06,73.71
X$13754 330 54 331 644 645 cell_1rw
* cell instance $13755 m0 *1 93.765,73.71
X$13755 332 54 333 644 645 cell_1rw
* cell instance $13756 m0 *1 94.47,73.71
X$13756 334 54 335 644 645 cell_1rw
* cell instance $13757 m0 *1 95.175,73.71
X$13757 336 54 337 644 645 cell_1rw
* cell instance $13758 m0 *1 95.88,73.71
X$13758 338 54 339 644 645 cell_1rw
* cell instance $13759 m0 *1 96.585,73.71
X$13759 340 54 341 644 645 cell_1rw
* cell instance $13760 m0 *1 97.29,73.71
X$13760 342 54 343 644 645 cell_1rw
* cell instance $13761 m0 *1 97.995,73.71
X$13761 344 54 345 644 645 cell_1rw
* cell instance $13762 m0 *1 98.7,73.71
X$13762 346 54 347 644 645 cell_1rw
* cell instance $13763 m0 *1 99.405,73.71
X$13763 348 54 349 644 645 cell_1rw
* cell instance $13764 m0 *1 100.11,73.71
X$13764 350 54 351 644 645 cell_1rw
* cell instance $13765 m0 *1 100.815,73.71
X$13765 352 54 353 644 645 cell_1rw
* cell instance $13766 m0 *1 101.52,73.71
X$13766 354 54 355 644 645 cell_1rw
* cell instance $13767 m0 *1 102.225,73.71
X$13767 356 54 357 644 645 cell_1rw
* cell instance $13768 m0 *1 102.93,73.71
X$13768 358 54 359 644 645 cell_1rw
* cell instance $13769 m0 *1 103.635,73.71
X$13769 360 54 361 644 645 cell_1rw
* cell instance $13770 m0 *1 104.34,73.71
X$13770 362 54 363 644 645 cell_1rw
* cell instance $13771 m0 *1 105.045,73.71
X$13771 364 54 365 644 645 cell_1rw
* cell instance $13772 m0 *1 105.75,73.71
X$13772 366 54 367 644 645 cell_1rw
* cell instance $13773 m0 *1 106.455,73.71
X$13773 368 54 369 644 645 cell_1rw
* cell instance $13774 m0 *1 107.16,73.71
X$13774 370 54 371 644 645 cell_1rw
* cell instance $13775 m0 *1 107.865,73.71
X$13775 372 54 373 644 645 cell_1rw
* cell instance $13776 m0 *1 108.57,73.71
X$13776 374 54 375 644 645 cell_1rw
* cell instance $13777 m0 *1 109.275,73.71
X$13777 376 54 377 644 645 cell_1rw
* cell instance $13778 m0 *1 109.98,73.71
X$13778 378 54 379 644 645 cell_1rw
* cell instance $13779 m0 *1 110.685,73.71
X$13779 380 54 381 644 645 cell_1rw
* cell instance $13780 m0 *1 111.39,73.71
X$13780 382 54 383 644 645 cell_1rw
* cell instance $13781 m0 *1 112.095,73.71
X$13781 384 54 385 644 645 cell_1rw
* cell instance $13782 m0 *1 112.8,73.71
X$13782 386 54 387 644 645 cell_1rw
* cell instance $13783 m0 *1 113.505,73.71
X$13783 388 54 389 644 645 cell_1rw
* cell instance $13784 m0 *1 114.21,73.71
X$13784 390 54 391 644 645 cell_1rw
* cell instance $13785 m0 *1 114.915,73.71
X$13785 392 54 393 644 645 cell_1rw
* cell instance $13786 m0 *1 115.62,73.71
X$13786 394 54 395 644 645 cell_1rw
* cell instance $13787 m0 *1 116.325,73.71
X$13787 396 54 397 644 645 cell_1rw
* cell instance $13788 m0 *1 117.03,73.71
X$13788 398 54 399 644 645 cell_1rw
* cell instance $13789 m0 *1 117.735,73.71
X$13789 400 54 401 644 645 cell_1rw
* cell instance $13790 m0 *1 118.44,73.71
X$13790 402 54 403 644 645 cell_1rw
* cell instance $13791 m0 *1 119.145,73.71
X$13791 404 54 405 644 645 cell_1rw
* cell instance $13792 m0 *1 119.85,73.71
X$13792 406 54 407 644 645 cell_1rw
* cell instance $13793 m0 *1 120.555,73.71
X$13793 408 54 409 644 645 cell_1rw
* cell instance $13794 m0 *1 121.26,73.71
X$13794 410 54 411 644 645 cell_1rw
* cell instance $13795 m0 *1 121.965,73.71
X$13795 412 54 413 644 645 cell_1rw
* cell instance $13796 m0 *1 122.67,73.71
X$13796 414 54 415 644 645 cell_1rw
* cell instance $13797 m0 *1 123.375,73.71
X$13797 416 54 417 644 645 cell_1rw
* cell instance $13798 m0 *1 124.08,73.71
X$13798 418 54 419 644 645 cell_1rw
* cell instance $13799 m0 *1 124.785,73.71
X$13799 420 54 421 644 645 cell_1rw
* cell instance $13800 m0 *1 125.49,73.71
X$13800 422 54 423 644 645 cell_1rw
* cell instance $13801 m0 *1 126.195,73.71
X$13801 424 54 425 644 645 cell_1rw
* cell instance $13802 m0 *1 126.9,73.71
X$13802 426 54 427 644 645 cell_1rw
* cell instance $13803 m0 *1 127.605,73.71
X$13803 428 54 429 644 645 cell_1rw
* cell instance $13804 m0 *1 128.31,73.71
X$13804 430 54 431 644 645 cell_1rw
* cell instance $13805 m0 *1 129.015,73.71
X$13805 432 54 433 644 645 cell_1rw
* cell instance $13806 m0 *1 129.72,73.71
X$13806 434 54 435 644 645 cell_1rw
* cell instance $13807 m0 *1 130.425,73.71
X$13807 436 54 437 644 645 cell_1rw
* cell instance $13808 m0 *1 131.13,73.71
X$13808 438 54 439 644 645 cell_1rw
* cell instance $13809 m0 *1 131.835,73.71
X$13809 440 54 441 644 645 cell_1rw
* cell instance $13810 m0 *1 132.54,73.71
X$13810 442 54 443 644 645 cell_1rw
* cell instance $13811 m0 *1 133.245,73.71
X$13811 444 54 445 644 645 cell_1rw
* cell instance $13812 m0 *1 133.95,73.71
X$13812 446 54 447 644 645 cell_1rw
* cell instance $13813 m0 *1 134.655,73.71
X$13813 448 54 449 644 645 cell_1rw
* cell instance $13814 m0 *1 135.36,73.71
X$13814 450 54 451 644 645 cell_1rw
* cell instance $13815 m0 *1 136.065,73.71
X$13815 452 54 453 644 645 cell_1rw
* cell instance $13816 m0 *1 136.77,73.71
X$13816 454 54 455 644 645 cell_1rw
* cell instance $13817 m0 *1 137.475,73.71
X$13817 456 54 457 644 645 cell_1rw
* cell instance $13818 m0 *1 138.18,73.71
X$13818 458 54 459 644 645 cell_1rw
* cell instance $13819 m0 *1 138.885,73.71
X$13819 460 54 461 644 645 cell_1rw
* cell instance $13820 m0 *1 139.59,73.71
X$13820 462 54 463 644 645 cell_1rw
* cell instance $13821 m0 *1 140.295,73.71
X$13821 464 54 465 644 645 cell_1rw
* cell instance $13822 m0 *1 141,73.71
X$13822 466 54 467 644 645 cell_1rw
* cell instance $13823 m0 *1 141.705,73.71
X$13823 468 54 469 644 645 cell_1rw
* cell instance $13824 m0 *1 142.41,73.71
X$13824 470 54 471 644 645 cell_1rw
* cell instance $13825 m0 *1 143.115,73.71
X$13825 472 54 473 644 645 cell_1rw
* cell instance $13826 m0 *1 143.82,73.71
X$13826 474 54 475 644 645 cell_1rw
* cell instance $13827 m0 *1 144.525,73.71
X$13827 476 54 477 644 645 cell_1rw
* cell instance $13828 m0 *1 145.23,73.71
X$13828 478 54 479 644 645 cell_1rw
* cell instance $13829 m0 *1 145.935,73.71
X$13829 480 54 481 644 645 cell_1rw
* cell instance $13830 m0 *1 146.64,73.71
X$13830 482 54 483 644 645 cell_1rw
* cell instance $13831 m0 *1 147.345,73.71
X$13831 484 54 485 644 645 cell_1rw
* cell instance $13832 m0 *1 148.05,73.71
X$13832 486 54 487 644 645 cell_1rw
* cell instance $13833 m0 *1 148.755,73.71
X$13833 488 54 489 644 645 cell_1rw
* cell instance $13834 m0 *1 149.46,73.71
X$13834 490 54 491 644 645 cell_1rw
* cell instance $13835 m0 *1 150.165,73.71
X$13835 492 54 493 644 645 cell_1rw
* cell instance $13836 m0 *1 150.87,73.71
X$13836 494 54 495 644 645 cell_1rw
* cell instance $13837 m0 *1 151.575,73.71
X$13837 496 54 497 644 645 cell_1rw
* cell instance $13838 m0 *1 152.28,73.71
X$13838 498 54 499 644 645 cell_1rw
* cell instance $13839 m0 *1 152.985,73.71
X$13839 500 54 501 644 645 cell_1rw
* cell instance $13840 m0 *1 153.69,73.71
X$13840 502 54 503 644 645 cell_1rw
* cell instance $13841 m0 *1 154.395,73.71
X$13841 504 54 505 644 645 cell_1rw
* cell instance $13842 m0 *1 155.1,73.71
X$13842 506 54 507 644 645 cell_1rw
* cell instance $13843 m0 *1 155.805,73.71
X$13843 508 54 509 644 645 cell_1rw
* cell instance $13844 m0 *1 156.51,73.71
X$13844 510 54 511 644 645 cell_1rw
* cell instance $13845 m0 *1 157.215,73.71
X$13845 512 54 513 644 645 cell_1rw
* cell instance $13846 m0 *1 157.92,73.71
X$13846 514 54 515 644 645 cell_1rw
* cell instance $13847 m0 *1 158.625,73.71
X$13847 516 54 517 644 645 cell_1rw
* cell instance $13848 m0 *1 159.33,73.71
X$13848 518 54 519 644 645 cell_1rw
* cell instance $13849 m0 *1 160.035,73.71
X$13849 520 54 521 644 645 cell_1rw
* cell instance $13850 m0 *1 160.74,73.71
X$13850 522 54 523 644 645 cell_1rw
* cell instance $13851 m0 *1 161.445,73.71
X$13851 524 54 525 644 645 cell_1rw
* cell instance $13852 m0 *1 162.15,73.71
X$13852 526 54 527 644 645 cell_1rw
* cell instance $13853 m0 *1 162.855,73.71
X$13853 528 54 529 644 645 cell_1rw
* cell instance $13854 m0 *1 163.56,73.71
X$13854 530 54 531 644 645 cell_1rw
* cell instance $13855 m0 *1 164.265,73.71
X$13855 532 54 533 644 645 cell_1rw
* cell instance $13856 m0 *1 164.97,73.71
X$13856 534 54 535 644 645 cell_1rw
* cell instance $13857 m0 *1 165.675,73.71
X$13857 536 54 537 644 645 cell_1rw
* cell instance $13858 m0 *1 166.38,73.71
X$13858 538 54 539 644 645 cell_1rw
* cell instance $13859 m0 *1 167.085,73.71
X$13859 540 54 541 644 645 cell_1rw
* cell instance $13860 m0 *1 167.79,73.71
X$13860 542 54 543 644 645 cell_1rw
* cell instance $13861 m0 *1 168.495,73.71
X$13861 544 54 545 644 645 cell_1rw
* cell instance $13862 m0 *1 169.2,73.71
X$13862 546 54 547 644 645 cell_1rw
* cell instance $13863 m0 *1 169.905,73.71
X$13863 548 54 549 644 645 cell_1rw
* cell instance $13864 m0 *1 170.61,73.71
X$13864 550 54 551 644 645 cell_1rw
* cell instance $13865 m0 *1 171.315,73.71
X$13865 552 54 553 644 645 cell_1rw
* cell instance $13866 m0 *1 172.02,73.71
X$13866 554 54 555 644 645 cell_1rw
* cell instance $13867 m0 *1 172.725,73.71
X$13867 556 54 557 644 645 cell_1rw
* cell instance $13868 m0 *1 173.43,73.71
X$13868 558 54 559 644 645 cell_1rw
* cell instance $13869 m0 *1 174.135,73.71
X$13869 560 54 561 644 645 cell_1rw
* cell instance $13870 m0 *1 174.84,73.71
X$13870 562 54 563 644 645 cell_1rw
* cell instance $13871 m0 *1 175.545,73.71
X$13871 564 54 565 644 645 cell_1rw
* cell instance $13872 m0 *1 176.25,73.71
X$13872 566 54 567 644 645 cell_1rw
* cell instance $13873 m0 *1 176.955,73.71
X$13873 568 54 569 644 645 cell_1rw
* cell instance $13874 m0 *1 177.66,73.71
X$13874 570 54 571 644 645 cell_1rw
* cell instance $13875 m0 *1 178.365,73.71
X$13875 572 54 573 644 645 cell_1rw
* cell instance $13876 m0 *1 179.07,73.71
X$13876 574 54 575 644 645 cell_1rw
* cell instance $13877 m0 *1 179.775,73.71
X$13877 576 54 577 644 645 cell_1rw
* cell instance $13878 m0 *1 180.48,73.71
X$13878 578 54 579 644 645 cell_1rw
* cell instance $13879 r0 *1 0.705,73.71
X$13879 67 55 68 644 645 cell_1rw
* cell instance $13880 r0 *1 0,73.71
X$13880 65 55 66 644 645 cell_1rw
* cell instance $13881 r0 *1 1.41,73.71
X$13881 69 55 70 644 645 cell_1rw
* cell instance $13882 r0 *1 2.115,73.71
X$13882 71 55 72 644 645 cell_1rw
* cell instance $13883 r0 *1 2.82,73.71
X$13883 73 55 74 644 645 cell_1rw
* cell instance $13884 r0 *1 3.525,73.71
X$13884 75 55 76 644 645 cell_1rw
* cell instance $13885 r0 *1 4.23,73.71
X$13885 77 55 78 644 645 cell_1rw
* cell instance $13886 r0 *1 4.935,73.71
X$13886 79 55 80 644 645 cell_1rw
* cell instance $13887 r0 *1 5.64,73.71
X$13887 81 55 82 644 645 cell_1rw
* cell instance $13888 r0 *1 6.345,73.71
X$13888 83 55 84 644 645 cell_1rw
* cell instance $13889 r0 *1 7.05,73.71
X$13889 85 55 86 644 645 cell_1rw
* cell instance $13890 r0 *1 7.755,73.71
X$13890 87 55 88 644 645 cell_1rw
* cell instance $13891 r0 *1 8.46,73.71
X$13891 89 55 90 644 645 cell_1rw
* cell instance $13892 r0 *1 9.165,73.71
X$13892 91 55 92 644 645 cell_1rw
* cell instance $13893 r0 *1 9.87,73.71
X$13893 93 55 94 644 645 cell_1rw
* cell instance $13894 r0 *1 10.575,73.71
X$13894 95 55 96 644 645 cell_1rw
* cell instance $13895 r0 *1 11.28,73.71
X$13895 97 55 98 644 645 cell_1rw
* cell instance $13896 r0 *1 11.985,73.71
X$13896 99 55 100 644 645 cell_1rw
* cell instance $13897 r0 *1 12.69,73.71
X$13897 101 55 102 644 645 cell_1rw
* cell instance $13898 r0 *1 13.395,73.71
X$13898 103 55 104 644 645 cell_1rw
* cell instance $13899 r0 *1 14.1,73.71
X$13899 105 55 106 644 645 cell_1rw
* cell instance $13900 r0 *1 14.805,73.71
X$13900 107 55 108 644 645 cell_1rw
* cell instance $13901 r0 *1 15.51,73.71
X$13901 109 55 110 644 645 cell_1rw
* cell instance $13902 r0 *1 16.215,73.71
X$13902 111 55 112 644 645 cell_1rw
* cell instance $13903 r0 *1 16.92,73.71
X$13903 113 55 114 644 645 cell_1rw
* cell instance $13904 r0 *1 17.625,73.71
X$13904 115 55 116 644 645 cell_1rw
* cell instance $13905 r0 *1 18.33,73.71
X$13905 117 55 118 644 645 cell_1rw
* cell instance $13906 r0 *1 19.035,73.71
X$13906 119 55 120 644 645 cell_1rw
* cell instance $13907 r0 *1 19.74,73.71
X$13907 121 55 122 644 645 cell_1rw
* cell instance $13908 r0 *1 20.445,73.71
X$13908 123 55 124 644 645 cell_1rw
* cell instance $13909 r0 *1 21.15,73.71
X$13909 125 55 126 644 645 cell_1rw
* cell instance $13910 r0 *1 21.855,73.71
X$13910 127 55 128 644 645 cell_1rw
* cell instance $13911 r0 *1 22.56,73.71
X$13911 129 55 130 644 645 cell_1rw
* cell instance $13912 r0 *1 23.265,73.71
X$13912 131 55 132 644 645 cell_1rw
* cell instance $13913 r0 *1 23.97,73.71
X$13913 133 55 134 644 645 cell_1rw
* cell instance $13914 r0 *1 24.675,73.71
X$13914 135 55 136 644 645 cell_1rw
* cell instance $13915 r0 *1 25.38,73.71
X$13915 137 55 138 644 645 cell_1rw
* cell instance $13916 r0 *1 26.085,73.71
X$13916 139 55 140 644 645 cell_1rw
* cell instance $13917 r0 *1 26.79,73.71
X$13917 141 55 142 644 645 cell_1rw
* cell instance $13918 r0 *1 27.495,73.71
X$13918 143 55 144 644 645 cell_1rw
* cell instance $13919 r0 *1 28.2,73.71
X$13919 145 55 146 644 645 cell_1rw
* cell instance $13920 r0 *1 28.905,73.71
X$13920 147 55 148 644 645 cell_1rw
* cell instance $13921 r0 *1 29.61,73.71
X$13921 149 55 150 644 645 cell_1rw
* cell instance $13922 r0 *1 30.315,73.71
X$13922 151 55 152 644 645 cell_1rw
* cell instance $13923 r0 *1 31.02,73.71
X$13923 153 55 154 644 645 cell_1rw
* cell instance $13924 r0 *1 31.725,73.71
X$13924 155 55 156 644 645 cell_1rw
* cell instance $13925 r0 *1 32.43,73.71
X$13925 157 55 158 644 645 cell_1rw
* cell instance $13926 r0 *1 33.135,73.71
X$13926 159 55 160 644 645 cell_1rw
* cell instance $13927 r0 *1 33.84,73.71
X$13927 161 55 162 644 645 cell_1rw
* cell instance $13928 r0 *1 34.545,73.71
X$13928 163 55 164 644 645 cell_1rw
* cell instance $13929 r0 *1 35.25,73.71
X$13929 165 55 166 644 645 cell_1rw
* cell instance $13930 r0 *1 35.955,73.71
X$13930 167 55 168 644 645 cell_1rw
* cell instance $13931 r0 *1 36.66,73.71
X$13931 169 55 170 644 645 cell_1rw
* cell instance $13932 r0 *1 37.365,73.71
X$13932 171 55 172 644 645 cell_1rw
* cell instance $13933 r0 *1 38.07,73.71
X$13933 173 55 174 644 645 cell_1rw
* cell instance $13934 r0 *1 38.775,73.71
X$13934 175 55 176 644 645 cell_1rw
* cell instance $13935 r0 *1 39.48,73.71
X$13935 177 55 178 644 645 cell_1rw
* cell instance $13936 r0 *1 40.185,73.71
X$13936 179 55 180 644 645 cell_1rw
* cell instance $13937 r0 *1 40.89,73.71
X$13937 181 55 182 644 645 cell_1rw
* cell instance $13938 r0 *1 41.595,73.71
X$13938 183 55 184 644 645 cell_1rw
* cell instance $13939 r0 *1 42.3,73.71
X$13939 185 55 186 644 645 cell_1rw
* cell instance $13940 r0 *1 43.005,73.71
X$13940 187 55 188 644 645 cell_1rw
* cell instance $13941 r0 *1 43.71,73.71
X$13941 189 55 190 644 645 cell_1rw
* cell instance $13942 r0 *1 44.415,73.71
X$13942 191 55 192 644 645 cell_1rw
* cell instance $13943 r0 *1 45.12,73.71
X$13943 193 55 194 644 645 cell_1rw
* cell instance $13944 r0 *1 45.825,73.71
X$13944 195 55 196 644 645 cell_1rw
* cell instance $13945 r0 *1 46.53,73.71
X$13945 197 55 198 644 645 cell_1rw
* cell instance $13946 r0 *1 47.235,73.71
X$13946 199 55 200 644 645 cell_1rw
* cell instance $13947 r0 *1 47.94,73.71
X$13947 201 55 202 644 645 cell_1rw
* cell instance $13948 r0 *1 48.645,73.71
X$13948 203 55 204 644 645 cell_1rw
* cell instance $13949 r0 *1 49.35,73.71
X$13949 205 55 206 644 645 cell_1rw
* cell instance $13950 r0 *1 50.055,73.71
X$13950 207 55 208 644 645 cell_1rw
* cell instance $13951 r0 *1 50.76,73.71
X$13951 209 55 210 644 645 cell_1rw
* cell instance $13952 r0 *1 51.465,73.71
X$13952 211 55 212 644 645 cell_1rw
* cell instance $13953 r0 *1 52.17,73.71
X$13953 213 55 214 644 645 cell_1rw
* cell instance $13954 r0 *1 52.875,73.71
X$13954 215 55 216 644 645 cell_1rw
* cell instance $13955 r0 *1 53.58,73.71
X$13955 217 55 218 644 645 cell_1rw
* cell instance $13956 r0 *1 54.285,73.71
X$13956 219 55 220 644 645 cell_1rw
* cell instance $13957 r0 *1 54.99,73.71
X$13957 221 55 222 644 645 cell_1rw
* cell instance $13958 r0 *1 55.695,73.71
X$13958 223 55 224 644 645 cell_1rw
* cell instance $13959 r0 *1 56.4,73.71
X$13959 225 55 226 644 645 cell_1rw
* cell instance $13960 r0 *1 57.105,73.71
X$13960 227 55 228 644 645 cell_1rw
* cell instance $13961 r0 *1 57.81,73.71
X$13961 229 55 230 644 645 cell_1rw
* cell instance $13962 r0 *1 58.515,73.71
X$13962 231 55 232 644 645 cell_1rw
* cell instance $13963 r0 *1 59.22,73.71
X$13963 233 55 234 644 645 cell_1rw
* cell instance $13964 r0 *1 59.925,73.71
X$13964 235 55 236 644 645 cell_1rw
* cell instance $13965 r0 *1 60.63,73.71
X$13965 237 55 238 644 645 cell_1rw
* cell instance $13966 r0 *1 61.335,73.71
X$13966 239 55 240 644 645 cell_1rw
* cell instance $13967 r0 *1 62.04,73.71
X$13967 241 55 242 644 645 cell_1rw
* cell instance $13968 r0 *1 62.745,73.71
X$13968 243 55 244 644 645 cell_1rw
* cell instance $13969 r0 *1 63.45,73.71
X$13969 245 55 246 644 645 cell_1rw
* cell instance $13970 r0 *1 64.155,73.71
X$13970 247 55 248 644 645 cell_1rw
* cell instance $13971 r0 *1 64.86,73.71
X$13971 249 55 250 644 645 cell_1rw
* cell instance $13972 r0 *1 65.565,73.71
X$13972 251 55 252 644 645 cell_1rw
* cell instance $13973 r0 *1 66.27,73.71
X$13973 253 55 254 644 645 cell_1rw
* cell instance $13974 r0 *1 66.975,73.71
X$13974 255 55 256 644 645 cell_1rw
* cell instance $13975 r0 *1 67.68,73.71
X$13975 257 55 258 644 645 cell_1rw
* cell instance $13976 r0 *1 68.385,73.71
X$13976 259 55 260 644 645 cell_1rw
* cell instance $13977 r0 *1 69.09,73.71
X$13977 261 55 262 644 645 cell_1rw
* cell instance $13978 r0 *1 69.795,73.71
X$13978 263 55 264 644 645 cell_1rw
* cell instance $13979 r0 *1 70.5,73.71
X$13979 265 55 266 644 645 cell_1rw
* cell instance $13980 r0 *1 71.205,73.71
X$13980 267 55 268 644 645 cell_1rw
* cell instance $13981 r0 *1 71.91,73.71
X$13981 269 55 270 644 645 cell_1rw
* cell instance $13982 r0 *1 72.615,73.71
X$13982 271 55 272 644 645 cell_1rw
* cell instance $13983 r0 *1 73.32,73.71
X$13983 273 55 274 644 645 cell_1rw
* cell instance $13984 r0 *1 74.025,73.71
X$13984 275 55 276 644 645 cell_1rw
* cell instance $13985 r0 *1 74.73,73.71
X$13985 277 55 278 644 645 cell_1rw
* cell instance $13986 r0 *1 75.435,73.71
X$13986 279 55 280 644 645 cell_1rw
* cell instance $13987 r0 *1 76.14,73.71
X$13987 281 55 282 644 645 cell_1rw
* cell instance $13988 r0 *1 76.845,73.71
X$13988 283 55 284 644 645 cell_1rw
* cell instance $13989 r0 *1 77.55,73.71
X$13989 285 55 286 644 645 cell_1rw
* cell instance $13990 r0 *1 78.255,73.71
X$13990 287 55 288 644 645 cell_1rw
* cell instance $13991 r0 *1 78.96,73.71
X$13991 289 55 290 644 645 cell_1rw
* cell instance $13992 r0 *1 79.665,73.71
X$13992 291 55 292 644 645 cell_1rw
* cell instance $13993 r0 *1 80.37,73.71
X$13993 293 55 294 644 645 cell_1rw
* cell instance $13994 r0 *1 81.075,73.71
X$13994 295 55 296 644 645 cell_1rw
* cell instance $13995 r0 *1 81.78,73.71
X$13995 297 55 298 644 645 cell_1rw
* cell instance $13996 r0 *1 82.485,73.71
X$13996 299 55 300 644 645 cell_1rw
* cell instance $13997 r0 *1 83.19,73.71
X$13997 301 55 302 644 645 cell_1rw
* cell instance $13998 r0 *1 83.895,73.71
X$13998 303 55 304 644 645 cell_1rw
* cell instance $13999 r0 *1 84.6,73.71
X$13999 305 55 306 644 645 cell_1rw
* cell instance $14000 r0 *1 85.305,73.71
X$14000 307 55 308 644 645 cell_1rw
* cell instance $14001 r0 *1 86.01,73.71
X$14001 309 55 310 644 645 cell_1rw
* cell instance $14002 r0 *1 86.715,73.71
X$14002 311 55 312 644 645 cell_1rw
* cell instance $14003 r0 *1 87.42,73.71
X$14003 313 55 314 644 645 cell_1rw
* cell instance $14004 r0 *1 88.125,73.71
X$14004 315 55 316 644 645 cell_1rw
* cell instance $14005 r0 *1 88.83,73.71
X$14005 317 55 318 644 645 cell_1rw
* cell instance $14006 r0 *1 89.535,73.71
X$14006 319 55 320 644 645 cell_1rw
* cell instance $14007 r0 *1 90.24,73.71
X$14007 321 55 323 644 645 cell_1rw
* cell instance $14008 r0 *1 90.945,73.71
X$14008 324 55 325 644 645 cell_1rw
* cell instance $14009 r0 *1 91.65,73.71
X$14009 326 55 327 644 645 cell_1rw
* cell instance $14010 r0 *1 92.355,73.71
X$14010 328 55 329 644 645 cell_1rw
* cell instance $14011 r0 *1 93.06,73.71
X$14011 330 55 331 644 645 cell_1rw
* cell instance $14012 r0 *1 93.765,73.71
X$14012 332 55 333 644 645 cell_1rw
* cell instance $14013 r0 *1 94.47,73.71
X$14013 334 55 335 644 645 cell_1rw
* cell instance $14014 r0 *1 95.175,73.71
X$14014 336 55 337 644 645 cell_1rw
* cell instance $14015 r0 *1 95.88,73.71
X$14015 338 55 339 644 645 cell_1rw
* cell instance $14016 r0 *1 96.585,73.71
X$14016 340 55 341 644 645 cell_1rw
* cell instance $14017 r0 *1 97.29,73.71
X$14017 342 55 343 644 645 cell_1rw
* cell instance $14018 r0 *1 97.995,73.71
X$14018 344 55 345 644 645 cell_1rw
* cell instance $14019 r0 *1 98.7,73.71
X$14019 346 55 347 644 645 cell_1rw
* cell instance $14020 r0 *1 99.405,73.71
X$14020 348 55 349 644 645 cell_1rw
* cell instance $14021 r0 *1 100.11,73.71
X$14021 350 55 351 644 645 cell_1rw
* cell instance $14022 r0 *1 100.815,73.71
X$14022 352 55 353 644 645 cell_1rw
* cell instance $14023 r0 *1 101.52,73.71
X$14023 354 55 355 644 645 cell_1rw
* cell instance $14024 r0 *1 102.225,73.71
X$14024 356 55 357 644 645 cell_1rw
* cell instance $14025 r0 *1 102.93,73.71
X$14025 358 55 359 644 645 cell_1rw
* cell instance $14026 r0 *1 103.635,73.71
X$14026 360 55 361 644 645 cell_1rw
* cell instance $14027 r0 *1 104.34,73.71
X$14027 362 55 363 644 645 cell_1rw
* cell instance $14028 r0 *1 105.045,73.71
X$14028 364 55 365 644 645 cell_1rw
* cell instance $14029 r0 *1 105.75,73.71
X$14029 366 55 367 644 645 cell_1rw
* cell instance $14030 r0 *1 106.455,73.71
X$14030 368 55 369 644 645 cell_1rw
* cell instance $14031 r0 *1 107.16,73.71
X$14031 370 55 371 644 645 cell_1rw
* cell instance $14032 r0 *1 107.865,73.71
X$14032 372 55 373 644 645 cell_1rw
* cell instance $14033 r0 *1 108.57,73.71
X$14033 374 55 375 644 645 cell_1rw
* cell instance $14034 r0 *1 109.275,73.71
X$14034 376 55 377 644 645 cell_1rw
* cell instance $14035 r0 *1 109.98,73.71
X$14035 378 55 379 644 645 cell_1rw
* cell instance $14036 r0 *1 110.685,73.71
X$14036 380 55 381 644 645 cell_1rw
* cell instance $14037 r0 *1 111.39,73.71
X$14037 382 55 383 644 645 cell_1rw
* cell instance $14038 r0 *1 112.095,73.71
X$14038 384 55 385 644 645 cell_1rw
* cell instance $14039 r0 *1 112.8,73.71
X$14039 386 55 387 644 645 cell_1rw
* cell instance $14040 r0 *1 113.505,73.71
X$14040 388 55 389 644 645 cell_1rw
* cell instance $14041 r0 *1 114.21,73.71
X$14041 390 55 391 644 645 cell_1rw
* cell instance $14042 r0 *1 114.915,73.71
X$14042 392 55 393 644 645 cell_1rw
* cell instance $14043 r0 *1 115.62,73.71
X$14043 394 55 395 644 645 cell_1rw
* cell instance $14044 r0 *1 116.325,73.71
X$14044 396 55 397 644 645 cell_1rw
* cell instance $14045 r0 *1 117.03,73.71
X$14045 398 55 399 644 645 cell_1rw
* cell instance $14046 r0 *1 117.735,73.71
X$14046 400 55 401 644 645 cell_1rw
* cell instance $14047 r0 *1 118.44,73.71
X$14047 402 55 403 644 645 cell_1rw
* cell instance $14048 r0 *1 119.145,73.71
X$14048 404 55 405 644 645 cell_1rw
* cell instance $14049 r0 *1 119.85,73.71
X$14049 406 55 407 644 645 cell_1rw
* cell instance $14050 r0 *1 120.555,73.71
X$14050 408 55 409 644 645 cell_1rw
* cell instance $14051 r0 *1 121.26,73.71
X$14051 410 55 411 644 645 cell_1rw
* cell instance $14052 r0 *1 121.965,73.71
X$14052 412 55 413 644 645 cell_1rw
* cell instance $14053 r0 *1 122.67,73.71
X$14053 414 55 415 644 645 cell_1rw
* cell instance $14054 r0 *1 123.375,73.71
X$14054 416 55 417 644 645 cell_1rw
* cell instance $14055 r0 *1 124.08,73.71
X$14055 418 55 419 644 645 cell_1rw
* cell instance $14056 r0 *1 124.785,73.71
X$14056 420 55 421 644 645 cell_1rw
* cell instance $14057 r0 *1 125.49,73.71
X$14057 422 55 423 644 645 cell_1rw
* cell instance $14058 r0 *1 126.195,73.71
X$14058 424 55 425 644 645 cell_1rw
* cell instance $14059 r0 *1 126.9,73.71
X$14059 426 55 427 644 645 cell_1rw
* cell instance $14060 r0 *1 127.605,73.71
X$14060 428 55 429 644 645 cell_1rw
* cell instance $14061 r0 *1 128.31,73.71
X$14061 430 55 431 644 645 cell_1rw
* cell instance $14062 r0 *1 129.015,73.71
X$14062 432 55 433 644 645 cell_1rw
* cell instance $14063 r0 *1 129.72,73.71
X$14063 434 55 435 644 645 cell_1rw
* cell instance $14064 r0 *1 130.425,73.71
X$14064 436 55 437 644 645 cell_1rw
* cell instance $14065 r0 *1 131.13,73.71
X$14065 438 55 439 644 645 cell_1rw
* cell instance $14066 r0 *1 131.835,73.71
X$14066 440 55 441 644 645 cell_1rw
* cell instance $14067 r0 *1 132.54,73.71
X$14067 442 55 443 644 645 cell_1rw
* cell instance $14068 r0 *1 133.245,73.71
X$14068 444 55 445 644 645 cell_1rw
* cell instance $14069 r0 *1 133.95,73.71
X$14069 446 55 447 644 645 cell_1rw
* cell instance $14070 r0 *1 134.655,73.71
X$14070 448 55 449 644 645 cell_1rw
* cell instance $14071 r0 *1 135.36,73.71
X$14071 450 55 451 644 645 cell_1rw
* cell instance $14072 r0 *1 136.065,73.71
X$14072 452 55 453 644 645 cell_1rw
* cell instance $14073 r0 *1 136.77,73.71
X$14073 454 55 455 644 645 cell_1rw
* cell instance $14074 r0 *1 137.475,73.71
X$14074 456 55 457 644 645 cell_1rw
* cell instance $14075 r0 *1 138.18,73.71
X$14075 458 55 459 644 645 cell_1rw
* cell instance $14076 r0 *1 138.885,73.71
X$14076 460 55 461 644 645 cell_1rw
* cell instance $14077 r0 *1 139.59,73.71
X$14077 462 55 463 644 645 cell_1rw
* cell instance $14078 r0 *1 140.295,73.71
X$14078 464 55 465 644 645 cell_1rw
* cell instance $14079 r0 *1 141,73.71
X$14079 466 55 467 644 645 cell_1rw
* cell instance $14080 r0 *1 141.705,73.71
X$14080 468 55 469 644 645 cell_1rw
* cell instance $14081 r0 *1 142.41,73.71
X$14081 470 55 471 644 645 cell_1rw
* cell instance $14082 r0 *1 143.115,73.71
X$14082 472 55 473 644 645 cell_1rw
* cell instance $14083 r0 *1 143.82,73.71
X$14083 474 55 475 644 645 cell_1rw
* cell instance $14084 r0 *1 144.525,73.71
X$14084 476 55 477 644 645 cell_1rw
* cell instance $14085 r0 *1 145.23,73.71
X$14085 478 55 479 644 645 cell_1rw
* cell instance $14086 r0 *1 145.935,73.71
X$14086 480 55 481 644 645 cell_1rw
* cell instance $14087 r0 *1 146.64,73.71
X$14087 482 55 483 644 645 cell_1rw
* cell instance $14088 r0 *1 147.345,73.71
X$14088 484 55 485 644 645 cell_1rw
* cell instance $14089 r0 *1 148.05,73.71
X$14089 486 55 487 644 645 cell_1rw
* cell instance $14090 r0 *1 148.755,73.71
X$14090 488 55 489 644 645 cell_1rw
* cell instance $14091 r0 *1 149.46,73.71
X$14091 490 55 491 644 645 cell_1rw
* cell instance $14092 r0 *1 150.165,73.71
X$14092 492 55 493 644 645 cell_1rw
* cell instance $14093 r0 *1 150.87,73.71
X$14093 494 55 495 644 645 cell_1rw
* cell instance $14094 r0 *1 151.575,73.71
X$14094 496 55 497 644 645 cell_1rw
* cell instance $14095 r0 *1 152.28,73.71
X$14095 498 55 499 644 645 cell_1rw
* cell instance $14096 r0 *1 152.985,73.71
X$14096 500 55 501 644 645 cell_1rw
* cell instance $14097 r0 *1 153.69,73.71
X$14097 502 55 503 644 645 cell_1rw
* cell instance $14098 r0 *1 154.395,73.71
X$14098 504 55 505 644 645 cell_1rw
* cell instance $14099 r0 *1 155.1,73.71
X$14099 506 55 507 644 645 cell_1rw
* cell instance $14100 r0 *1 155.805,73.71
X$14100 508 55 509 644 645 cell_1rw
* cell instance $14101 r0 *1 156.51,73.71
X$14101 510 55 511 644 645 cell_1rw
* cell instance $14102 r0 *1 157.215,73.71
X$14102 512 55 513 644 645 cell_1rw
* cell instance $14103 r0 *1 157.92,73.71
X$14103 514 55 515 644 645 cell_1rw
* cell instance $14104 r0 *1 158.625,73.71
X$14104 516 55 517 644 645 cell_1rw
* cell instance $14105 r0 *1 159.33,73.71
X$14105 518 55 519 644 645 cell_1rw
* cell instance $14106 r0 *1 160.035,73.71
X$14106 520 55 521 644 645 cell_1rw
* cell instance $14107 r0 *1 160.74,73.71
X$14107 522 55 523 644 645 cell_1rw
* cell instance $14108 r0 *1 161.445,73.71
X$14108 524 55 525 644 645 cell_1rw
* cell instance $14109 r0 *1 162.15,73.71
X$14109 526 55 527 644 645 cell_1rw
* cell instance $14110 r0 *1 162.855,73.71
X$14110 528 55 529 644 645 cell_1rw
* cell instance $14111 r0 *1 163.56,73.71
X$14111 530 55 531 644 645 cell_1rw
* cell instance $14112 r0 *1 164.265,73.71
X$14112 532 55 533 644 645 cell_1rw
* cell instance $14113 r0 *1 164.97,73.71
X$14113 534 55 535 644 645 cell_1rw
* cell instance $14114 r0 *1 165.675,73.71
X$14114 536 55 537 644 645 cell_1rw
* cell instance $14115 r0 *1 166.38,73.71
X$14115 538 55 539 644 645 cell_1rw
* cell instance $14116 r0 *1 167.085,73.71
X$14116 540 55 541 644 645 cell_1rw
* cell instance $14117 r0 *1 167.79,73.71
X$14117 542 55 543 644 645 cell_1rw
* cell instance $14118 r0 *1 168.495,73.71
X$14118 544 55 545 644 645 cell_1rw
* cell instance $14119 r0 *1 169.2,73.71
X$14119 546 55 547 644 645 cell_1rw
* cell instance $14120 r0 *1 169.905,73.71
X$14120 548 55 549 644 645 cell_1rw
* cell instance $14121 r0 *1 170.61,73.71
X$14121 550 55 551 644 645 cell_1rw
* cell instance $14122 r0 *1 171.315,73.71
X$14122 552 55 553 644 645 cell_1rw
* cell instance $14123 r0 *1 172.02,73.71
X$14123 554 55 555 644 645 cell_1rw
* cell instance $14124 r0 *1 172.725,73.71
X$14124 556 55 557 644 645 cell_1rw
* cell instance $14125 r0 *1 173.43,73.71
X$14125 558 55 559 644 645 cell_1rw
* cell instance $14126 r0 *1 174.135,73.71
X$14126 560 55 561 644 645 cell_1rw
* cell instance $14127 r0 *1 174.84,73.71
X$14127 562 55 563 644 645 cell_1rw
* cell instance $14128 r0 *1 175.545,73.71
X$14128 564 55 565 644 645 cell_1rw
* cell instance $14129 r0 *1 176.25,73.71
X$14129 566 55 567 644 645 cell_1rw
* cell instance $14130 r0 *1 176.955,73.71
X$14130 568 55 569 644 645 cell_1rw
* cell instance $14131 r0 *1 177.66,73.71
X$14131 570 55 571 644 645 cell_1rw
* cell instance $14132 r0 *1 178.365,73.71
X$14132 572 55 573 644 645 cell_1rw
* cell instance $14133 r0 *1 179.07,73.71
X$14133 574 55 575 644 645 cell_1rw
* cell instance $14134 r0 *1 179.775,73.71
X$14134 576 55 577 644 645 cell_1rw
* cell instance $14135 r0 *1 180.48,73.71
X$14135 578 55 579 644 645 cell_1rw
* cell instance $14136 m0 *1 0.705,76.44
X$14136 67 56 68 644 645 cell_1rw
* cell instance $14137 m0 *1 0,76.44
X$14137 65 56 66 644 645 cell_1rw
* cell instance $14138 m0 *1 1.41,76.44
X$14138 69 56 70 644 645 cell_1rw
* cell instance $14139 m0 *1 2.115,76.44
X$14139 71 56 72 644 645 cell_1rw
* cell instance $14140 m0 *1 2.82,76.44
X$14140 73 56 74 644 645 cell_1rw
* cell instance $14141 m0 *1 3.525,76.44
X$14141 75 56 76 644 645 cell_1rw
* cell instance $14142 m0 *1 4.23,76.44
X$14142 77 56 78 644 645 cell_1rw
* cell instance $14143 m0 *1 4.935,76.44
X$14143 79 56 80 644 645 cell_1rw
* cell instance $14144 m0 *1 5.64,76.44
X$14144 81 56 82 644 645 cell_1rw
* cell instance $14145 m0 *1 6.345,76.44
X$14145 83 56 84 644 645 cell_1rw
* cell instance $14146 m0 *1 7.05,76.44
X$14146 85 56 86 644 645 cell_1rw
* cell instance $14147 m0 *1 7.755,76.44
X$14147 87 56 88 644 645 cell_1rw
* cell instance $14148 m0 *1 8.46,76.44
X$14148 89 56 90 644 645 cell_1rw
* cell instance $14149 m0 *1 9.165,76.44
X$14149 91 56 92 644 645 cell_1rw
* cell instance $14150 m0 *1 9.87,76.44
X$14150 93 56 94 644 645 cell_1rw
* cell instance $14151 m0 *1 10.575,76.44
X$14151 95 56 96 644 645 cell_1rw
* cell instance $14152 m0 *1 11.28,76.44
X$14152 97 56 98 644 645 cell_1rw
* cell instance $14153 m0 *1 11.985,76.44
X$14153 99 56 100 644 645 cell_1rw
* cell instance $14154 m0 *1 12.69,76.44
X$14154 101 56 102 644 645 cell_1rw
* cell instance $14155 m0 *1 13.395,76.44
X$14155 103 56 104 644 645 cell_1rw
* cell instance $14156 m0 *1 14.1,76.44
X$14156 105 56 106 644 645 cell_1rw
* cell instance $14157 m0 *1 14.805,76.44
X$14157 107 56 108 644 645 cell_1rw
* cell instance $14158 m0 *1 15.51,76.44
X$14158 109 56 110 644 645 cell_1rw
* cell instance $14159 m0 *1 16.215,76.44
X$14159 111 56 112 644 645 cell_1rw
* cell instance $14160 m0 *1 16.92,76.44
X$14160 113 56 114 644 645 cell_1rw
* cell instance $14161 m0 *1 17.625,76.44
X$14161 115 56 116 644 645 cell_1rw
* cell instance $14162 m0 *1 18.33,76.44
X$14162 117 56 118 644 645 cell_1rw
* cell instance $14163 m0 *1 19.035,76.44
X$14163 119 56 120 644 645 cell_1rw
* cell instance $14164 m0 *1 19.74,76.44
X$14164 121 56 122 644 645 cell_1rw
* cell instance $14165 m0 *1 20.445,76.44
X$14165 123 56 124 644 645 cell_1rw
* cell instance $14166 m0 *1 21.15,76.44
X$14166 125 56 126 644 645 cell_1rw
* cell instance $14167 m0 *1 21.855,76.44
X$14167 127 56 128 644 645 cell_1rw
* cell instance $14168 m0 *1 22.56,76.44
X$14168 129 56 130 644 645 cell_1rw
* cell instance $14169 m0 *1 23.265,76.44
X$14169 131 56 132 644 645 cell_1rw
* cell instance $14170 m0 *1 23.97,76.44
X$14170 133 56 134 644 645 cell_1rw
* cell instance $14171 m0 *1 24.675,76.44
X$14171 135 56 136 644 645 cell_1rw
* cell instance $14172 m0 *1 25.38,76.44
X$14172 137 56 138 644 645 cell_1rw
* cell instance $14173 m0 *1 26.085,76.44
X$14173 139 56 140 644 645 cell_1rw
* cell instance $14174 m0 *1 26.79,76.44
X$14174 141 56 142 644 645 cell_1rw
* cell instance $14175 m0 *1 27.495,76.44
X$14175 143 56 144 644 645 cell_1rw
* cell instance $14176 m0 *1 28.2,76.44
X$14176 145 56 146 644 645 cell_1rw
* cell instance $14177 m0 *1 28.905,76.44
X$14177 147 56 148 644 645 cell_1rw
* cell instance $14178 m0 *1 29.61,76.44
X$14178 149 56 150 644 645 cell_1rw
* cell instance $14179 m0 *1 30.315,76.44
X$14179 151 56 152 644 645 cell_1rw
* cell instance $14180 m0 *1 31.02,76.44
X$14180 153 56 154 644 645 cell_1rw
* cell instance $14181 m0 *1 31.725,76.44
X$14181 155 56 156 644 645 cell_1rw
* cell instance $14182 m0 *1 32.43,76.44
X$14182 157 56 158 644 645 cell_1rw
* cell instance $14183 m0 *1 33.135,76.44
X$14183 159 56 160 644 645 cell_1rw
* cell instance $14184 m0 *1 33.84,76.44
X$14184 161 56 162 644 645 cell_1rw
* cell instance $14185 m0 *1 34.545,76.44
X$14185 163 56 164 644 645 cell_1rw
* cell instance $14186 m0 *1 35.25,76.44
X$14186 165 56 166 644 645 cell_1rw
* cell instance $14187 m0 *1 35.955,76.44
X$14187 167 56 168 644 645 cell_1rw
* cell instance $14188 m0 *1 36.66,76.44
X$14188 169 56 170 644 645 cell_1rw
* cell instance $14189 m0 *1 37.365,76.44
X$14189 171 56 172 644 645 cell_1rw
* cell instance $14190 m0 *1 38.07,76.44
X$14190 173 56 174 644 645 cell_1rw
* cell instance $14191 m0 *1 38.775,76.44
X$14191 175 56 176 644 645 cell_1rw
* cell instance $14192 m0 *1 39.48,76.44
X$14192 177 56 178 644 645 cell_1rw
* cell instance $14193 m0 *1 40.185,76.44
X$14193 179 56 180 644 645 cell_1rw
* cell instance $14194 m0 *1 40.89,76.44
X$14194 181 56 182 644 645 cell_1rw
* cell instance $14195 m0 *1 41.595,76.44
X$14195 183 56 184 644 645 cell_1rw
* cell instance $14196 m0 *1 42.3,76.44
X$14196 185 56 186 644 645 cell_1rw
* cell instance $14197 m0 *1 43.005,76.44
X$14197 187 56 188 644 645 cell_1rw
* cell instance $14198 m0 *1 43.71,76.44
X$14198 189 56 190 644 645 cell_1rw
* cell instance $14199 m0 *1 44.415,76.44
X$14199 191 56 192 644 645 cell_1rw
* cell instance $14200 m0 *1 45.12,76.44
X$14200 193 56 194 644 645 cell_1rw
* cell instance $14201 m0 *1 45.825,76.44
X$14201 195 56 196 644 645 cell_1rw
* cell instance $14202 m0 *1 46.53,76.44
X$14202 197 56 198 644 645 cell_1rw
* cell instance $14203 m0 *1 47.235,76.44
X$14203 199 56 200 644 645 cell_1rw
* cell instance $14204 m0 *1 47.94,76.44
X$14204 201 56 202 644 645 cell_1rw
* cell instance $14205 m0 *1 48.645,76.44
X$14205 203 56 204 644 645 cell_1rw
* cell instance $14206 m0 *1 49.35,76.44
X$14206 205 56 206 644 645 cell_1rw
* cell instance $14207 m0 *1 50.055,76.44
X$14207 207 56 208 644 645 cell_1rw
* cell instance $14208 m0 *1 50.76,76.44
X$14208 209 56 210 644 645 cell_1rw
* cell instance $14209 m0 *1 51.465,76.44
X$14209 211 56 212 644 645 cell_1rw
* cell instance $14210 m0 *1 52.17,76.44
X$14210 213 56 214 644 645 cell_1rw
* cell instance $14211 m0 *1 52.875,76.44
X$14211 215 56 216 644 645 cell_1rw
* cell instance $14212 m0 *1 53.58,76.44
X$14212 217 56 218 644 645 cell_1rw
* cell instance $14213 m0 *1 54.285,76.44
X$14213 219 56 220 644 645 cell_1rw
* cell instance $14214 m0 *1 54.99,76.44
X$14214 221 56 222 644 645 cell_1rw
* cell instance $14215 m0 *1 55.695,76.44
X$14215 223 56 224 644 645 cell_1rw
* cell instance $14216 m0 *1 56.4,76.44
X$14216 225 56 226 644 645 cell_1rw
* cell instance $14217 m0 *1 57.105,76.44
X$14217 227 56 228 644 645 cell_1rw
* cell instance $14218 m0 *1 57.81,76.44
X$14218 229 56 230 644 645 cell_1rw
* cell instance $14219 m0 *1 58.515,76.44
X$14219 231 56 232 644 645 cell_1rw
* cell instance $14220 m0 *1 59.22,76.44
X$14220 233 56 234 644 645 cell_1rw
* cell instance $14221 m0 *1 59.925,76.44
X$14221 235 56 236 644 645 cell_1rw
* cell instance $14222 m0 *1 60.63,76.44
X$14222 237 56 238 644 645 cell_1rw
* cell instance $14223 m0 *1 61.335,76.44
X$14223 239 56 240 644 645 cell_1rw
* cell instance $14224 m0 *1 62.04,76.44
X$14224 241 56 242 644 645 cell_1rw
* cell instance $14225 m0 *1 62.745,76.44
X$14225 243 56 244 644 645 cell_1rw
* cell instance $14226 m0 *1 63.45,76.44
X$14226 245 56 246 644 645 cell_1rw
* cell instance $14227 m0 *1 64.155,76.44
X$14227 247 56 248 644 645 cell_1rw
* cell instance $14228 m0 *1 64.86,76.44
X$14228 249 56 250 644 645 cell_1rw
* cell instance $14229 m0 *1 65.565,76.44
X$14229 251 56 252 644 645 cell_1rw
* cell instance $14230 m0 *1 66.27,76.44
X$14230 253 56 254 644 645 cell_1rw
* cell instance $14231 m0 *1 66.975,76.44
X$14231 255 56 256 644 645 cell_1rw
* cell instance $14232 m0 *1 67.68,76.44
X$14232 257 56 258 644 645 cell_1rw
* cell instance $14233 m0 *1 68.385,76.44
X$14233 259 56 260 644 645 cell_1rw
* cell instance $14234 m0 *1 69.09,76.44
X$14234 261 56 262 644 645 cell_1rw
* cell instance $14235 m0 *1 69.795,76.44
X$14235 263 56 264 644 645 cell_1rw
* cell instance $14236 m0 *1 70.5,76.44
X$14236 265 56 266 644 645 cell_1rw
* cell instance $14237 m0 *1 71.205,76.44
X$14237 267 56 268 644 645 cell_1rw
* cell instance $14238 m0 *1 71.91,76.44
X$14238 269 56 270 644 645 cell_1rw
* cell instance $14239 m0 *1 72.615,76.44
X$14239 271 56 272 644 645 cell_1rw
* cell instance $14240 m0 *1 73.32,76.44
X$14240 273 56 274 644 645 cell_1rw
* cell instance $14241 m0 *1 74.025,76.44
X$14241 275 56 276 644 645 cell_1rw
* cell instance $14242 m0 *1 74.73,76.44
X$14242 277 56 278 644 645 cell_1rw
* cell instance $14243 m0 *1 75.435,76.44
X$14243 279 56 280 644 645 cell_1rw
* cell instance $14244 m0 *1 76.14,76.44
X$14244 281 56 282 644 645 cell_1rw
* cell instance $14245 m0 *1 76.845,76.44
X$14245 283 56 284 644 645 cell_1rw
* cell instance $14246 m0 *1 77.55,76.44
X$14246 285 56 286 644 645 cell_1rw
* cell instance $14247 m0 *1 78.255,76.44
X$14247 287 56 288 644 645 cell_1rw
* cell instance $14248 m0 *1 78.96,76.44
X$14248 289 56 290 644 645 cell_1rw
* cell instance $14249 m0 *1 79.665,76.44
X$14249 291 56 292 644 645 cell_1rw
* cell instance $14250 m0 *1 80.37,76.44
X$14250 293 56 294 644 645 cell_1rw
* cell instance $14251 m0 *1 81.075,76.44
X$14251 295 56 296 644 645 cell_1rw
* cell instance $14252 m0 *1 81.78,76.44
X$14252 297 56 298 644 645 cell_1rw
* cell instance $14253 m0 *1 82.485,76.44
X$14253 299 56 300 644 645 cell_1rw
* cell instance $14254 m0 *1 83.19,76.44
X$14254 301 56 302 644 645 cell_1rw
* cell instance $14255 m0 *1 83.895,76.44
X$14255 303 56 304 644 645 cell_1rw
* cell instance $14256 m0 *1 84.6,76.44
X$14256 305 56 306 644 645 cell_1rw
* cell instance $14257 m0 *1 85.305,76.44
X$14257 307 56 308 644 645 cell_1rw
* cell instance $14258 m0 *1 86.01,76.44
X$14258 309 56 310 644 645 cell_1rw
* cell instance $14259 m0 *1 86.715,76.44
X$14259 311 56 312 644 645 cell_1rw
* cell instance $14260 m0 *1 87.42,76.44
X$14260 313 56 314 644 645 cell_1rw
* cell instance $14261 m0 *1 88.125,76.44
X$14261 315 56 316 644 645 cell_1rw
* cell instance $14262 m0 *1 88.83,76.44
X$14262 317 56 318 644 645 cell_1rw
* cell instance $14263 m0 *1 89.535,76.44
X$14263 319 56 320 644 645 cell_1rw
* cell instance $14264 m0 *1 90.24,76.44
X$14264 321 56 323 644 645 cell_1rw
* cell instance $14265 m0 *1 90.945,76.44
X$14265 324 56 325 644 645 cell_1rw
* cell instance $14266 m0 *1 91.65,76.44
X$14266 326 56 327 644 645 cell_1rw
* cell instance $14267 m0 *1 92.355,76.44
X$14267 328 56 329 644 645 cell_1rw
* cell instance $14268 m0 *1 93.06,76.44
X$14268 330 56 331 644 645 cell_1rw
* cell instance $14269 m0 *1 93.765,76.44
X$14269 332 56 333 644 645 cell_1rw
* cell instance $14270 m0 *1 94.47,76.44
X$14270 334 56 335 644 645 cell_1rw
* cell instance $14271 m0 *1 95.175,76.44
X$14271 336 56 337 644 645 cell_1rw
* cell instance $14272 m0 *1 95.88,76.44
X$14272 338 56 339 644 645 cell_1rw
* cell instance $14273 m0 *1 96.585,76.44
X$14273 340 56 341 644 645 cell_1rw
* cell instance $14274 m0 *1 97.29,76.44
X$14274 342 56 343 644 645 cell_1rw
* cell instance $14275 m0 *1 97.995,76.44
X$14275 344 56 345 644 645 cell_1rw
* cell instance $14276 m0 *1 98.7,76.44
X$14276 346 56 347 644 645 cell_1rw
* cell instance $14277 m0 *1 99.405,76.44
X$14277 348 56 349 644 645 cell_1rw
* cell instance $14278 m0 *1 100.11,76.44
X$14278 350 56 351 644 645 cell_1rw
* cell instance $14279 m0 *1 100.815,76.44
X$14279 352 56 353 644 645 cell_1rw
* cell instance $14280 m0 *1 101.52,76.44
X$14280 354 56 355 644 645 cell_1rw
* cell instance $14281 m0 *1 102.225,76.44
X$14281 356 56 357 644 645 cell_1rw
* cell instance $14282 m0 *1 102.93,76.44
X$14282 358 56 359 644 645 cell_1rw
* cell instance $14283 m0 *1 103.635,76.44
X$14283 360 56 361 644 645 cell_1rw
* cell instance $14284 m0 *1 104.34,76.44
X$14284 362 56 363 644 645 cell_1rw
* cell instance $14285 m0 *1 105.045,76.44
X$14285 364 56 365 644 645 cell_1rw
* cell instance $14286 m0 *1 105.75,76.44
X$14286 366 56 367 644 645 cell_1rw
* cell instance $14287 m0 *1 106.455,76.44
X$14287 368 56 369 644 645 cell_1rw
* cell instance $14288 m0 *1 107.16,76.44
X$14288 370 56 371 644 645 cell_1rw
* cell instance $14289 m0 *1 107.865,76.44
X$14289 372 56 373 644 645 cell_1rw
* cell instance $14290 m0 *1 108.57,76.44
X$14290 374 56 375 644 645 cell_1rw
* cell instance $14291 m0 *1 109.275,76.44
X$14291 376 56 377 644 645 cell_1rw
* cell instance $14292 m0 *1 109.98,76.44
X$14292 378 56 379 644 645 cell_1rw
* cell instance $14293 m0 *1 110.685,76.44
X$14293 380 56 381 644 645 cell_1rw
* cell instance $14294 m0 *1 111.39,76.44
X$14294 382 56 383 644 645 cell_1rw
* cell instance $14295 m0 *1 112.095,76.44
X$14295 384 56 385 644 645 cell_1rw
* cell instance $14296 m0 *1 112.8,76.44
X$14296 386 56 387 644 645 cell_1rw
* cell instance $14297 m0 *1 113.505,76.44
X$14297 388 56 389 644 645 cell_1rw
* cell instance $14298 m0 *1 114.21,76.44
X$14298 390 56 391 644 645 cell_1rw
* cell instance $14299 m0 *1 114.915,76.44
X$14299 392 56 393 644 645 cell_1rw
* cell instance $14300 m0 *1 115.62,76.44
X$14300 394 56 395 644 645 cell_1rw
* cell instance $14301 m0 *1 116.325,76.44
X$14301 396 56 397 644 645 cell_1rw
* cell instance $14302 m0 *1 117.03,76.44
X$14302 398 56 399 644 645 cell_1rw
* cell instance $14303 m0 *1 117.735,76.44
X$14303 400 56 401 644 645 cell_1rw
* cell instance $14304 m0 *1 118.44,76.44
X$14304 402 56 403 644 645 cell_1rw
* cell instance $14305 m0 *1 119.145,76.44
X$14305 404 56 405 644 645 cell_1rw
* cell instance $14306 m0 *1 119.85,76.44
X$14306 406 56 407 644 645 cell_1rw
* cell instance $14307 m0 *1 120.555,76.44
X$14307 408 56 409 644 645 cell_1rw
* cell instance $14308 m0 *1 121.26,76.44
X$14308 410 56 411 644 645 cell_1rw
* cell instance $14309 m0 *1 121.965,76.44
X$14309 412 56 413 644 645 cell_1rw
* cell instance $14310 m0 *1 122.67,76.44
X$14310 414 56 415 644 645 cell_1rw
* cell instance $14311 m0 *1 123.375,76.44
X$14311 416 56 417 644 645 cell_1rw
* cell instance $14312 m0 *1 124.08,76.44
X$14312 418 56 419 644 645 cell_1rw
* cell instance $14313 m0 *1 124.785,76.44
X$14313 420 56 421 644 645 cell_1rw
* cell instance $14314 m0 *1 125.49,76.44
X$14314 422 56 423 644 645 cell_1rw
* cell instance $14315 m0 *1 126.195,76.44
X$14315 424 56 425 644 645 cell_1rw
* cell instance $14316 m0 *1 126.9,76.44
X$14316 426 56 427 644 645 cell_1rw
* cell instance $14317 m0 *1 127.605,76.44
X$14317 428 56 429 644 645 cell_1rw
* cell instance $14318 m0 *1 128.31,76.44
X$14318 430 56 431 644 645 cell_1rw
* cell instance $14319 m0 *1 129.015,76.44
X$14319 432 56 433 644 645 cell_1rw
* cell instance $14320 m0 *1 129.72,76.44
X$14320 434 56 435 644 645 cell_1rw
* cell instance $14321 m0 *1 130.425,76.44
X$14321 436 56 437 644 645 cell_1rw
* cell instance $14322 m0 *1 131.13,76.44
X$14322 438 56 439 644 645 cell_1rw
* cell instance $14323 m0 *1 131.835,76.44
X$14323 440 56 441 644 645 cell_1rw
* cell instance $14324 m0 *1 132.54,76.44
X$14324 442 56 443 644 645 cell_1rw
* cell instance $14325 m0 *1 133.245,76.44
X$14325 444 56 445 644 645 cell_1rw
* cell instance $14326 m0 *1 133.95,76.44
X$14326 446 56 447 644 645 cell_1rw
* cell instance $14327 m0 *1 134.655,76.44
X$14327 448 56 449 644 645 cell_1rw
* cell instance $14328 m0 *1 135.36,76.44
X$14328 450 56 451 644 645 cell_1rw
* cell instance $14329 m0 *1 136.065,76.44
X$14329 452 56 453 644 645 cell_1rw
* cell instance $14330 m0 *1 136.77,76.44
X$14330 454 56 455 644 645 cell_1rw
* cell instance $14331 m0 *1 137.475,76.44
X$14331 456 56 457 644 645 cell_1rw
* cell instance $14332 m0 *1 138.18,76.44
X$14332 458 56 459 644 645 cell_1rw
* cell instance $14333 m0 *1 138.885,76.44
X$14333 460 56 461 644 645 cell_1rw
* cell instance $14334 m0 *1 139.59,76.44
X$14334 462 56 463 644 645 cell_1rw
* cell instance $14335 m0 *1 140.295,76.44
X$14335 464 56 465 644 645 cell_1rw
* cell instance $14336 m0 *1 141,76.44
X$14336 466 56 467 644 645 cell_1rw
* cell instance $14337 m0 *1 141.705,76.44
X$14337 468 56 469 644 645 cell_1rw
* cell instance $14338 m0 *1 142.41,76.44
X$14338 470 56 471 644 645 cell_1rw
* cell instance $14339 m0 *1 143.115,76.44
X$14339 472 56 473 644 645 cell_1rw
* cell instance $14340 m0 *1 143.82,76.44
X$14340 474 56 475 644 645 cell_1rw
* cell instance $14341 m0 *1 144.525,76.44
X$14341 476 56 477 644 645 cell_1rw
* cell instance $14342 m0 *1 145.23,76.44
X$14342 478 56 479 644 645 cell_1rw
* cell instance $14343 m0 *1 145.935,76.44
X$14343 480 56 481 644 645 cell_1rw
* cell instance $14344 m0 *1 146.64,76.44
X$14344 482 56 483 644 645 cell_1rw
* cell instance $14345 m0 *1 147.345,76.44
X$14345 484 56 485 644 645 cell_1rw
* cell instance $14346 m0 *1 148.05,76.44
X$14346 486 56 487 644 645 cell_1rw
* cell instance $14347 m0 *1 148.755,76.44
X$14347 488 56 489 644 645 cell_1rw
* cell instance $14348 m0 *1 149.46,76.44
X$14348 490 56 491 644 645 cell_1rw
* cell instance $14349 m0 *1 150.165,76.44
X$14349 492 56 493 644 645 cell_1rw
* cell instance $14350 m0 *1 150.87,76.44
X$14350 494 56 495 644 645 cell_1rw
* cell instance $14351 m0 *1 151.575,76.44
X$14351 496 56 497 644 645 cell_1rw
* cell instance $14352 m0 *1 152.28,76.44
X$14352 498 56 499 644 645 cell_1rw
* cell instance $14353 m0 *1 152.985,76.44
X$14353 500 56 501 644 645 cell_1rw
* cell instance $14354 m0 *1 153.69,76.44
X$14354 502 56 503 644 645 cell_1rw
* cell instance $14355 m0 *1 154.395,76.44
X$14355 504 56 505 644 645 cell_1rw
* cell instance $14356 m0 *1 155.1,76.44
X$14356 506 56 507 644 645 cell_1rw
* cell instance $14357 m0 *1 155.805,76.44
X$14357 508 56 509 644 645 cell_1rw
* cell instance $14358 m0 *1 156.51,76.44
X$14358 510 56 511 644 645 cell_1rw
* cell instance $14359 m0 *1 157.215,76.44
X$14359 512 56 513 644 645 cell_1rw
* cell instance $14360 m0 *1 157.92,76.44
X$14360 514 56 515 644 645 cell_1rw
* cell instance $14361 m0 *1 158.625,76.44
X$14361 516 56 517 644 645 cell_1rw
* cell instance $14362 m0 *1 159.33,76.44
X$14362 518 56 519 644 645 cell_1rw
* cell instance $14363 m0 *1 160.035,76.44
X$14363 520 56 521 644 645 cell_1rw
* cell instance $14364 m0 *1 160.74,76.44
X$14364 522 56 523 644 645 cell_1rw
* cell instance $14365 m0 *1 161.445,76.44
X$14365 524 56 525 644 645 cell_1rw
* cell instance $14366 m0 *1 162.15,76.44
X$14366 526 56 527 644 645 cell_1rw
* cell instance $14367 m0 *1 162.855,76.44
X$14367 528 56 529 644 645 cell_1rw
* cell instance $14368 m0 *1 163.56,76.44
X$14368 530 56 531 644 645 cell_1rw
* cell instance $14369 m0 *1 164.265,76.44
X$14369 532 56 533 644 645 cell_1rw
* cell instance $14370 m0 *1 164.97,76.44
X$14370 534 56 535 644 645 cell_1rw
* cell instance $14371 m0 *1 165.675,76.44
X$14371 536 56 537 644 645 cell_1rw
* cell instance $14372 m0 *1 166.38,76.44
X$14372 538 56 539 644 645 cell_1rw
* cell instance $14373 m0 *1 167.085,76.44
X$14373 540 56 541 644 645 cell_1rw
* cell instance $14374 m0 *1 167.79,76.44
X$14374 542 56 543 644 645 cell_1rw
* cell instance $14375 m0 *1 168.495,76.44
X$14375 544 56 545 644 645 cell_1rw
* cell instance $14376 m0 *1 169.2,76.44
X$14376 546 56 547 644 645 cell_1rw
* cell instance $14377 m0 *1 169.905,76.44
X$14377 548 56 549 644 645 cell_1rw
* cell instance $14378 m0 *1 170.61,76.44
X$14378 550 56 551 644 645 cell_1rw
* cell instance $14379 m0 *1 171.315,76.44
X$14379 552 56 553 644 645 cell_1rw
* cell instance $14380 m0 *1 172.02,76.44
X$14380 554 56 555 644 645 cell_1rw
* cell instance $14381 m0 *1 172.725,76.44
X$14381 556 56 557 644 645 cell_1rw
* cell instance $14382 m0 *1 173.43,76.44
X$14382 558 56 559 644 645 cell_1rw
* cell instance $14383 m0 *1 174.135,76.44
X$14383 560 56 561 644 645 cell_1rw
* cell instance $14384 m0 *1 174.84,76.44
X$14384 562 56 563 644 645 cell_1rw
* cell instance $14385 m0 *1 175.545,76.44
X$14385 564 56 565 644 645 cell_1rw
* cell instance $14386 m0 *1 176.25,76.44
X$14386 566 56 567 644 645 cell_1rw
* cell instance $14387 m0 *1 176.955,76.44
X$14387 568 56 569 644 645 cell_1rw
* cell instance $14388 m0 *1 177.66,76.44
X$14388 570 56 571 644 645 cell_1rw
* cell instance $14389 m0 *1 178.365,76.44
X$14389 572 56 573 644 645 cell_1rw
* cell instance $14390 m0 *1 179.07,76.44
X$14390 574 56 575 644 645 cell_1rw
* cell instance $14391 m0 *1 179.775,76.44
X$14391 576 56 577 644 645 cell_1rw
* cell instance $14392 m0 *1 180.48,76.44
X$14392 578 56 579 644 645 cell_1rw
* cell instance $14393 r0 *1 0.705,76.44
X$14393 67 57 68 644 645 cell_1rw
* cell instance $14394 r0 *1 0,76.44
X$14394 65 57 66 644 645 cell_1rw
* cell instance $14395 r0 *1 1.41,76.44
X$14395 69 57 70 644 645 cell_1rw
* cell instance $14396 r0 *1 2.115,76.44
X$14396 71 57 72 644 645 cell_1rw
* cell instance $14397 r0 *1 2.82,76.44
X$14397 73 57 74 644 645 cell_1rw
* cell instance $14398 r0 *1 3.525,76.44
X$14398 75 57 76 644 645 cell_1rw
* cell instance $14399 r0 *1 4.23,76.44
X$14399 77 57 78 644 645 cell_1rw
* cell instance $14400 r0 *1 4.935,76.44
X$14400 79 57 80 644 645 cell_1rw
* cell instance $14401 r0 *1 5.64,76.44
X$14401 81 57 82 644 645 cell_1rw
* cell instance $14402 r0 *1 6.345,76.44
X$14402 83 57 84 644 645 cell_1rw
* cell instance $14403 r0 *1 7.05,76.44
X$14403 85 57 86 644 645 cell_1rw
* cell instance $14404 r0 *1 7.755,76.44
X$14404 87 57 88 644 645 cell_1rw
* cell instance $14405 r0 *1 8.46,76.44
X$14405 89 57 90 644 645 cell_1rw
* cell instance $14406 r0 *1 9.165,76.44
X$14406 91 57 92 644 645 cell_1rw
* cell instance $14407 r0 *1 9.87,76.44
X$14407 93 57 94 644 645 cell_1rw
* cell instance $14408 r0 *1 10.575,76.44
X$14408 95 57 96 644 645 cell_1rw
* cell instance $14409 r0 *1 11.28,76.44
X$14409 97 57 98 644 645 cell_1rw
* cell instance $14410 r0 *1 11.985,76.44
X$14410 99 57 100 644 645 cell_1rw
* cell instance $14411 r0 *1 12.69,76.44
X$14411 101 57 102 644 645 cell_1rw
* cell instance $14412 r0 *1 13.395,76.44
X$14412 103 57 104 644 645 cell_1rw
* cell instance $14413 r0 *1 14.1,76.44
X$14413 105 57 106 644 645 cell_1rw
* cell instance $14414 r0 *1 14.805,76.44
X$14414 107 57 108 644 645 cell_1rw
* cell instance $14415 r0 *1 15.51,76.44
X$14415 109 57 110 644 645 cell_1rw
* cell instance $14416 r0 *1 16.215,76.44
X$14416 111 57 112 644 645 cell_1rw
* cell instance $14417 r0 *1 16.92,76.44
X$14417 113 57 114 644 645 cell_1rw
* cell instance $14418 r0 *1 17.625,76.44
X$14418 115 57 116 644 645 cell_1rw
* cell instance $14419 r0 *1 18.33,76.44
X$14419 117 57 118 644 645 cell_1rw
* cell instance $14420 r0 *1 19.035,76.44
X$14420 119 57 120 644 645 cell_1rw
* cell instance $14421 r0 *1 19.74,76.44
X$14421 121 57 122 644 645 cell_1rw
* cell instance $14422 r0 *1 20.445,76.44
X$14422 123 57 124 644 645 cell_1rw
* cell instance $14423 r0 *1 21.15,76.44
X$14423 125 57 126 644 645 cell_1rw
* cell instance $14424 r0 *1 21.855,76.44
X$14424 127 57 128 644 645 cell_1rw
* cell instance $14425 r0 *1 22.56,76.44
X$14425 129 57 130 644 645 cell_1rw
* cell instance $14426 r0 *1 23.265,76.44
X$14426 131 57 132 644 645 cell_1rw
* cell instance $14427 r0 *1 23.97,76.44
X$14427 133 57 134 644 645 cell_1rw
* cell instance $14428 r0 *1 24.675,76.44
X$14428 135 57 136 644 645 cell_1rw
* cell instance $14429 r0 *1 25.38,76.44
X$14429 137 57 138 644 645 cell_1rw
* cell instance $14430 r0 *1 26.085,76.44
X$14430 139 57 140 644 645 cell_1rw
* cell instance $14431 r0 *1 26.79,76.44
X$14431 141 57 142 644 645 cell_1rw
* cell instance $14432 r0 *1 27.495,76.44
X$14432 143 57 144 644 645 cell_1rw
* cell instance $14433 r0 *1 28.2,76.44
X$14433 145 57 146 644 645 cell_1rw
* cell instance $14434 r0 *1 28.905,76.44
X$14434 147 57 148 644 645 cell_1rw
* cell instance $14435 r0 *1 29.61,76.44
X$14435 149 57 150 644 645 cell_1rw
* cell instance $14436 r0 *1 30.315,76.44
X$14436 151 57 152 644 645 cell_1rw
* cell instance $14437 r0 *1 31.02,76.44
X$14437 153 57 154 644 645 cell_1rw
* cell instance $14438 r0 *1 31.725,76.44
X$14438 155 57 156 644 645 cell_1rw
* cell instance $14439 r0 *1 32.43,76.44
X$14439 157 57 158 644 645 cell_1rw
* cell instance $14440 r0 *1 33.135,76.44
X$14440 159 57 160 644 645 cell_1rw
* cell instance $14441 r0 *1 33.84,76.44
X$14441 161 57 162 644 645 cell_1rw
* cell instance $14442 r0 *1 34.545,76.44
X$14442 163 57 164 644 645 cell_1rw
* cell instance $14443 r0 *1 35.25,76.44
X$14443 165 57 166 644 645 cell_1rw
* cell instance $14444 r0 *1 35.955,76.44
X$14444 167 57 168 644 645 cell_1rw
* cell instance $14445 r0 *1 36.66,76.44
X$14445 169 57 170 644 645 cell_1rw
* cell instance $14446 r0 *1 37.365,76.44
X$14446 171 57 172 644 645 cell_1rw
* cell instance $14447 r0 *1 38.07,76.44
X$14447 173 57 174 644 645 cell_1rw
* cell instance $14448 r0 *1 38.775,76.44
X$14448 175 57 176 644 645 cell_1rw
* cell instance $14449 r0 *1 39.48,76.44
X$14449 177 57 178 644 645 cell_1rw
* cell instance $14450 r0 *1 40.185,76.44
X$14450 179 57 180 644 645 cell_1rw
* cell instance $14451 r0 *1 40.89,76.44
X$14451 181 57 182 644 645 cell_1rw
* cell instance $14452 r0 *1 41.595,76.44
X$14452 183 57 184 644 645 cell_1rw
* cell instance $14453 r0 *1 42.3,76.44
X$14453 185 57 186 644 645 cell_1rw
* cell instance $14454 r0 *1 43.005,76.44
X$14454 187 57 188 644 645 cell_1rw
* cell instance $14455 r0 *1 43.71,76.44
X$14455 189 57 190 644 645 cell_1rw
* cell instance $14456 r0 *1 44.415,76.44
X$14456 191 57 192 644 645 cell_1rw
* cell instance $14457 r0 *1 45.12,76.44
X$14457 193 57 194 644 645 cell_1rw
* cell instance $14458 r0 *1 45.825,76.44
X$14458 195 57 196 644 645 cell_1rw
* cell instance $14459 r0 *1 46.53,76.44
X$14459 197 57 198 644 645 cell_1rw
* cell instance $14460 r0 *1 47.235,76.44
X$14460 199 57 200 644 645 cell_1rw
* cell instance $14461 r0 *1 47.94,76.44
X$14461 201 57 202 644 645 cell_1rw
* cell instance $14462 r0 *1 48.645,76.44
X$14462 203 57 204 644 645 cell_1rw
* cell instance $14463 r0 *1 49.35,76.44
X$14463 205 57 206 644 645 cell_1rw
* cell instance $14464 r0 *1 50.055,76.44
X$14464 207 57 208 644 645 cell_1rw
* cell instance $14465 r0 *1 50.76,76.44
X$14465 209 57 210 644 645 cell_1rw
* cell instance $14466 r0 *1 51.465,76.44
X$14466 211 57 212 644 645 cell_1rw
* cell instance $14467 r0 *1 52.17,76.44
X$14467 213 57 214 644 645 cell_1rw
* cell instance $14468 r0 *1 52.875,76.44
X$14468 215 57 216 644 645 cell_1rw
* cell instance $14469 r0 *1 53.58,76.44
X$14469 217 57 218 644 645 cell_1rw
* cell instance $14470 r0 *1 54.285,76.44
X$14470 219 57 220 644 645 cell_1rw
* cell instance $14471 r0 *1 54.99,76.44
X$14471 221 57 222 644 645 cell_1rw
* cell instance $14472 r0 *1 55.695,76.44
X$14472 223 57 224 644 645 cell_1rw
* cell instance $14473 r0 *1 56.4,76.44
X$14473 225 57 226 644 645 cell_1rw
* cell instance $14474 r0 *1 57.105,76.44
X$14474 227 57 228 644 645 cell_1rw
* cell instance $14475 r0 *1 57.81,76.44
X$14475 229 57 230 644 645 cell_1rw
* cell instance $14476 r0 *1 58.515,76.44
X$14476 231 57 232 644 645 cell_1rw
* cell instance $14477 r0 *1 59.22,76.44
X$14477 233 57 234 644 645 cell_1rw
* cell instance $14478 r0 *1 59.925,76.44
X$14478 235 57 236 644 645 cell_1rw
* cell instance $14479 r0 *1 60.63,76.44
X$14479 237 57 238 644 645 cell_1rw
* cell instance $14480 r0 *1 61.335,76.44
X$14480 239 57 240 644 645 cell_1rw
* cell instance $14481 r0 *1 62.04,76.44
X$14481 241 57 242 644 645 cell_1rw
* cell instance $14482 r0 *1 62.745,76.44
X$14482 243 57 244 644 645 cell_1rw
* cell instance $14483 r0 *1 63.45,76.44
X$14483 245 57 246 644 645 cell_1rw
* cell instance $14484 r0 *1 64.155,76.44
X$14484 247 57 248 644 645 cell_1rw
* cell instance $14485 r0 *1 64.86,76.44
X$14485 249 57 250 644 645 cell_1rw
* cell instance $14486 r0 *1 65.565,76.44
X$14486 251 57 252 644 645 cell_1rw
* cell instance $14487 r0 *1 66.27,76.44
X$14487 253 57 254 644 645 cell_1rw
* cell instance $14488 r0 *1 66.975,76.44
X$14488 255 57 256 644 645 cell_1rw
* cell instance $14489 r0 *1 67.68,76.44
X$14489 257 57 258 644 645 cell_1rw
* cell instance $14490 r0 *1 68.385,76.44
X$14490 259 57 260 644 645 cell_1rw
* cell instance $14491 r0 *1 69.09,76.44
X$14491 261 57 262 644 645 cell_1rw
* cell instance $14492 r0 *1 69.795,76.44
X$14492 263 57 264 644 645 cell_1rw
* cell instance $14493 r0 *1 70.5,76.44
X$14493 265 57 266 644 645 cell_1rw
* cell instance $14494 r0 *1 71.205,76.44
X$14494 267 57 268 644 645 cell_1rw
* cell instance $14495 r0 *1 71.91,76.44
X$14495 269 57 270 644 645 cell_1rw
* cell instance $14496 r0 *1 72.615,76.44
X$14496 271 57 272 644 645 cell_1rw
* cell instance $14497 r0 *1 73.32,76.44
X$14497 273 57 274 644 645 cell_1rw
* cell instance $14498 r0 *1 74.025,76.44
X$14498 275 57 276 644 645 cell_1rw
* cell instance $14499 r0 *1 74.73,76.44
X$14499 277 57 278 644 645 cell_1rw
* cell instance $14500 r0 *1 75.435,76.44
X$14500 279 57 280 644 645 cell_1rw
* cell instance $14501 r0 *1 76.14,76.44
X$14501 281 57 282 644 645 cell_1rw
* cell instance $14502 r0 *1 76.845,76.44
X$14502 283 57 284 644 645 cell_1rw
* cell instance $14503 r0 *1 77.55,76.44
X$14503 285 57 286 644 645 cell_1rw
* cell instance $14504 r0 *1 78.255,76.44
X$14504 287 57 288 644 645 cell_1rw
* cell instance $14505 r0 *1 78.96,76.44
X$14505 289 57 290 644 645 cell_1rw
* cell instance $14506 r0 *1 79.665,76.44
X$14506 291 57 292 644 645 cell_1rw
* cell instance $14507 r0 *1 80.37,76.44
X$14507 293 57 294 644 645 cell_1rw
* cell instance $14508 r0 *1 81.075,76.44
X$14508 295 57 296 644 645 cell_1rw
* cell instance $14509 r0 *1 81.78,76.44
X$14509 297 57 298 644 645 cell_1rw
* cell instance $14510 r0 *1 82.485,76.44
X$14510 299 57 300 644 645 cell_1rw
* cell instance $14511 r0 *1 83.19,76.44
X$14511 301 57 302 644 645 cell_1rw
* cell instance $14512 r0 *1 83.895,76.44
X$14512 303 57 304 644 645 cell_1rw
* cell instance $14513 r0 *1 84.6,76.44
X$14513 305 57 306 644 645 cell_1rw
* cell instance $14514 r0 *1 85.305,76.44
X$14514 307 57 308 644 645 cell_1rw
* cell instance $14515 r0 *1 86.01,76.44
X$14515 309 57 310 644 645 cell_1rw
* cell instance $14516 r0 *1 86.715,76.44
X$14516 311 57 312 644 645 cell_1rw
* cell instance $14517 r0 *1 87.42,76.44
X$14517 313 57 314 644 645 cell_1rw
* cell instance $14518 r0 *1 88.125,76.44
X$14518 315 57 316 644 645 cell_1rw
* cell instance $14519 r0 *1 88.83,76.44
X$14519 317 57 318 644 645 cell_1rw
* cell instance $14520 r0 *1 89.535,76.44
X$14520 319 57 320 644 645 cell_1rw
* cell instance $14521 r0 *1 90.24,76.44
X$14521 321 57 323 644 645 cell_1rw
* cell instance $14522 r0 *1 90.945,76.44
X$14522 324 57 325 644 645 cell_1rw
* cell instance $14523 r0 *1 91.65,76.44
X$14523 326 57 327 644 645 cell_1rw
* cell instance $14524 r0 *1 92.355,76.44
X$14524 328 57 329 644 645 cell_1rw
* cell instance $14525 r0 *1 93.06,76.44
X$14525 330 57 331 644 645 cell_1rw
* cell instance $14526 r0 *1 93.765,76.44
X$14526 332 57 333 644 645 cell_1rw
* cell instance $14527 r0 *1 94.47,76.44
X$14527 334 57 335 644 645 cell_1rw
* cell instance $14528 r0 *1 95.175,76.44
X$14528 336 57 337 644 645 cell_1rw
* cell instance $14529 r0 *1 95.88,76.44
X$14529 338 57 339 644 645 cell_1rw
* cell instance $14530 r0 *1 96.585,76.44
X$14530 340 57 341 644 645 cell_1rw
* cell instance $14531 r0 *1 97.29,76.44
X$14531 342 57 343 644 645 cell_1rw
* cell instance $14532 r0 *1 97.995,76.44
X$14532 344 57 345 644 645 cell_1rw
* cell instance $14533 r0 *1 98.7,76.44
X$14533 346 57 347 644 645 cell_1rw
* cell instance $14534 r0 *1 99.405,76.44
X$14534 348 57 349 644 645 cell_1rw
* cell instance $14535 r0 *1 100.11,76.44
X$14535 350 57 351 644 645 cell_1rw
* cell instance $14536 r0 *1 100.815,76.44
X$14536 352 57 353 644 645 cell_1rw
* cell instance $14537 r0 *1 101.52,76.44
X$14537 354 57 355 644 645 cell_1rw
* cell instance $14538 r0 *1 102.225,76.44
X$14538 356 57 357 644 645 cell_1rw
* cell instance $14539 r0 *1 102.93,76.44
X$14539 358 57 359 644 645 cell_1rw
* cell instance $14540 r0 *1 103.635,76.44
X$14540 360 57 361 644 645 cell_1rw
* cell instance $14541 r0 *1 104.34,76.44
X$14541 362 57 363 644 645 cell_1rw
* cell instance $14542 r0 *1 105.045,76.44
X$14542 364 57 365 644 645 cell_1rw
* cell instance $14543 r0 *1 105.75,76.44
X$14543 366 57 367 644 645 cell_1rw
* cell instance $14544 r0 *1 106.455,76.44
X$14544 368 57 369 644 645 cell_1rw
* cell instance $14545 r0 *1 107.16,76.44
X$14545 370 57 371 644 645 cell_1rw
* cell instance $14546 r0 *1 107.865,76.44
X$14546 372 57 373 644 645 cell_1rw
* cell instance $14547 r0 *1 108.57,76.44
X$14547 374 57 375 644 645 cell_1rw
* cell instance $14548 r0 *1 109.275,76.44
X$14548 376 57 377 644 645 cell_1rw
* cell instance $14549 r0 *1 109.98,76.44
X$14549 378 57 379 644 645 cell_1rw
* cell instance $14550 r0 *1 110.685,76.44
X$14550 380 57 381 644 645 cell_1rw
* cell instance $14551 r0 *1 111.39,76.44
X$14551 382 57 383 644 645 cell_1rw
* cell instance $14552 r0 *1 112.095,76.44
X$14552 384 57 385 644 645 cell_1rw
* cell instance $14553 r0 *1 112.8,76.44
X$14553 386 57 387 644 645 cell_1rw
* cell instance $14554 r0 *1 113.505,76.44
X$14554 388 57 389 644 645 cell_1rw
* cell instance $14555 r0 *1 114.21,76.44
X$14555 390 57 391 644 645 cell_1rw
* cell instance $14556 r0 *1 114.915,76.44
X$14556 392 57 393 644 645 cell_1rw
* cell instance $14557 r0 *1 115.62,76.44
X$14557 394 57 395 644 645 cell_1rw
* cell instance $14558 r0 *1 116.325,76.44
X$14558 396 57 397 644 645 cell_1rw
* cell instance $14559 r0 *1 117.03,76.44
X$14559 398 57 399 644 645 cell_1rw
* cell instance $14560 r0 *1 117.735,76.44
X$14560 400 57 401 644 645 cell_1rw
* cell instance $14561 r0 *1 118.44,76.44
X$14561 402 57 403 644 645 cell_1rw
* cell instance $14562 r0 *1 119.145,76.44
X$14562 404 57 405 644 645 cell_1rw
* cell instance $14563 r0 *1 119.85,76.44
X$14563 406 57 407 644 645 cell_1rw
* cell instance $14564 r0 *1 120.555,76.44
X$14564 408 57 409 644 645 cell_1rw
* cell instance $14565 r0 *1 121.26,76.44
X$14565 410 57 411 644 645 cell_1rw
* cell instance $14566 r0 *1 121.965,76.44
X$14566 412 57 413 644 645 cell_1rw
* cell instance $14567 r0 *1 122.67,76.44
X$14567 414 57 415 644 645 cell_1rw
* cell instance $14568 r0 *1 123.375,76.44
X$14568 416 57 417 644 645 cell_1rw
* cell instance $14569 r0 *1 124.08,76.44
X$14569 418 57 419 644 645 cell_1rw
* cell instance $14570 r0 *1 124.785,76.44
X$14570 420 57 421 644 645 cell_1rw
* cell instance $14571 r0 *1 125.49,76.44
X$14571 422 57 423 644 645 cell_1rw
* cell instance $14572 r0 *1 126.195,76.44
X$14572 424 57 425 644 645 cell_1rw
* cell instance $14573 r0 *1 126.9,76.44
X$14573 426 57 427 644 645 cell_1rw
* cell instance $14574 r0 *1 127.605,76.44
X$14574 428 57 429 644 645 cell_1rw
* cell instance $14575 r0 *1 128.31,76.44
X$14575 430 57 431 644 645 cell_1rw
* cell instance $14576 r0 *1 129.015,76.44
X$14576 432 57 433 644 645 cell_1rw
* cell instance $14577 r0 *1 129.72,76.44
X$14577 434 57 435 644 645 cell_1rw
* cell instance $14578 r0 *1 130.425,76.44
X$14578 436 57 437 644 645 cell_1rw
* cell instance $14579 r0 *1 131.13,76.44
X$14579 438 57 439 644 645 cell_1rw
* cell instance $14580 r0 *1 131.835,76.44
X$14580 440 57 441 644 645 cell_1rw
* cell instance $14581 r0 *1 132.54,76.44
X$14581 442 57 443 644 645 cell_1rw
* cell instance $14582 r0 *1 133.245,76.44
X$14582 444 57 445 644 645 cell_1rw
* cell instance $14583 r0 *1 133.95,76.44
X$14583 446 57 447 644 645 cell_1rw
* cell instance $14584 r0 *1 134.655,76.44
X$14584 448 57 449 644 645 cell_1rw
* cell instance $14585 r0 *1 135.36,76.44
X$14585 450 57 451 644 645 cell_1rw
* cell instance $14586 r0 *1 136.065,76.44
X$14586 452 57 453 644 645 cell_1rw
* cell instance $14587 r0 *1 136.77,76.44
X$14587 454 57 455 644 645 cell_1rw
* cell instance $14588 r0 *1 137.475,76.44
X$14588 456 57 457 644 645 cell_1rw
* cell instance $14589 r0 *1 138.18,76.44
X$14589 458 57 459 644 645 cell_1rw
* cell instance $14590 r0 *1 138.885,76.44
X$14590 460 57 461 644 645 cell_1rw
* cell instance $14591 r0 *1 139.59,76.44
X$14591 462 57 463 644 645 cell_1rw
* cell instance $14592 r0 *1 140.295,76.44
X$14592 464 57 465 644 645 cell_1rw
* cell instance $14593 r0 *1 141,76.44
X$14593 466 57 467 644 645 cell_1rw
* cell instance $14594 r0 *1 141.705,76.44
X$14594 468 57 469 644 645 cell_1rw
* cell instance $14595 r0 *1 142.41,76.44
X$14595 470 57 471 644 645 cell_1rw
* cell instance $14596 r0 *1 143.115,76.44
X$14596 472 57 473 644 645 cell_1rw
* cell instance $14597 r0 *1 143.82,76.44
X$14597 474 57 475 644 645 cell_1rw
* cell instance $14598 r0 *1 144.525,76.44
X$14598 476 57 477 644 645 cell_1rw
* cell instance $14599 r0 *1 145.23,76.44
X$14599 478 57 479 644 645 cell_1rw
* cell instance $14600 r0 *1 145.935,76.44
X$14600 480 57 481 644 645 cell_1rw
* cell instance $14601 r0 *1 146.64,76.44
X$14601 482 57 483 644 645 cell_1rw
* cell instance $14602 r0 *1 147.345,76.44
X$14602 484 57 485 644 645 cell_1rw
* cell instance $14603 r0 *1 148.05,76.44
X$14603 486 57 487 644 645 cell_1rw
* cell instance $14604 r0 *1 148.755,76.44
X$14604 488 57 489 644 645 cell_1rw
* cell instance $14605 r0 *1 149.46,76.44
X$14605 490 57 491 644 645 cell_1rw
* cell instance $14606 r0 *1 150.165,76.44
X$14606 492 57 493 644 645 cell_1rw
* cell instance $14607 r0 *1 150.87,76.44
X$14607 494 57 495 644 645 cell_1rw
* cell instance $14608 r0 *1 151.575,76.44
X$14608 496 57 497 644 645 cell_1rw
* cell instance $14609 r0 *1 152.28,76.44
X$14609 498 57 499 644 645 cell_1rw
* cell instance $14610 r0 *1 152.985,76.44
X$14610 500 57 501 644 645 cell_1rw
* cell instance $14611 r0 *1 153.69,76.44
X$14611 502 57 503 644 645 cell_1rw
* cell instance $14612 r0 *1 154.395,76.44
X$14612 504 57 505 644 645 cell_1rw
* cell instance $14613 r0 *1 155.1,76.44
X$14613 506 57 507 644 645 cell_1rw
* cell instance $14614 r0 *1 155.805,76.44
X$14614 508 57 509 644 645 cell_1rw
* cell instance $14615 r0 *1 156.51,76.44
X$14615 510 57 511 644 645 cell_1rw
* cell instance $14616 r0 *1 157.215,76.44
X$14616 512 57 513 644 645 cell_1rw
* cell instance $14617 r0 *1 157.92,76.44
X$14617 514 57 515 644 645 cell_1rw
* cell instance $14618 r0 *1 158.625,76.44
X$14618 516 57 517 644 645 cell_1rw
* cell instance $14619 r0 *1 159.33,76.44
X$14619 518 57 519 644 645 cell_1rw
* cell instance $14620 r0 *1 160.035,76.44
X$14620 520 57 521 644 645 cell_1rw
* cell instance $14621 r0 *1 160.74,76.44
X$14621 522 57 523 644 645 cell_1rw
* cell instance $14622 r0 *1 161.445,76.44
X$14622 524 57 525 644 645 cell_1rw
* cell instance $14623 r0 *1 162.15,76.44
X$14623 526 57 527 644 645 cell_1rw
* cell instance $14624 r0 *1 162.855,76.44
X$14624 528 57 529 644 645 cell_1rw
* cell instance $14625 r0 *1 163.56,76.44
X$14625 530 57 531 644 645 cell_1rw
* cell instance $14626 r0 *1 164.265,76.44
X$14626 532 57 533 644 645 cell_1rw
* cell instance $14627 r0 *1 164.97,76.44
X$14627 534 57 535 644 645 cell_1rw
* cell instance $14628 r0 *1 165.675,76.44
X$14628 536 57 537 644 645 cell_1rw
* cell instance $14629 r0 *1 166.38,76.44
X$14629 538 57 539 644 645 cell_1rw
* cell instance $14630 r0 *1 167.085,76.44
X$14630 540 57 541 644 645 cell_1rw
* cell instance $14631 r0 *1 167.79,76.44
X$14631 542 57 543 644 645 cell_1rw
* cell instance $14632 r0 *1 168.495,76.44
X$14632 544 57 545 644 645 cell_1rw
* cell instance $14633 r0 *1 169.2,76.44
X$14633 546 57 547 644 645 cell_1rw
* cell instance $14634 r0 *1 169.905,76.44
X$14634 548 57 549 644 645 cell_1rw
* cell instance $14635 r0 *1 170.61,76.44
X$14635 550 57 551 644 645 cell_1rw
* cell instance $14636 r0 *1 171.315,76.44
X$14636 552 57 553 644 645 cell_1rw
* cell instance $14637 r0 *1 172.02,76.44
X$14637 554 57 555 644 645 cell_1rw
* cell instance $14638 r0 *1 172.725,76.44
X$14638 556 57 557 644 645 cell_1rw
* cell instance $14639 r0 *1 173.43,76.44
X$14639 558 57 559 644 645 cell_1rw
* cell instance $14640 r0 *1 174.135,76.44
X$14640 560 57 561 644 645 cell_1rw
* cell instance $14641 r0 *1 174.84,76.44
X$14641 562 57 563 644 645 cell_1rw
* cell instance $14642 r0 *1 175.545,76.44
X$14642 564 57 565 644 645 cell_1rw
* cell instance $14643 r0 *1 176.25,76.44
X$14643 566 57 567 644 645 cell_1rw
* cell instance $14644 r0 *1 176.955,76.44
X$14644 568 57 569 644 645 cell_1rw
* cell instance $14645 r0 *1 177.66,76.44
X$14645 570 57 571 644 645 cell_1rw
* cell instance $14646 r0 *1 178.365,76.44
X$14646 572 57 573 644 645 cell_1rw
* cell instance $14647 r0 *1 179.07,76.44
X$14647 574 57 575 644 645 cell_1rw
* cell instance $14648 r0 *1 179.775,76.44
X$14648 576 57 577 644 645 cell_1rw
* cell instance $14649 r0 *1 180.48,76.44
X$14649 578 57 579 644 645 cell_1rw
* cell instance $14650 m0 *1 0.705,79.17
X$14650 67 58 68 644 645 cell_1rw
* cell instance $14651 m0 *1 0,79.17
X$14651 65 58 66 644 645 cell_1rw
* cell instance $14652 m0 *1 1.41,79.17
X$14652 69 58 70 644 645 cell_1rw
* cell instance $14653 m0 *1 2.115,79.17
X$14653 71 58 72 644 645 cell_1rw
* cell instance $14654 m0 *1 2.82,79.17
X$14654 73 58 74 644 645 cell_1rw
* cell instance $14655 m0 *1 3.525,79.17
X$14655 75 58 76 644 645 cell_1rw
* cell instance $14656 m0 *1 4.23,79.17
X$14656 77 58 78 644 645 cell_1rw
* cell instance $14657 m0 *1 4.935,79.17
X$14657 79 58 80 644 645 cell_1rw
* cell instance $14658 m0 *1 5.64,79.17
X$14658 81 58 82 644 645 cell_1rw
* cell instance $14659 m0 *1 6.345,79.17
X$14659 83 58 84 644 645 cell_1rw
* cell instance $14660 m0 *1 7.05,79.17
X$14660 85 58 86 644 645 cell_1rw
* cell instance $14661 m0 *1 7.755,79.17
X$14661 87 58 88 644 645 cell_1rw
* cell instance $14662 m0 *1 8.46,79.17
X$14662 89 58 90 644 645 cell_1rw
* cell instance $14663 m0 *1 9.165,79.17
X$14663 91 58 92 644 645 cell_1rw
* cell instance $14664 m0 *1 9.87,79.17
X$14664 93 58 94 644 645 cell_1rw
* cell instance $14665 m0 *1 10.575,79.17
X$14665 95 58 96 644 645 cell_1rw
* cell instance $14666 m0 *1 11.28,79.17
X$14666 97 58 98 644 645 cell_1rw
* cell instance $14667 m0 *1 11.985,79.17
X$14667 99 58 100 644 645 cell_1rw
* cell instance $14668 m0 *1 12.69,79.17
X$14668 101 58 102 644 645 cell_1rw
* cell instance $14669 m0 *1 13.395,79.17
X$14669 103 58 104 644 645 cell_1rw
* cell instance $14670 m0 *1 14.1,79.17
X$14670 105 58 106 644 645 cell_1rw
* cell instance $14671 m0 *1 14.805,79.17
X$14671 107 58 108 644 645 cell_1rw
* cell instance $14672 m0 *1 15.51,79.17
X$14672 109 58 110 644 645 cell_1rw
* cell instance $14673 m0 *1 16.215,79.17
X$14673 111 58 112 644 645 cell_1rw
* cell instance $14674 m0 *1 16.92,79.17
X$14674 113 58 114 644 645 cell_1rw
* cell instance $14675 m0 *1 17.625,79.17
X$14675 115 58 116 644 645 cell_1rw
* cell instance $14676 m0 *1 18.33,79.17
X$14676 117 58 118 644 645 cell_1rw
* cell instance $14677 m0 *1 19.035,79.17
X$14677 119 58 120 644 645 cell_1rw
* cell instance $14678 m0 *1 19.74,79.17
X$14678 121 58 122 644 645 cell_1rw
* cell instance $14679 m0 *1 20.445,79.17
X$14679 123 58 124 644 645 cell_1rw
* cell instance $14680 m0 *1 21.15,79.17
X$14680 125 58 126 644 645 cell_1rw
* cell instance $14681 m0 *1 21.855,79.17
X$14681 127 58 128 644 645 cell_1rw
* cell instance $14682 m0 *1 22.56,79.17
X$14682 129 58 130 644 645 cell_1rw
* cell instance $14683 m0 *1 23.265,79.17
X$14683 131 58 132 644 645 cell_1rw
* cell instance $14684 m0 *1 23.97,79.17
X$14684 133 58 134 644 645 cell_1rw
* cell instance $14685 m0 *1 24.675,79.17
X$14685 135 58 136 644 645 cell_1rw
* cell instance $14686 m0 *1 25.38,79.17
X$14686 137 58 138 644 645 cell_1rw
* cell instance $14687 m0 *1 26.085,79.17
X$14687 139 58 140 644 645 cell_1rw
* cell instance $14688 m0 *1 26.79,79.17
X$14688 141 58 142 644 645 cell_1rw
* cell instance $14689 m0 *1 27.495,79.17
X$14689 143 58 144 644 645 cell_1rw
* cell instance $14690 m0 *1 28.2,79.17
X$14690 145 58 146 644 645 cell_1rw
* cell instance $14691 m0 *1 28.905,79.17
X$14691 147 58 148 644 645 cell_1rw
* cell instance $14692 m0 *1 29.61,79.17
X$14692 149 58 150 644 645 cell_1rw
* cell instance $14693 m0 *1 30.315,79.17
X$14693 151 58 152 644 645 cell_1rw
* cell instance $14694 m0 *1 31.02,79.17
X$14694 153 58 154 644 645 cell_1rw
* cell instance $14695 m0 *1 31.725,79.17
X$14695 155 58 156 644 645 cell_1rw
* cell instance $14696 m0 *1 32.43,79.17
X$14696 157 58 158 644 645 cell_1rw
* cell instance $14697 m0 *1 33.135,79.17
X$14697 159 58 160 644 645 cell_1rw
* cell instance $14698 m0 *1 33.84,79.17
X$14698 161 58 162 644 645 cell_1rw
* cell instance $14699 m0 *1 34.545,79.17
X$14699 163 58 164 644 645 cell_1rw
* cell instance $14700 m0 *1 35.25,79.17
X$14700 165 58 166 644 645 cell_1rw
* cell instance $14701 m0 *1 35.955,79.17
X$14701 167 58 168 644 645 cell_1rw
* cell instance $14702 m0 *1 36.66,79.17
X$14702 169 58 170 644 645 cell_1rw
* cell instance $14703 m0 *1 37.365,79.17
X$14703 171 58 172 644 645 cell_1rw
* cell instance $14704 m0 *1 38.07,79.17
X$14704 173 58 174 644 645 cell_1rw
* cell instance $14705 m0 *1 38.775,79.17
X$14705 175 58 176 644 645 cell_1rw
* cell instance $14706 m0 *1 39.48,79.17
X$14706 177 58 178 644 645 cell_1rw
* cell instance $14707 m0 *1 40.185,79.17
X$14707 179 58 180 644 645 cell_1rw
* cell instance $14708 m0 *1 40.89,79.17
X$14708 181 58 182 644 645 cell_1rw
* cell instance $14709 m0 *1 41.595,79.17
X$14709 183 58 184 644 645 cell_1rw
* cell instance $14710 m0 *1 42.3,79.17
X$14710 185 58 186 644 645 cell_1rw
* cell instance $14711 m0 *1 43.005,79.17
X$14711 187 58 188 644 645 cell_1rw
* cell instance $14712 m0 *1 43.71,79.17
X$14712 189 58 190 644 645 cell_1rw
* cell instance $14713 m0 *1 44.415,79.17
X$14713 191 58 192 644 645 cell_1rw
* cell instance $14714 m0 *1 45.12,79.17
X$14714 193 58 194 644 645 cell_1rw
* cell instance $14715 m0 *1 45.825,79.17
X$14715 195 58 196 644 645 cell_1rw
* cell instance $14716 m0 *1 46.53,79.17
X$14716 197 58 198 644 645 cell_1rw
* cell instance $14717 m0 *1 47.235,79.17
X$14717 199 58 200 644 645 cell_1rw
* cell instance $14718 m0 *1 47.94,79.17
X$14718 201 58 202 644 645 cell_1rw
* cell instance $14719 m0 *1 48.645,79.17
X$14719 203 58 204 644 645 cell_1rw
* cell instance $14720 m0 *1 49.35,79.17
X$14720 205 58 206 644 645 cell_1rw
* cell instance $14721 m0 *1 50.055,79.17
X$14721 207 58 208 644 645 cell_1rw
* cell instance $14722 m0 *1 50.76,79.17
X$14722 209 58 210 644 645 cell_1rw
* cell instance $14723 m0 *1 51.465,79.17
X$14723 211 58 212 644 645 cell_1rw
* cell instance $14724 m0 *1 52.17,79.17
X$14724 213 58 214 644 645 cell_1rw
* cell instance $14725 m0 *1 52.875,79.17
X$14725 215 58 216 644 645 cell_1rw
* cell instance $14726 m0 *1 53.58,79.17
X$14726 217 58 218 644 645 cell_1rw
* cell instance $14727 m0 *1 54.285,79.17
X$14727 219 58 220 644 645 cell_1rw
* cell instance $14728 m0 *1 54.99,79.17
X$14728 221 58 222 644 645 cell_1rw
* cell instance $14729 m0 *1 55.695,79.17
X$14729 223 58 224 644 645 cell_1rw
* cell instance $14730 m0 *1 56.4,79.17
X$14730 225 58 226 644 645 cell_1rw
* cell instance $14731 m0 *1 57.105,79.17
X$14731 227 58 228 644 645 cell_1rw
* cell instance $14732 m0 *1 57.81,79.17
X$14732 229 58 230 644 645 cell_1rw
* cell instance $14733 m0 *1 58.515,79.17
X$14733 231 58 232 644 645 cell_1rw
* cell instance $14734 m0 *1 59.22,79.17
X$14734 233 58 234 644 645 cell_1rw
* cell instance $14735 m0 *1 59.925,79.17
X$14735 235 58 236 644 645 cell_1rw
* cell instance $14736 m0 *1 60.63,79.17
X$14736 237 58 238 644 645 cell_1rw
* cell instance $14737 m0 *1 61.335,79.17
X$14737 239 58 240 644 645 cell_1rw
* cell instance $14738 m0 *1 62.04,79.17
X$14738 241 58 242 644 645 cell_1rw
* cell instance $14739 m0 *1 62.745,79.17
X$14739 243 58 244 644 645 cell_1rw
* cell instance $14740 m0 *1 63.45,79.17
X$14740 245 58 246 644 645 cell_1rw
* cell instance $14741 m0 *1 64.155,79.17
X$14741 247 58 248 644 645 cell_1rw
* cell instance $14742 m0 *1 64.86,79.17
X$14742 249 58 250 644 645 cell_1rw
* cell instance $14743 m0 *1 65.565,79.17
X$14743 251 58 252 644 645 cell_1rw
* cell instance $14744 m0 *1 66.27,79.17
X$14744 253 58 254 644 645 cell_1rw
* cell instance $14745 m0 *1 66.975,79.17
X$14745 255 58 256 644 645 cell_1rw
* cell instance $14746 m0 *1 67.68,79.17
X$14746 257 58 258 644 645 cell_1rw
* cell instance $14747 m0 *1 68.385,79.17
X$14747 259 58 260 644 645 cell_1rw
* cell instance $14748 m0 *1 69.09,79.17
X$14748 261 58 262 644 645 cell_1rw
* cell instance $14749 m0 *1 69.795,79.17
X$14749 263 58 264 644 645 cell_1rw
* cell instance $14750 m0 *1 70.5,79.17
X$14750 265 58 266 644 645 cell_1rw
* cell instance $14751 m0 *1 71.205,79.17
X$14751 267 58 268 644 645 cell_1rw
* cell instance $14752 m0 *1 71.91,79.17
X$14752 269 58 270 644 645 cell_1rw
* cell instance $14753 m0 *1 72.615,79.17
X$14753 271 58 272 644 645 cell_1rw
* cell instance $14754 m0 *1 73.32,79.17
X$14754 273 58 274 644 645 cell_1rw
* cell instance $14755 m0 *1 74.025,79.17
X$14755 275 58 276 644 645 cell_1rw
* cell instance $14756 m0 *1 74.73,79.17
X$14756 277 58 278 644 645 cell_1rw
* cell instance $14757 m0 *1 75.435,79.17
X$14757 279 58 280 644 645 cell_1rw
* cell instance $14758 m0 *1 76.14,79.17
X$14758 281 58 282 644 645 cell_1rw
* cell instance $14759 m0 *1 76.845,79.17
X$14759 283 58 284 644 645 cell_1rw
* cell instance $14760 m0 *1 77.55,79.17
X$14760 285 58 286 644 645 cell_1rw
* cell instance $14761 m0 *1 78.255,79.17
X$14761 287 58 288 644 645 cell_1rw
* cell instance $14762 m0 *1 78.96,79.17
X$14762 289 58 290 644 645 cell_1rw
* cell instance $14763 m0 *1 79.665,79.17
X$14763 291 58 292 644 645 cell_1rw
* cell instance $14764 m0 *1 80.37,79.17
X$14764 293 58 294 644 645 cell_1rw
* cell instance $14765 m0 *1 81.075,79.17
X$14765 295 58 296 644 645 cell_1rw
* cell instance $14766 m0 *1 81.78,79.17
X$14766 297 58 298 644 645 cell_1rw
* cell instance $14767 m0 *1 82.485,79.17
X$14767 299 58 300 644 645 cell_1rw
* cell instance $14768 m0 *1 83.19,79.17
X$14768 301 58 302 644 645 cell_1rw
* cell instance $14769 m0 *1 83.895,79.17
X$14769 303 58 304 644 645 cell_1rw
* cell instance $14770 m0 *1 84.6,79.17
X$14770 305 58 306 644 645 cell_1rw
* cell instance $14771 m0 *1 85.305,79.17
X$14771 307 58 308 644 645 cell_1rw
* cell instance $14772 m0 *1 86.01,79.17
X$14772 309 58 310 644 645 cell_1rw
* cell instance $14773 m0 *1 86.715,79.17
X$14773 311 58 312 644 645 cell_1rw
* cell instance $14774 m0 *1 87.42,79.17
X$14774 313 58 314 644 645 cell_1rw
* cell instance $14775 m0 *1 88.125,79.17
X$14775 315 58 316 644 645 cell_1rw
* cell instance $14776 m0 *1 88.83,79.17
X$14776 317 58 318 644 645 cell_1rw
* cell instance $14777 m0 *1 89.535,79.17
X$14777 319 58 320 644 645 cell_1rw
* cell instance $14778 m0 *1 90.24,79.17
X$14778 321 58 323 644 645 cell_1rw
* cell instance $14779 m0 *1 90.945,79.17
X$14779 324 58 325 644 645 cell_1rw
* cell instance $14780 m0 *1 91.65,79.17
X$14780 326 58 327 644 645 cell_1rw
* cell instance $14781 m0 *1 92.355,79.17
X$14781 328 58 329 644 645 cell_1rw
* cell instance $14782 m0 *1 93.06,79.17
X$14782 330 58 331 644 645 cell_1rw
* cell instance $14783 m0 *1 93.765,79.17
X$14783 332 58 333 644 645 cell_1rw
* cell instance $14784 m0 *1 94.47,79.17
X$14784 334 58 335 644 645 cell_1rw
* cell instance $14785 m0 *1 95.175,79.17
X$14785 336 58 337 644 645 cell_1rw
* cell instance $14786 m0 *1 95.88,79.17
X$14786 338 58 339 644 645 cell_1rw
* cell instance $14787 m0 *1 96.585,79.17
X$14787 340 58 341 644 645 cell_1rw
* cell instance $14788 m0 *1 97.29,79.17
X$14788 342 58 343 644 645 cell_1rw
* cell instance $14789 m0 *1 97.995,79.17
X$14789 344 58 345 644 645 cell_1rw
* cell instance $14790 m0 *1 98.7,79.17
X$14790 346 58 347 644 645 cell_1rw
* cell instance $14791 m0 *1 99.405,79.17
X$14791 348 58 349 644 645 cell_1rw
* cell instance $14792 m0 *1 100.11,79.17
X$14792 350 58 351 644 645 cell_1rw
* cell instance $14793 m0 *1 100.815,79.17
X$14793 352 58 353 644 645 cell_1rw
* cell instance $14794 m0 *1 101.52,79.17
X$14794 354 58 355 644 645 cell_1rw
* cell instance $14795 m0 *1 102.225,79.17
X$14795 356 58 357 644 645 cell_1rw
* cell instance $14796 m0 *1 102.93,79.17
X$14796 358 58 359 644 645 cell_1rw
* cell instance $14797 m0 *1 103.635,79.17
X$14797 360 58 361 644 645 cell_1rw
* cell instance $14798 m0 *1 104.34,79.17
X$14798 362 58 363 644 645 cell_1rw
* cell instance $14799 m0 *1 105.045,79.17
X$14799 364 58 365 644 645 cell_1rw
* cell instance $14800 m0 *1 105.75,79.17
X$14800 366 58 367 644 645 cell_1rw
* cell instance $14801 m0 *1 106.455,79.17
X$14801 368 58 369 644 645 cell_1rw
* cell instance $14802 m0 *1 107.16,79.17
X$14802 370 58 371 644 645 cell_1rw
* cell instance $14803 m0 *1 107.865,79.17
X$14803 372 58 373 644 645 cell_1rw
* cell instance $14804 m0 *1 108.57,79.17
X$14804 374 58 375 644 645 cell_1rw
* cell instance $14805 m0 *1 109.275,79.17
X$14805 376 58 377 644 645 cell_1rw
* cell instance $14806 m0 *1 109.98,79.17
X$14806 378 58 379 644 645 cell_1rw
* cell instance $14807 m0 *1 110.685,79.17
X$14807 380 58 381 644 645 cell_1rw
* cell instance $14808 m0 *1 111.39,79.17
X$14808 382 58 383 644 645 cell_1rw
* cell instance $14809 m0 *1 112.095,79.17
X$14809 384 58 385 644 645 cell_1rw
* cell instance $14810 m0 *1 112.8,79.17
X$14810 386 58 387 644 645 cell_1rw
* cell instance $14811 m0 *1 113.505,79.17
X$14811 388 58 389 644 645 cell_1rw
* cell instance $14812 m0 *1 114.21,79.17
X$14812 390 58 391 644 645 cell_1rw
* cell instance $14813 m0 *1 114.915,79.17
X$14813 392 58 393 644 645 cell_1rw
* cell instance $14814 m0 *1 115.62,79.17
X$14814 394 58 395 644 645 cell_1rw
* cell instance $14815 m0 *1 116.325,79.17
X$14815 396 58 397 644 645 cell_1rw
* cell instance $14816 m0 *1 117.03,79.17
X$14816 398 58 399 644 645 cell_1rw
* cell instance $14817 m0 *1 117.735,79.17
X$14817 400 58 401 644 645 cell_1rw
* cell instance $14818 m0 *1 118.44,79.17
X$14818 402 58 403 644 645 cell_1rw
* cell instance $14819 m0 *1 119.145,79.17
X$14819 404 58 405 644 645 cell_1rw
* cell instance $14820 m0 *1 119.85,79.17
X$14820 406 58 407 644 645 cell_1rw
* cell instance $14821 m0 *1 120.555,79.17
X$14821 408 58 409 644 645 cell_1rw
* cell instance $14822 m0 *1 121.26,79.17
X$14822 410 58 411 644 645 cell_1rw
* cell instance $14823 m0 *1 121.965,79.17
X$14823 412 58 413 644 645 cell_1rw
* cell instance $14824 m0 *1 122.67,79.17
X$14824 414 58 415 644 645 cell_1rw
* cell instance $14825 m0 *1 123.375,79.17
X$14825 416 58 417 644 645 cell_1rw
* cell instance $14826 m0 *1 124.08,79.17
X$14826 418 58 419 644 645 cell_1rw
* cell instance $14827 m0 *1 124.785,79.17
X$14827 420 58 421 644 645 cell_1rw
* cell instance $14828 m0 *1 125.49,79.17
X$14828 422 58 423 644 645 cell_1rw
* cell instance $14829 m0 *1 126.195,79.17
X$14829 424 58 425 644 645 cell_1rw
* cell instance $14830 m0 *1 126.9,79.17
X$14830 426 58 427 644 645 cell_1rw
* cell instance $14831 m0 *1 127.605,79.17
X$14831 428 58 429 644 645 cell_1rw
* cell instance $14832 m0 *1 128.31,79.17
X$14832 430 58 431 644 645 cell_1rw
* cell instance $14833 m0 *1 129.015,79.17
X$14833 432 58 433 644 645 cell_1rw
* cell instance $14834 m0 *1 129.72,79.17
X$14834 434 58 435 644 645 cell_1rw
* cell instance $14835 m0 *1 130.425,79.17
X$14835 436 58 437 644 645 cell_1rw
* cell instance $14836 m0 *1 131.13,79.17
X$14836 438 58 439 644 645 cell_1rw
* cell instance $14837 m0 *1 131.835,79.17
X$14837 440 58 441 644 645 cell_1rw
* cell instance $14838 m0 *1 132.54,79.17
X$14838 442 58 443 644 645 cell_1rw
* cell instance $14839 m0 *1 133.245,79.17
X$14839 444 58 445 644 645 cell_1rw
* cell instance $14840 m0 *1 133.95,79.17
X$14840 446 58 447 644 645 cell_1rw
* cell instance $14841 m0 *1 134.655,79.17
X$14841 448 58 449 644 645 cell_1rw
* cell instance $14842 m0 *1 135.36,79.17
X$14842 450 58 451 644 645 cell_1rw
* cell instance $14843 m0 *1 136.065,79.17
X$14843 452 58 453 644 645 cell_1rw
* cell instance $14844 m0 *1 136.77,79.17
X$14844 454 58 455 644 645 cell_1rw
* cell instance $14845 m0 *1 137.475,79.17
X$14845 456 58 457 644 645 cell_1rw
* cell instance $14846 m0 *1 138.18,79.17
X$14846 458 58 459 644 645 cell_1rw
* cell instance $14847 m0 *1 138.885,79.17
X$14847 460 58 461 644 645 cell_1rw
* cell instance $14848 m0 *1 139.59,79.17
X$14848 462 58 463 644 645 cell_1rw
* cell instance $14849 m0 *1 140.295,79.17
X$14849 464 58 465 644 645 cell_1rw
* cell instance $14850 m0 *1 141,79.17
X$14850 466 58 467 644 645 cell_1rw
* cell instance $14851 m0 *1 141.705,79.17
X$14851 468 58 469 644 645 cell_1rw
* cell instance $14852 m0 *1 142.41,79.17
X$14852 470 58 471 644 645 cell_1rw
* cell instance $14853 m0 *1 143.115,79.17
X$14853 472 58 473 644 645 cell_1rw
* cell instance $14854 m0 *1 143.82,79.17
X$14854 474 58 475 644 645 cell_1rw
* cell instance $14855 m0 *1 144.525,79.17
X$14855 476 58 477 644 645 cell_1rw
* cell instance $14856 m0 *1 145.23,79.17
X$14856 478 58 479 644 645 cell_1rw
* cell instance $14857 m0 *1 145.935,79.17
X$14857 480 58 481 644 645 cell_1rw
* cell instance $14858 m0 *1 146.64,79.17
X$14858 482 58 483 644 645 cell_1rw
* cell instance $14859 m0 *1 147.345,79.17
X$14859 484 58 485 644 645 cell_1rw
* cell instance $14860 m0 *1 148.05,79.17
X$14860 486 58 487 644 645 cell_1rw
* cell instance $14861 m0 *1 148.755,79.17
X$14861 488 58 489 644 645 cell_1rw
* cell instance $14862 m0 *1 149.46,79.17
X$14862 490 58 491 644 645 cell_1rw
* cell instance $14863 m0 *1 150.165,79.17
X$14863 492 58 493 644 645 cell_1rw
* cell instance $14864 m0 *1 150.87,79.17
X$14864 494 58 495 644 645 cell_1rw
* cell instance $14865 m0 *1 151.575,79.17
X$14865 496 58 497 644 645 cell_1rw
* cell instance $14866 m0 *1 152.28,79.17
X$14866 498 58 499 644 645 cell_1rw
* cell instance $14867 m0 *1 152.985,79.17
X$14867 500 58 501 644 645 cell_1rw
* cell instance $14868 m0 *1 153.69,79.17
X$14868 502 58 503 644 645 cell_1rw
* cell instance $14869 m0 *1 154.395,79.17
X$14869 504 58 505 644 645 cell_1rw
* cell instance $14870 m0 *1 155.1,79.17
X$14870 506 58 507 644 645 cell_1rw
* cell instance $14871 m0 *1 155.805,79.17
X$14871 508 58 509 644 645 cell_1rw
* cell instance $14872 m0 *1 156.51,79.17
X$14872 510 58 511 644 645 cell_1rw
* cell instance $14873 m0 *1 157.215,79.17
X$14873 512 58 513 644 645 cell_1rw
* cell instance $14874 m0 *1 157.92,79.17
X$14874 514 58 515 644 645 cell_1rw
* cell instance $14875 m0 *1 158.625,79.17
X$14875 516 58 517 644 645 cell_1rw
* cell instance $14876 m0 *1 159.33,79.17
X$14876 518 58 519 644 645 cell_1rw
* cell instance $14877 m0 *1 160.035,79.17
X$14877 520 58 521 644 645 cell_1rw
* cell instance $14878 m0 *1 160.74,79.17
X$14878 522 58 523 644 645 cell_1rw
* cell instance $14879 m0 *1 161.445,79.17
X$14879 524 58 525 644 645 cell_1rw
* cell instance $14880 m0 *1 162.15,79.17
X$14880 526 58 527 644 645 cell_1rw
* cell instance $14881 m0 *1 162.855,79.17
X$14881 528 58 529 644 645 cell_1rw
* cell instance $14882 m0 *1 163.56,79.17
X$14882 530 58 531 644 645 cell_1rw
* cell instance $14883 m0 *1 164.265,79.17
X$14883 532 58 533 644 645 cell_1rw
* cell instance $14884 m0 *1 164.97,79.17
X$14884 534 58 535 644 645 cell_1rw
* cell instance $14885 m0 *1 165.675,79.17
X$14885 536 58 537 644 645 cell_1rw
* cell instance $14886 m0 *1 166.38,79.17
X$14886 538 58 539 644 645 cell_1rw
* cell instance $14887 m0 *1 167.085,79.17
X$14887 540 58 541 644 645 cell_1rw
* cell instance $14888 m0 *1 167.79,79.17
X$14888 542 58 543 644 645 cell_1rw
* cell instance $14889 m0 *1 168.495,79.17
X$14889 544 58 545 644 645 cell_1rw
* cell instance $14890 m0 *1 169.2,79.17
X$14890 546 58 547 644 645 cell_1rw
* cell instance $14891 m0 *1 169.905,79.17
X$14891 548 58 549 644 645 cell_1rw
* cell instance $14892 m0 *1 170.61,79.17
X$14892 550 58 551 644 645 cell_1rw
* cell instance $14893 m0 *1 171.315,79.17
X$14893 552 58 553 644 645 cell_1rw
* cell instance $14894 m0 *1 172.02,79.17
X$14894 554 58 555 644 645 cell_1rw
* cell instance $14895 m0 *1 172.725,79.17
X$14895 556 58 557 644 645 cell_1rw
* cell instance $14896 m0 *1 173.43,79.17
X$14896 558 58 559 644 645 cell_1rw
* cell instance $14897 m0 *1 174.135,79.17
X$14897 560 58 561 644 645 cell_1rw
* cell instance $14898 m0 *1 174.84,79.17
X$14898 562 58 563 644 645 cell_1rw
* cell instance $14899 m0 *1 175.545,79.17
X$14899 564 58 565 644 645 cell_1rw
* cell instance $14900 m0 *1 176.25,79.17
X$14900 566 58 567 644 645 cell_1rw
* cell instance $14901 m0 *1 176.955,79.17
X$14901 568 58 569 644 645 cell_1rw
* cell instance $14902 m0 *1 177.66,79.17
X$14902 570 58 571 644 645 cell_1rw
* cell instance $14903 m0 *1 178.365,79.17
X$14903 572 58 573 644 645 cell_1rw
* cell instance $14904 m0 *1 179.07,79.17
X$14904 574 58 575 644 645 cell_1rw
* cell instance $14905 m0 *1 179.775,79.17
X$14905 576 58 577 644 645 cell_1rw
* cell instance $14906 m0 *1 180.48,79.17
X$14906 578 58 579 644 645 cell_1rw
* cell instance $14907 r0 *1 0.705,79.17
X$14907 67 59 68 644 645 cell_1rw
* cell instance $14908 r0 *1 0,79.17
X$14908 65 59 66 644 645 cell_1rw
* cell instance $14909 r0 *1 1.41,79.17
X$14909 69 59 70 644 645 cell_1rw
* cell instance $14910 r0 *1 2.115,79.17
X$14910 71 59 72 644 645 cell_1rw
* cell instance $14911 r0 *1 2.82,79.17
X$14911 73 59 74 644 645 cell_1rw
* cell instance $14912 r0 *1 3.525,79.17
X$14912 75 59 76 644 645 cell_1rw
* cell instance $14913 r0 *1 4.23,79.17
X$14913 77 59 78 644 645 cell_1rw
* cell instance $14914 r0 *1 4.935,79.17
X$14914 79 59 80 644 645 cell_1rw
* cell instance $14915 r0 *1 5.64,79.17
X$14915 81 59 82 644 645 cell_1rw
* cell instance $14916 r0 *1 6.345,79.17
X$14916 83 59 84 644 645 cell_1rw
* cell instance $14917 r0 *1 7.05,79.17
X$14917 85 59 86 644 645 cell_1rw
* cell instance $14918 r0 *1 7.755,79.17
X$14918 87 59 88 644 645 cell_1rw
* cell instance $14919 r0 *1 8.46,79.17
X$14919 89 59 90 644 645 cell_1rw
* cell instance $14920 r0 *1 9.165,79.17
X$14920 91 59 92 644 645 cell_1rw
* cell instance $14921 r0 *1 9.87,79.17
X$14921 93 59 94 644 645 cell_1rw
* cell instance $14922 r0 *1 10.575,79.17
X$14922 95 59 96 644 645 cell_1rw
* cell instance $14923 r0 *1 11.28,79.17
X$14923 97 59 98 644 645 cell_1rw
* cell instance $14924 r0 *1 11.985,79.17
X$14924 99 59 100 644 645 cell_1rw
* cell instance $14925 r0 *1 12.69,79.17
X$14925 101 59 102 644 645 cell_1rw
* cell instance $14926 r0 *1 13.395,79.17
X$14926 103 59 104 644 645 cell_1rw
* cell instance $14927 r0 *1 14.1,79.17
X$14927 105 59 106 644 645 cell_1rw
* cell instance $14928 r0 *1 14.805,79.17
X$14928 107 59 108 644 645 cell_1rw
* cell instance $14929 r0 *1 15.51,79.17
X$14929 109 59 110 644 645 cell_1rw
* cell instance $14930 r0 *1 16.215,79.17
X$14930 111 59 112 644 645 cell_1rw
* cell instance $14931 r0 *1 16.92,79.17
X$14931 113 59 114 644 645 cell_1rw
* cell instance $14932 r0 *1 17.625,79.17
X$14932 115 59 116 644 645 cell_1rw
* cell instance $14933 r0 *1 18.33,79.17
X$14933 117 59 118 644 645 cell_1rw
* cell instance $14934 r0 *1 19.035,79.17
X$14934 119 59 120 644 645 cell_1rw
* cell instance $14935 r0 *1 19.74,79.17
X$14935 121 59 122 644 645 cell_1rw
* cell instance $14936 r0 *1 20.445,79.17
X$14936 123 59 124 644 645 cell_1rw
* cell instance $14937 r0 *1 21.15,79.17
X$14937 125 59 126 644 645 cell_1rw
* cell instance $14938 r0 *1 21.855,79.17
X$14938 127 59 128 644 645 cell_1rw
* cell instance $14939 r0 *1 22.56,79.17
X$14939 129 59 130 644 645 cell_1rw
* cell instance $14940 r0 *1 23.265,79.17
X$14940 131 59 132 644 645 cell_1rw
* cell instance $14941 r0 *1 23.97,79.17
X$14941 133 59 134 644 645 cell_1rw
* cell instance $14942 r0 *1 24.675,79.17
X$14942 135 59 136 644 645 cell_1rw
* cell instance $14943 r0 *1 25.38,79.17
X$14943 137 59 138 644 645 cell_1rw
* cell instance $14944 r0 *1 26.085,79.17
X$14944 139 59 140 644 645 cell_1rw
* cell instance $14945 r0 *1 26.79,79.17
X$14945 141 59 142 644 645 cell_1rw
* cell instance $14946 r0 *1 27.495,79.17
X$14946 143 59 144 644 645 cell_1rw
* cell instance $14947 r0 *1 28.2,79.17
X$14947 145 59 146 644 645 cell_1rw
* cell instance $14948 r0 *1 28.905,79.17
X$14948 147 59 148 644 645 cell_1rw
* cell instance $14949 r0 *1 29.61,79.17
X$14949 149 59 150 644 645 cell_1rw
* cell instance $14950 r0 *1 30.315,79.17
X$14950 151 59 152 644 645 cell_1rw
* cell instance $14951 r0 *1 31.02,79.17
X$14951 153 59 154 644 645 cell_1rw
* cell instance $14952 r0 *1 31.725,79.17
X$14952 155 59 156 644 645 cell_1rw
* cell instance $14953 r0 *1 32.43,79.17
X$14953 157 59 158 644 645 cell_1rw
* cell instance $14954 r0 *1 33.135,79.17
X$14954 159 59 160 644 645 cell_1rw
* cell instance $14955 r0 *1 33.84,79.17
X$14955 161 59 162 644 645 cell_1rw
* cell instance $14956 r0 *1 34.545,79.17
X$14956 163 59 164 644 645 cell_1rw
* cell instance $14957 r0 *1 35.25,79.17
X$14957 165 59 166 644 645 cell_1rw
* cell instance $14958 r0 *1 35.955,79.17
X$14958 167 59 168 644 645 cell_1rw
* cell instance $14959 r0 *1 36.66,79.17
X$14959 169 59 170 644 645 cell_1rw
* cell instance $14960 r0 *1 37.365,79.17
X$14960 171 59 172 644 645 cell_1rw
* cell instance $14961 r0 *1 38.07,79.17
X$14961 173 59 174 644 645 cell_1rw
* cell instance $14962 r0 *1 38.775,79.17
X$14962 175 59 176 644 645 cell_1rw
* cell instance $14963 r0 *1 39.48,79.17
X$14963 177 59 178 644 645 cell_1rw
* cell instance $14964 r0 *1 40.185,79.17
X$14964 179 59 180 644 645 cell_1rw
* cell instance $14965 r0 *1 40.89,79.17
X$14965 181 59 182 644 645 cell_1rw
* cell instance $14966 r0 *1 41.595,79.17
X$14966 183 59 184 644 645 cell_1rw
* cell instance $14967 r0 *1 42.3,79.17
X$14967 185 59 186 644 645 cell_1rw
* cell instance $14968 r0 *1 43.005,79.17
X$14968 187 59 188 644 645 cell_1rw
* cell instance $14969 r0 *1 43.71,79.17
X$14969 189 59 190 644 645 cell_1rw
* cell instance $14970 r0 *1 44.415,79.17
X$14970 191 59 192 644 645 cell_1rw
* cell instance $14971 r0 *1 45.12,79.17
X$14971 193 59 194 644 645 cell_1rw
* cell instance $14972 r0 *1 45.825,79.17
X$14972 195 59 196 644 645 cell_1rw
* cell instance $14973 r0 *1 46.53,79.17
X$14973 197 59 198 644 645 cell_1rw
* cell instance $14974 r0 *1 47.235,79.17
X$14974 199 59 200 644 645 cell_1rw
* cell instance $14975 r0 *1 47.94,79.17
X$14975 201 59 202 644 645 cell_1rw
* cell instance $14976 r0 *1 48.645,79.17
X$14976 203 59 204 644 645 cell_1rw
* cell instance $14977 r0 *1 49.35,79.17
X$14977 205 59 206 644 645 cell_1rw
* cell instance $14978 r0 *1 50.055,79.17
X$14978 207 59 208 644 645 cell_1rw
* cell instance $14979 r0 *1 50.76,79.17
X$14979 209 59 210 644 645 cell_1rw
* cell instance $14980 r0 *1 51.465,79.17
X$14980 211 59 212 644 645 cell_1rw
* cell instance $14981 r0 *1 52.17,79.17
X$14981 213 59 214 644 645 cell_1rw
* cell instance $14982 r0 *1 52.875,79.17
X$14982 215 59 216 644 645 cell_1rw
* cell instance $14983 r0 *1 53.58,79.17
X$14983 217 59 218 644 645 cell_1rw
* cell instance $14984 r0 *1 54.285,79.17
X$14984 219 59 220 644 645 cell_1rw
* cell instance $14985 r0 *1 54.99,79.17
X$14985 221 59 222 644 645 cell_1rw
* cell instance $14986 r0 *1 55.695,79.17
X$14986 223 59 224 644 645 cell_1rw
* cell instance $14987 r0 *1 56.4,79.17
X$14987 225 59 226 644 645 cell_1rw
* cell instance $14988 r0 *1 57.105,79.17
X$14988 227 59 228 644 645 cell_1rw
* cell instance $14989 r0 *1 57.81,79.17
X$14989 229 59 230 644 645 cell_1rw
* cell instance $14990 r0 *1 58.515,79.17
X$14990 231 59 232 644 645 cell_1rw
* cell instance $14991 r0 *1 59.22,79.17
X$14991 233 59 234 644 645 cell_1rw
* cell instance $14992 r0 *1 59.925,79.17
X$14992 235 59 236 644 645 cell_1rw
* cell instance $14993 r0 *1 60.63,79.17
X$14993 237 59 238 644 645 cell_1rw
* cell instance $14994 r0 *1 61.335,79.17
X$14994 239 59 240 644 645 cell_1rw
* cell instance $14995 r0 *1 62.04,79.17
X$14995 241 59 242 644 645 cell_1rw
* cell instance $14996 r0 *1 62.745,79.17
X$14996 243 59 244 644 645 cell_1rw
* cell instance $14997 r0 *1 63.45,79.17
X$14997 245 59 246 644 645 cell_1rw
* cell instance $14998 r0 *1 64.155,79.17
X$14998 247 59 248 644 645 cell_1rw
* cell instance $14999 r0 *1 64.86,79.17
X$14999 249 59 250 644 645 cell_1rw
* cell instance $15000 r0 *1 65.565,79.17
X$15000 251 59 252 644 645 cell_1rw
* cell instance $15001 r0 *1 66.27,79.17
X$15001 253 59 254 644 645 cell_1rw
* cell instance $15002 r0 *1 66.975,79.17
X$15002 255 59 256 644 645 cell_1rw
* cell instance $15003 r0 *1 67.68,79.17
X$15003 257 59 258 644 645 cell_1rw
* cell instance $15004 r0 *1 68.385,79.17
X$15004 259 59 260 644 645 cell_1rw
* cell instance $15005 r0 *1 69.09,79.17
X$15005 261 59 262 644 645 cell_1rw
* cell instance $15006 r0 *1 69.795,79.17
X$15006 263 59 264 644 645 cell_1rw
* cell instance $15007 r0 *1 70.5,79.17
X$15007 265 59 266 644 645 cell_1rw
* cell instance $15008 r0 *1 71.205,79.17
X$15008 267 59 268 644 645 cell_1rw
* cell instance $15009 r0 *1 71.91,79.17
X$15009 269 59 270 644 645 cell_1rw
* cell instance $15010 r0 *1 72.615,79.17
X$15010 271 59 272 644 645 cell_1rw
* cell instance $15011 r0 *1 73.32,79.17
X$15011 273 59 274 644 645 cell_1rw
* cell instance $15012 r0 *1 74.025,79.17
X$15012 275 59 276 644 645 cell_1rw
* cell instance $15013 r0 *1 74.73,79.17
X$15013 277 59 278 644 645 cell_1rw
* cell instance $15014 r0 *1 75.435,79.17
X$15014 279 59 280 644 645 cell_1rw
* cell instance $15015 r0 *1 76.14,79.17
X$15015 281 59 282 644 645 cell_1rw
* cell instance $15016 r0 *1 76.845,79.17
X$15016 283 59 284 644 645 cell_1rw
* cell instance $15017 r0 *1 77.55,79.17
X$15017 285 59 286 644 645 cell_1rw
* cell instance $15018 r0 *1 78.255,79.17
X$15018 287 59 288 644 645 cell_1rw
* cell instance $15019 r0 *1 78.96,79.17
X$15019 289 59 290 644 645 cell_1rw
* cell instance $15020 r0 *1 79.665,79.17
X$15020 291 59 292 644 645 cell_1rw
* cell instance $15021 r0 *1 80.37,79.17
X$15021 293 59 294 644 645 cell_1rw
* cell instance $15022 r0 *1 81.075,79.17
X$15022 295 59 296 644 645 cell_1rw
* cell instance $15023 r0 *1 81.78,79.17
X$15023 297 59 298 644 645 cell_1rw
* cell instance $15024 r0 *1 82.485,79.17
X$15024 299 59 300 644 645 cell_1rw
* cell instance $15025 r0 *1 83.19,79.17
X$15025 301 59 302 644 645 cell_1rw
* cell instance $15026 r0 *1 83.895,79.17
X$15026 303 59 304 644 645 cell_1rw
* cell instance $15027 r0 *1 84.6,79.17
X$15027 305 59 306 644 645 cell_1rw
* cell instance $15028 r0 *1 85.305,79.17
X$15028 307 59 308 644 645 cell_1rw
* cell instance $15029 r0 *1 86.01,79.17
X$15029 309 59 310 644 645 cell_1rw
* cell instance $15030 r0 *1 86.715,79.17
X$15030 311 59 312 644 645 cell_1rw
* cell instance $15031 r0 *1 87.42,79.17
X$15031 313 59 314 644 645 cell_1rw
* cell instance $15032 r0 *1 88.125,79.17
X$15032 315 59 316 644 645 cell_1rw
* cell instance $15033 r0 *1 88.83,79.17
X$15033 317 59 318 644 645 cell_1rw
* cell instance $15034 r0 *1 89.535,79.17
X$15034 319 59 320 644 645 cell_1rw
* cell instance $15035 r0 *1 90.24,79.17
X$15035 321 59 323 644 645 cell_1rw
* cell instance $15036 r0 *1 90.945,79.17
X$15036 324 59 325 644 645 cell_1rw
* cell instance $15037 r0 *1 91.65,79.17
X$15037 326 59 327 644 645 cell_1rw
* cell instance $15038 r0 *1 92.355,79.17
X$15038 328 59 329 644 645 cell_1rw
* cell instance $15039 r0 *1 93.06,79.17
X$15039 330 59 331 644 645 cell_1rw
* cell instance $15040 r0 *1 93.765,79.17
X$15040 332 59 333 644 645 cell_1rw
* cell instance $15041 r0 *1 94.47,79.17
X$15041 334 59 335 644 645 cell_1rw
* cell instance $15042 r0 *1 95.175,79.17
X$15042 336 59 337 644 645 cell_1rw
* cell instance $15043 r0 *1 95.88,79.17
X$15043 338 59 339 644 645 cell_1rw
* cell instance $15044 r0 *1 96.585,79.17
X$15044 340 59 341 644 645 cell_1rw
* cell instance $15045 r0 *1 97.29,79.17
X$15045 342 59 343 644 645 cell_1rw
* cell instance $15046 r0 *1 97.995,79.17
X$15046 344 59 345 644 645 cell_1rw
* cell instance $15047 r0 *1 98.7,79.17
X$15047 346 59 347 644 645 cell_1rw
* cell instance $15048 r0 *1 99.405,79.17
X$15048 348 59 349 644 645 cell_1rw
* cell instance $15049 r0 *1 100.11,79.17
X$15049 350 59 351 644 645 cell_1rw
* cell instance $15050 r0 *1 100.815,79.17
X$15050 352 59 353 644 645 cell_1rw
* cell instance $15051 r0 *1 101.52,79.17
X$15051 354 59 355 644 645 cell_1rw
* cell instance $15052 r0 *1 102.225,79.17
X$15052 356 59 357 644 645 cell_1rw
* cell instance $15053 r0 *1 102.93,79.17
X$15053 358 59 359 644 645 cell_1rw
* cell instance $15054 r0 *1 103.635,79.17
X$15054 360 59 361 644 645 cell_1rw
* cell instance $15055 r0 *1 104.34,79.17
X$15055 362 59 363 644 645 cell_1rw
* cell instance $15056 r0 *1 105.045,79.17
X$15056 364 59 365 644 645 cell_1rw
* cell instance $15057 r0 *1 105.75,79.17
X$15057 366 59 367 644 645 cell_1rw
* cell instance $15058 r0 *1 106.455,79.17
X$15058 368 59 369 644 645 cell_1rw
* cell instance $15059 r0 *1 107.16,79.17
X$15059 370 59 371 644 645 cell_1rw
* cell instance $15060 r0 *1 107.865,79.17
X$15060 372 59 373 644 645 cell_1rw
* cell instance $15061 r0 *1 108.57,79.17
X$15061 374 59 375 644 645 cell_1rw
* cell instance $15062 r0 *1 109.275,79.17
X$15062 376 59 377 644 645 cell_1rw
* cell instance $15063 r0 *1 109.98,79.17
X$15063 378 59 379 644 645 cell_1rw
* cell instance $15064 r0 *1 110.685,79.17
X$15064 380 59 381 644 645 cell_1rw
* cell instance $15065 r0 *1 111.39,79.17
X$15065 382 59 383 644 645 cell_1rw
* cell instance $15066 r0 *1 112.095,79.17
X$15066 384 59 385 644 645 cell_1rw
* cell instance $15067 r0 *1 112.8,79.17
X$15067 386 59 387 644 645 cell_1rw
* cell instance $15068 r0 *1 113.505,79.17
X$15068 388 59 389 644 645 cell_1rw
* cell instance $15069 r0 *1 114.21,79.17
X$15069 390 59 391 644 645 cell_1rw
* cell instance $15070 r0 *1 114.915,79.17
X$15070 392 59 393 644 645 cell_1rw
* cell instance $15071 r0 *1 115.62,79.17
X$15071 394 59 395 644 645 cell_1rw
* cell instance $15072 r0 *1 116.325,79.17
X$15072 396 59 397 644 645 cell_1rw
* cell instance $15073 r0 *1 117.03,79.17
X$15073 398 59 399 644 645 cell_1rw
* cell instance $15074 r0 *1 117.735,79.17
X$15074 400 59 401 644 645 cell_1rw
* cell instance $15075 r0 *1 118.44,79.17
X$15075 402 59 403 644 645 cell_1rw
* cell instance $15076 r0 *1 119.145,79.17
X$15076 404 59 405 644 645 cell_1rw
* cell instance $15077 r0 *1 119.85,79.17
X$15077 406 59 407 644 645 cell_1rw
* cell instance $15078 r0 *1 120.555,79.17
X$15078 408 59 409 644 645 cell_1rw
* cell instance $15079 r0 *1 121.26,79.17
X$15079 410 59 411 644 645 cell_1rw
* cell instance $15080 r0 *1 121.965,79.17
X$15080 412 59 413 644 645 cell_1rw
* cell instance $15081 r0 *1 122.67,79.17
X$15081 414 59 415 644 645 cell_1rw
* cell instance $15082 r0 *1 123.375,79.17
X$15082 416 59 417 644 645 cell_1rw
* cell instance $15083 r0 *1 124.08,79.17
X$15083 418 59 419 644 645 cell_1rw
* cell instance $15084 r0 *1 124.785,79.17
X$15084 420 59 421 644 645 cell_1rw
* cell instance $15085 r0 *1 125.49,79.17
X$15085 422 59 423 644 645 cell_1rw
* cell instance $15086 r0 *1 126.195,79.17
X$15086 424 59 425 644 645 cell_1rw
* cell instance $15087 r0 *1 126.9,79.17
X$15087 426 59 427 644 645 cell_1rw
* cell instance $15088 r0 *1 127.605,79.17
X$15088 428 59 429 644 645 cell_1rw
* cell instance $15089 r0 *1 128.31,79.17
X$15089 430 59 431 644 645 cell_1rw
* cell instance $15090 r0 *1 129.015,79.17
X$15090 432 59 433 644 645 cell_1rw
* cell instance $15091 r0 *1 129.72,79.17
X$15091 434 59 435 644 645 cell_1rw
* cell instance $15092 r0 *1 130.425,79.17
X$15092 436 59 437 644 645 cell_1rw
* cell instance $15093 r0 *1 131.13,79.17
X$15093 438 59 439 644 645 cell_1rw
* cell instance $15094 r0 *1 131.835,79.17
X$15094 440 59 441 644 645 cell_1rw
* cell instance $15095 r0 *1 132.54,79.17
X$15095 442 59 443 644 645 cell_1rw
* cell instance $15096 r0 *1 133.245,79.17
X$15096 444 59 445 644 645 cell_1rw
* cell instance $15097 r0 *1 133.95,79.17
X$15097 446 59 447 644 645 cell_1rw
* cell instance $15098 r0 *1 134.655,79.17
X$15098 448 59 449 644 645 cell_1rw
* cell instance $15099 r0 *1 135.36,79.17
X$15099 450 59 451 644 645 cell_1rw
* cell instance $15100 r0 *1 136.065,79.17
X$15100 452 59 453 644 645 cell_1rw
* cell instance $15101 r0 *1 136.77,79.17
X$15101 454 59 455 644 645 cell_1rw
* cell instance $15102 r0 *1 137.475,79.17
X$15102 456 59 457 644 645 cell_1rw
* cell instance $15103 r0 *1 138.18,79.17
X$15103 458 59 459 644 645 cell_1rw
* cell instance $15104 r0 *1 138.885,79.17
X$15104 460 59 461 644 645 cell_1rw
* cell instance $15105 r0 *1 139.59,79.17
X$15105 462 59 463 644 645 cell_1rw
* cell instance $15106 r0 *1 140.295,79.17
X$15106 464 59 465 644 645 cell_1rw
* cell instance $15107 r0 *1 141,79.17
X$15107 466 59 467 644 645 cell_1rw
* cell instance $15108 r0 *1 141.705,79.17
X$15108 468 59 469 644 645 cell_1rw
* cell instance $15109 r0 *1 142.41,79.17
X$15109 470 59 471 644 645 cell_1rw
* cell instance $15110 r0 *1 143.115,79.17
X$15110 472 59 473 644 645 cell_1rw
* cell instance $15111 r0 *1 143.82,79.17
X$15111 474 59 475 644 645 cell_1rw
* cell instance $15112 r0 *1 144.525,79.17
X$15112 476 59 477 644 645 cell_1rw
* cell instance $15113 r0 *1 145.23,79.17
X$15113 478 59 479 644 645 cell_1rw
* cell instance $15114 r0 *1 145.935,79.17
X$15114 480 59 481 644 645 cell_1rw
* cell instance $15115 r0 *1 146.64,79.17
X$15115 482 59 483 644 645 cell_1rw
* cell instance $15116 r0 *1 147.345,79.17
X$15116 484 59 485 644 645 cell_1rw
* cell instance $15117 r0 *1 148.05,79.17
X$15117 486 59 487 644 645 cell_1rw
* cell instance $15118 r0 *1 148.755,79.17
X$15118 488 59 489 644 645 cell_1rw
* cell instance $15119 r0 *1 149.46,79.17
X$15119 490 59 491 644 645 cell_1rw
* cell instance $15120 r0 *1 150.165,79.17
X$15120 492 59 493 644 645 cell_1rw
* cell instance $15121 r0 *1 150.87,79.17
X$15121 494 59 495 644 645 cell_1rw
* cell instance $15122 r0 *1 151.575,79.17
X$15122 496 59 497 644 645 cell_1rw
* cell instance $15123 r0 *1 152.28,79.17
X$15123 498 59 499 644 645 cell_1rw
* cell instance $15124 r0 *1 152.985,79.17
X$15124 500 59 501 644 645 cell_1rw
* cell instance $15125 r0 *1 153.69,79.17
X$15125 502 59 503 644 645 cell_1rw
* cell instance $15126 r0 *1 154.395,79.17
X$15126 504 59 505 644 645 cell_1rw
* cell instance $15127 r0 *1 155.1,79.17
X$15127 506 59 507 644 645 cell_1rw
* cell instance $15128 r0 *1 155.805,79.17
X$15128 508 59 509 644 645 cell_1rw
* cell instance $15129 r0 *1 156.51,79.17
X$15129 510 59 511 644 645 cell_1rw
* cell instance $15130 r0 *1 157.215,79.17
X$15130 512 59 513 644 645 cell_1rw
* cell instance $15131 r0 *1 157.92,79.17
X$15131 514 59 515 644 645 cell_1rw
* cell instance $15132 r0 *1 158.625,79.17
X$15132 516 59 517 644 645 cell_1rw
* cell instance $15133 r0 *1 159.33,79.17
X$15133 518 59 519 644 645 cell_1rw
* cell instance $15134 r0 *1 160.035,79.17
X$15134 520 59 521 644 645 cell_1rw
* cell instance $15135 r0 *1 160.74,79.17
X$15135 522 59 523 644 645 cell_1rw
* cell instance $15136 r0 *1 161.445,79.17
X$15136 524 59 525 644 645 cell_1rw
* cell instance $15137 r0 *1 162.15,79.17
X$15137 526 59 527 644 645 cell_1rw
* cell instance $15138 r0 *1 162.855,79.17
X$15138 528 59 529 644 645 cell_1rw
* cell instance $15139 r0 *1 163.56,79.17
X$15139 530 59 531 644 645 cell_1rw
* cell instance $15140 r0 *1 164.265,79.17
X$15140 532 59 533 644 645 cell_1rw
* cell instance $15141 r0 *1 164.97,79.17
X$15141 534 59 535 644 645 cell_1rw
* cell instance $15142 r0 *1 165.675,79.17
X$15142 536 59 537 644 645 cell_1rw
* cell instance $15143 r0 *1 166.38,79.17
X$15143 538 59 539 644 645 cell_1rw
* cell instance $15144 r0 *1 167.085,79.17
X$15144 540 59 541 644 645 cell_1rw
* cell instance $15145 r0 *1 167.79,79.17
X$15145 542 59 543 644 645 cell_1rw
* cell instance $15146 r0 *1 168.495,79.17
X$15146 544 59 545 644 645 cell_1rw
* cell instance $15147 r0 *1 169.2,79.17
X$15147 546 59 547 644 645 cell_1rw
* cell instance $15148 r0 *1 169.905,79.17
X$15148 548 59 549 644 645 cell_1rw
* cell instance $15149 r0 *1 170.61,79.17
X$15149 550 59 551 644 645 cell_1rw
* cell instance $15150 r0 *1 171.315,79.17
X$15150 552 59 553 644 645 cell_1rw
* cell instance $15151 r0 *1 172.02,79.17
X$15151 554 59 555 644 645 cell_1rw
* cell instance $15152 r0 *1 172.725,79.17
X$15152 556 59 557 644 645 cell_1rw
* cell instance $15153 r0 *1 173.43,79.17
X$15153 558 59 559 644 645 cell_1rw
* cell instance $15154 r0 *1 174.135,79.17
X$15154 560 59 561 644 645 cell_1rw
* cell instance $15155 r0 *1 174.84,79.17
X$15155 562 59 563 644 645 cell_1rw
* cell instance $15156 r0 *1 175.545,79.17
X$15156 564 59 565 644 645 cell_1rw
* cell instance $15157 r0 *1 176.25,79.17
X$15157 566 59 567 644 645 cell_1rw
* cell instance $15158 r0 *1 176.955,79.17
X$15158 568 59 569 644 645 cell_1rw
* cell instance $15159 r0 *1 177.66,79.17
X$15159 570 59 571 644 645 cell_1rw
* cell instance $15160 r0 *1 178.365,79.17
X$15160 572 59 573 644 645 cell_1rw
* cell instance $15161 r0 *1 179.07,79.17
X$15161 574 59 575 644 645 cell_1rw
* cell instance $15162 r0 *1 179.775,79.17
X$15162 576 59 577 644 645 cell_1rw
* cell instance $15163 r0 *1 180.48,79.17
X$15163 578 59 579 644 645 cell_1rw
* cell instance $15164 m0 *1 0.705,81.9
X$15164 67 60 68 644 645 cell_1rw
* cell instance $15165 m0 *1 0,81.9
X$15165 65 60 66 644 645 cell_1rw
* cell instance $15166 m0 *1 1.41,81.9
X$15166 69 60 70 644 645 cell_1rw
* cell instance $15167 m0 *1 2.115,81.9
X$15167 71 60 72 644 645 cell_1rw
* cell instance $15168 m0 *1 2.82,81.9
X$15168 73 60 74 644 645 cell_1rw
* cell instance $15169 m0 *1 3.525,81.9
X$15169 75 60 76 644 645 cell_1rw
* cell instance $15170 m0 *1 4.23,81.9
X$15170 77 60 78 644 645 cell_1rw
* cell instance $15171 m0 *1 4.935,81.9
X$15171 79 60 80 644 645 cell_1rw
* cell instance $15172 m0 *1 5.64,81.9
X$15172 81 60 82 644 645 cell_1rw
* cell instance $15173 m0 *1 6.345,81.9
X$15173 83 60 84 644 645 cell_1rw
* cell instance $15174 m0 *1 7.05,81.9
X$15174 85 60 86 644 645 cell_1rw
* cell instance $15175 m0 *1 7.755,81.9
X$15175 87 60 88 644 645 cell_1rw
* cell instance $15176 m0 *1 8.46,81.9
X$15176 89 60 90 644 645 cell_1rw
* cell instance $15177 m0 *1 9.165,81.9
X$15177 91 60 92 644 645 cell_1rw
* cell instance $15178 m0 *1 9.87,81.9
X$15178 93 60 94 644 645 cell_1rw
* cell instance $15179 m0 *1 10.575,81.9
X$15179 95 60 96 644 645 cell_1rw
* cell instance $15180 m0 *1 11.28,81.9
X$15180 97 60 98 644 645 cell_1rw
* cell instance $15181 m0 *1 11.985,81.9
X$15181 99 60 100 644 645 cell_1rw
* cell instance $15182 m0 *1 12.69,81.9
X$15182 101 60 102 644 645 cell_1rw
* cell instance $15183 m0 *1 13.395,81.9
X$15183 103 60 104 644 645 cell_1rw
* cell instance $15184 m0 *1 14.1,81.9
X$15184 105 60 106 644 645 cell_1rw
* cell instance $15185 m0 *1 14.805,81.9
X$15185 107 60 108 644 645 cell_1rw
* cell instance $15186 m0 *1 15.51,81.9
X$15186 109 60 110 644 645 cell_1rw
* cell instance $15187 m0 *1 16.215,81.9
X$15187 111 60 112 644 645 cell_1rw
* cell instance $15188 m0 *1 16.92,81.9
X$15188 113 60 114 644 645 cell_1rw
* cell instance $15189 m0 *1 17.625,81.9
X$15189 115 60 116 644 645 cell_1rw
* cell instance $15190 m0 *1 18.33,81.9
X$15190 117 60 118 644 645 cell_1rw
* cell instance $15191 m0 *1 19.035,81.9
X$15191 119 60 120 644 645 cell_1rw
* cell instance $15192 m0 *1 19.74,81.9
X$15192 121 60 122 644 645 cell_1rw
* cell instance $15193 m0 *1 20.445,81.9
X$15193 123 60 124 644 645 cell_1rw
* cell instance $15194 m0 *1 21.15,81.9
X$15194 125 60 126 644 645 cell_1rw
* cell instance $15195 m0 *1 21.855,81.9
X$15195 127 60 128 644 645 cell_1rw
* cell instance $15196 m0 *1 22.56,81.9
X$15196 129 60 130 644 645 cell_1rw
* cell instance $15197 m0 *1 23.265,81.9
X$15197 131 60 132 644 645 cell_1rw
* cell instance $15198 m0 *1 23.97,81.9
X$15198 133 60 134 644 645 cell_1rw
* cell instance $15199 m0 *1 24.675,81.9
X$15199 135 60 136 644 645 cell_1rw
* cell instance $15200 m0 *1 25.38,81.9
X$15200 137 60 138 644 645 cell_1rw
* cell instance $15201 m0 *1 26.085,81.9
X$15201 139 60 140 644 645 cell_1rw
* cell instance $15202 m0 *1 26.79,81.9
X$15202 141 60 142 644 645 cell_1rw
* cell instance $15203 m0 *1 27.495,81.9
X$15203 143 60 144 644 645 cell_1rw
* cell instance $15204 m0 *1 28.2,81.9
X$15204 145 60 146 644 645 cell_1rw
* cell instance $15205 m0 *1 28.905,81.9
X$15205 147 60 148 644 645 cell_1rw
* cell instance $15206 m0 *1 29.61,81.9
X$15206 149 60 150 644 645 cell_1rw
* cell instance $15207 m0 *1 30.315,81.9
X$15207 151 60 152 644 645 cell_1rw
* cell instance $15208 m0 *1 31.02,81.9
X$15208 153 60 154 644 645 cell_1rw
* cell instance $15209 m0 *1 31.725,81.9
X$15209 155 60 156 644 645 cell_1rw
* cell instance $15210 m0 *1 32.43,81.9
X$15210 157 60 158 644 645 cell_1rw
* cell instance $15211 m0 *1 33.135,81.9
X$15211 159 60 160 644 645 cell_1rw
* cell instance $15212 m0 *1 33.84,81.9
X$15212 161 60 162 644 645 cell_1rw
* cell instance $15213 m0 *1 34.545,81.9
X$15213 163 60 164 644 645 cell_1rw
* cell instance $15214 m0 *1 35.25,81.9
X$15214 165 60 166 644 645 cell_1rw
* cell instance $15215 m0 *1 35.955,81.9
X$15215 167 60 168 644 645 cell_1rw
* cell instance $15216 m0 *1 36.66,81.9
X$15216 169 60 170 644 645 cell_1rw
* cell instance $15217 m0 *1 37.365,81.9
X$15217 171 60 172 644 645 cell_1rw
* cell instance $15218 m0 *1 38.07,81.9
X$15218 173 60 174 644 645 cell_1rw
* cell instance $15219 m0 *1 38.775,81.9
X$15219 175 60 176 644 645 cell_1rw
* cell instance $15220 m0 *1 39.48,81.9
X$15220 177 60 178 644 645 cell_1rw
* cell instance $15221 m0 *1 40.185,81.9
X$15221 179 60 180 644 645 cell_1rw
* cell instance $15222 m0 *1 40.89,81.9
X$15222 181 60 182 644 645 cell_1rw
* cell instance $15223 m0 *1 41.595,81.9
X$15223 183 60 184 644 645 cell_1rw
* cell instance $15224 m0 *1 42.3,81.9
X$15224 185 60 186 644 645 cell_1rw
* cell instance $15225 m0 *1 43.005,81.9
X$15225 187 60 188 644 645 cell_1rw
* cell instance $15226 m0 *1 43.71,81.9
X$15226 189 60 190 644 645 cell_1rw
* cell instance $15227 m0 *1 44.415,81.9
X$15227 191 60 192 644 645 cell_1rw
* cell instance $15228 m0 *1 45.12,81.9
X$15228 193 60 194 644 645 cell_1rw
* cell instance $15229 m0 *1 45.825,81.9
X$15229 195 60 196 644 645 cell_1rw
* cell instance $15230 m0 *1 46.53,81.9
X$15230 197 60 198 644 645 cell_1rw
* cell instance $15231 m0 *1 47.235,81.9
X$15231 199 60 200 644 645 cell_1rw
* cell instance $15232 m0 *1 47.94,81.9
X$15232 201 60 202 644 645 cell_1rw
* cell instance $15233 m0 *1 48.645,81.9
X$15233 203 60 204 644 645 cell_1rw
* cell instance $15234 m0 *1 49.35,81.9
X$15234 205 60 206 644 645 cell_1rw
* cell instance $15235 m0 *1 50.055,81.9
X$15235 207 60 208 644 645 cell_1rw
* cell instance $15236 m0 *1 50.76,81.9
X$15236 209 60 210 644 645 cell_1rw
* cell instance $15237 m0 *1 51.465,81.9
X$15237 211 60 212 644 645 cell_1rw
* cell instance $15238 m0 *1 52.17,81.9
X$15238 213 60 214 644 645 cell_1rw
* cell instance $15239 m0 *1 52.875,81.9
X$15239 215 60 216 644 645 cell_1rw
* cell instance $15240 m0 *1 53.58,81.9
X$15240 217 60 218 644 645 cell_1rw
* cell instance $15241 m0 *1 54.285,81.9
X$15241 219 60 220 644 645 cell_1rw
* cell instance $15242 m0 *1 54.99,81.9
X$15242 221 60 222 644 645 cell_1rw
* cell instance $15243 m0 *1 55.695,81.9
X$15243 223 60 224 644 645 cell_1rw
* cell instance $15244 m0 *1 56.4,81.9
X$15244 225 60 226 644 645 cell_1rw
* cell instance $15245 m0 *1 57.105,81.9
X$15245 227 60 228 644 645 cell_1rw
* cell instance $15246 m0 *1 57.81,81.9
X$15246 229 60 230 644 645 cell_1rw
* cell instance $15247 m0 *1 58.515,81.9
X$15247 231 60 232 644 645 cell_1rw
* cell instance $15248 m0 *1 59.22,81.9
X$15248 233 60 234 644 645 cell_1rw
* cell instance $15249 m0 *1 59.925,81.9
X$15249 235 60 236 644 645 cell_1rw
* cell instance $15250 m0 *1 60.63,81.9
X$15250 237 60 238 644 645 cell_1rw
* cell instance $15251 m0 *1 61.335,81.9
X$15251 239 60 240 644 645 cell_1rw
* cell instance $15252 m0 *1 62.04,81.9
X$15252 241 60 242 644 645 cell_1rw
* cell instance $15253 m0 *1 62.745,81.9
X$15253 243 60 244 644 645 cell_1rw
* cell instance $15254 m0 *1 63.45,81.9
X$15254 245 60 246 644 645 cell_1rw
* cell instance $15255 m0 *1 64.155,81.9
X$15255 247 60 248 644 645 cell_1rw
* cell instance $15256 m0 *1 64.86,81.9
X$15256 249 60 250 644 645 cell_1rw
* cell instance $15257 m0 *1 65.565,81.9
X$15257 251 60 252 644 645 cell_1rw
* cell instance $15258 m0 *1 66.27,81.9
X$15258 253 60 254 644 645 cell_1rw
* cell instance $15259 m0 *1 66.975,81.9
X$15259 255 60 256 644 645 cell_1rw
* cell instance $15260 m0 *1 67.68,81.9
X$15260 257 60 258 644 645 cell_1rw
* cell instance $15261 m0 *1 68.385,81.9
X$15261 259 60 260 644 645 cell_1rw
* cell instance $15262 m0 *1 69.09,81.9
X$15262 261 60 262 644 645 cell_1rw
* cell instance $15263 m0 *1 69.795,81.9
X$15263 263 60 264 644 645 cell_1rw
* cell instance $15264 m0 *1 70.5,81.9
X$15264 265 60 266 644 645 cell_1rw
* cell instance $15265 m0 *1 71.205,81.9
X$15265 267 60 268 644 645 cell_1rw
* cell instance $15266 m0 *1 71.91,81.9
X$15266 269 60 270 644 645 cell_1rw
* cell instance $15267 m0 *1 72.615,81.9
X$15267 271 60 272 644 645 cell_1rw
* cell instance $15268 m0 *1 73.32,81.9
X$15268 273 60 274 644 645 cell_1rw
* cell instance $15269 m0 *1 74.025,81.9
X$15269 275 60 276 644 645 cell_1rw
* cell instance $15270 m0 *1 74.73,81.9
X$15270 277 60 278 644 645 cell_1rw
* cell instance $15271 m0 *1 75.435,81.9
X$15271 279 60 280 644 645 cell_1rw
* cell instance $15272 m0 *1 76.14,81.9
X$15272 281 60 282 644 645 cell_1rw
* cell instance $15273 m0 *1 76.845,81.9
X$15273 283 60 284 644 645 cell_1rw
* cell instance $15274 m0 *1 77.55,81.9
X$15274 285 60 286 644 645 cell_1rw
* cell instance $15275 m0 *1 78.255,81.9
X$15275 287 60 288 644 645 cell_1rw
* cell instance $15276 m0 *1 78.96,81.9
X$15276 289 60 290 644 645 cell_1rw
* cell instance $15277 m0 *1 79.665,81.9
X$15277 291 60 292 644 645 cell_1rw
* cell instance $15278 m0 *1 80.37,81.9
X$15278 293 60 294 644 645 cell_1rw
* cell instance $15279 m0 *1 81.075,81.9
X$15279 295 60 296 644 645 cell_1rw
* cell instance $15280 m0 *1 81.78,81.9
X$15280 297 60 298 644 645 cell_1rw
* cell instance $15281 m0 *1 82.485,81.9
X$15281 299 60 300 644 645 cell_1rw
* cell instance $15282 m0 *1 83.19,81.9
X$15282 301 60 302 644 645 cell_1rw
* cell instance $15283 m0 *1 83.895,81.9
X$15283 303 60 304 644 645 cell_1rw
* cell instance $15284 m0 *1 84.6,81.9
X$15284 305 60 306 644 645 cell_1rw
* cell instance $15285 m0 *1 85.305,81.9
X$15285 307 60 308 644 645 cell_1rw
* cell instance $15286 m0 *1 86.01,81.9
X$15286 309 60 310 644 645 cell_1rw
* cell instance $15287 m0 *1 86.715,81.9
X$15287 311 60 312 644 645 cell_1rw
* cell instance $15288 m0 *1 87.42,81.9
X$15288 313 60 314 644 645 cell_1rw
* cell instance $15289 m0 *1 88.125,81.9
X$15289 315 60 316 644 645 cell_1rw
* cell instance $15290 m0 *1 88.83,81.9
X$15290 317 60 318 644 645 cell_1rw
* cell instance $15291 m0 *1 89.535,81.9
X$15291 319 60 320 644 645 cell_1rw
* cell instance $15292 m0 *1 90.24,81.9
X$15292 321 60 323 644 645 cell_1rw
* cell instance $15293 m0 *1 90.945,81.9
X$15293 324 60 325 644 645 cell_1rw
* cell instance $15294 m0 *1 91.65,81.9
X$15294 326 60 327 644 645 cell_1rw
* cell instance $15295 m0 *1 92.355,81.9
X$15295 328 60 329 644 645 cell_1rw
* cell instance $15296 m0 *1 93.06,81.9
X$15296 330 60 331 644 645 cell_1rw
* cell instance $15297 m0 *1 93.765,81.9
X$15297 332 60 333 644 645 cell_1rw
* cell instance $15298 m0 *1 94.47,81.9
X$15298 334 60 335 644 645 cell_1rw
* cell instance $15299 m0 *1 95.175,81.9
X$15299 336 60 337 644 645 cell_1rw
* cell instance $15300 m0 *1 95.88,81.9
X$15300 338 60 339 644 645 cell_1rw
* cell instance $15301 m0 *1 96.585,81.9
X$15301 340 60 341 644 645 cell_1rw
* cell instance $15302 m0 *1 97.29,81.9
X$15302 342 60 343 644 645 cell_1rw
* cell instance $15303 m0 *1 97.995,81.9
X$15303 344 60 345 644 645 cell_1rw
* cell instance $15304 m0 *1 98.7,81.9
X$15304 346 60 347 644 645 cell_1rw
* cell instance $15305 m0 *1 99.405,81.9
X$15305 348 60 349 644 645 cell_1rw
* cell instance $15306 m0 *1 100.11,81.9
X$15306 350 60 351 644 645 cell_1rw
* cell instance $15307 m0 *1 100.815,81.9
X$15307 352 60 353 644 645 cell_1rw
* cell instance $15308 m0 *1 101.52,81.9
X$15308 354 60 355 644 645 cell_1rw
* cell instance $15309 m0 *1 102.225,81.9
X$15309 356 60 357 644 645 cell_1rw
* cell instance $15310 m0 *1 102.93,81.9
X$15310 358 60 359 644 645 cell_1rw
* cell instance $15311 m0 *1 103.635,81.9
X$15311 360 60 361 644 645 cell_1rw
* cell instance $15312 m0 *1 104.34,81.9
X$15312 362 60 363 644 645 cell_1rw
* cell instance $15313 m0 *1 105.045,81.9
X$15313 364 60 365 644 645 cell_1rw
* cell instance $15314 m0 *1 105.75,81.9
X$15314 366 60 367 644 645 cell_1rw
* cell instance $15315 m0 *1 106.455,81.9
X$15315 368 60 369 644 645 cell_1rw
* cell instance $15316 m0 *1 107.16,81.9
X$15316 370 60 371 644 645 cell_1rw
* cell instance $15317 m0 *1 107.865,81.9
X$15317 372 60 373 644 645 cell_1rw
* cell instance $15318 m0 *1 108.57,81.9
X$15318 374 60 375 644 645 cell_1rw
* cell instance $15319 m0 *1 109.275,81.9
X$15319 376 60 377 644 645 cell_1rw
* cell instance $15320 m0 *1 109.98,81.9
X$15320 378 60 379 644 645 cell_1rw
* cell instance $15321 m0 *1 110.685,81.9
X$15321 380 60 381 644 645 cell_1rw
* cell instance $15322 m0 *1 111.39,81.9
X$15322 382 60 383 644 645 cell_1rw
* cell instance $15323 m0 *1 112.095,81.9
X$15323 384 60 385 644 645 cell_1rw
* cell instance $15324 m0 *1 112.8,81.9
X$15324 386 60 387 644 645 cell_1rw
* cell instance $15325 m0 *1 113.505,81.9
X$15325 388 60 389 644 645 cell_1rw
* cell instance $15326 m0 *1 114.21,81.9
X$15326 390 60 391 644 645 cell_1rw
* cell instance $15327 m0 *1 114.915,81.9
X$15327 392 60 393 644 645 cell_1rw
* cell instance $15328 m0 *1 115.62,81.9
X$15328 394 60 395 644 645 cell_1rw
* cell instance $15329 m0 *1 116.325,81.9
X$15329 396 60 397 644 645 cell_1rw
* cell instance $15330 m0 *1 117.03,81.9
X$15330 398 60 399 644 645 cell_1rw
* cell instance $15331 m0 *1 117.735,81.9
X$15331 400 60 401 644 645 cell_1rw
* cell instance $15332 m0 *1 118.44,81.9
X$15332 402 60 403 644 645 cell_1rw
* cell instance $15333 m0 *1 119.145,81.9
X$15333 404 60 405 644 645 cell_1rw
* cell instance $15334 m0 *1 119.85,81.9
X$15334 406 60 407 644 645 cell_1rw
* cell instance $15335 m0 *1 120.555,81.9
X$15335 408 60 409 644 645 cell_1rw
* cell instance $15336 m0 *1 121.26,81.9
X$15336 410 60 411 644 645 cell_1rw
* cell instance $15337 m0 *1 121.965,81.9
X$15337 412 60 413 644 645 cell_1rw
* cell instance $15338 m0 *1 122.67,81.9
X$15338 414 60 415 644 645 cell_1rw
* cell instance $15339 m0 *1 123.375,81.9
X$15339 416 60 417 644 645 cell_1rw
* cell instance $15340 m0 *1 124.08,81.9
X$15340 418 60 419 644 645 cell_1rw
* cell instance $15341 m0 *1 124.785,81.9
X$15341 420 60 421 644 645 cell_1rw
* cell instance $15342 m0 *1 125.49,81.9
X$15342 422 60 423 644 645 cell_1rw
* cell instance $15343 m0 *1 126.195,81.9
X$15343 424 60 425 644 645 cell_1rw
* cell instance $15344 m0 *1 126.9,81.9
X$15344 426 60 427 644 645 cell_1rw
* cell instance $15345 m0 *1 127.605,81.9
X$15345 428 60 429 644 645 cell_1rw
* cell instance $15346 m0 *1 128.31,81.9
X$15346 430 60 431 644 645 cell_1rw
* cell instance $15347 m0 *1 129.015,81.9
X$15347 432 60 433 644 645 cell_1rw
* cell instance $15348 m0 *1 129.72,81.9
X$15348 434 60 435 644 645 cell_1rw
* cell instance $15349 m0 *1 130.425,81.9
X$15349 436 60 437 644 645 cell_1rw
* cell instance $15350 m0 *1 131.13,81.9
X$15350 438 60 439 644 645 cell_1rw
* cell instance $15351 m0 *1 131.835,81.9
X$15351 440 60 441 644 645 cell_1rw
* cell instance $15352 m0 *1 132.54,81.9
X$15352 442 60 443 644 645 cell_1rw
* cell instance $15353 m0 *1 133.245,81.9
X$15353 444 60 445 644 645 cell_1rw
* cell instance $15354 m0 *1 133.95,81.9
X$15354 446 60 447 644 645 cell_1rw
* cell instance $15355 m0 *1 134.655,81.9
X$15355 448 60 449 644 645 cell_1rw
* cell instance $15356 m0 *1 135.36,81.9
X$15356 450 60 451 644 645 cell_1rw
* cell instance $15357 m0 *1 136.065,81.9
X$15357 452 60 453 644 645 cell_1rw
* cell instance $15358 m0 *1 136.77,81.9
X$15358 454 60 455 644 645 cell_1rw
* cell instance $15359 m0 *1 137.475,81.9
X$15359 456 60 457 644 645 cell_1rw
* cell instance $15360 m0 *1 138.18,81.9
X$15360 458 60 459 644 645 cell_1rw
* cell instance $15361 m0 *1 138.885,81.9
X$15361 460 60 461 644 645 cell_1rw
* cell instance $15362 m0 *1 139.59,81.9
X$15362 462 60 463 644 645 cell_1rw
* cell instance $15363 m0 *1 140.295,81.9
X$15363 464 60 465 644 645 cell_1rw
* cell instance $15364 m0 *1 141,81.9
X$15364 466 60 467 644 645 cell_1rw
* cell instance $15365 m0 *1 141.705,81.9
X$15365 468 60 469 644 645 cell_1rw
* cell instance $15366 m0 *1 142.41,81.9
X$15366 470 60 471 644 645 cell_1rw
* cell instance $15367 m0 *1 143.115,81.9
X$15367 472 60 473 644 645 cell_1rw
* cell instance $15368 m0 *1 143.82,81.9
X$15368 474 60 475 644 645 cell_1rw
* cell instance $15369 m0 *1 144.525,81.9
X$15369 476 60 477 644 645 cell_1rw
* cell instance $15370 m0 *1 145.23,81.9
X$15370 478 60 479 644 645 cell_1rw
* cell instance $15371 m0 *1 145.935,81.9
X$15371 480 60 481 644 645 cell_1rw
* cell instance $15372 m0 *1 146.64,81.9
X$15372 482 60 483 644 645 cell_1rw
* cell instance $15373 m0 *1 147.345,81.9
X$15373 484 60 485 644 645 cell_1rw
* cell instance $15374 m0 *1 148.05,81.9
X$15374 486 60 487 644 645 cell_1rw
* cell instance $15375 m0 *1 148.755,81.9
X$15375 488 60 489 644 645 cell_1rw
* cell instance $15376 m0 *1 149.46,81.9
X$15376 490 60 491 644 645 cell_1rw
* cell instance $15377 m0 *1 150.165,81.9
X$15377 492 60 493 644 645 cell_1rw
* cell instance $15378 m0 *1 150.87,81.9
X$15378 494 60 495 644 645 cell_1rw
* cell instance $15379 m0 *1 151.575,81.9
X$15379 496 60 497 644 645 cell_1rw
* cell instance $15380 m0 *1 152.28,81.9
X$15380 498 60 499 644 645 cell_1rw
* cell instance $15381 m0 *1 152.985,81.9
X$15381 500 60 501 644 645 cell_1rw
* cell instance $15382 m0 *1 153.69,81.9
X$15382 502 60 503 644 645 cell_1rw
* cell instance $15383 m0 *1 154.395,81.9
X$15383 504 60 505 644 645 cell_1rw
* cell instance $15384 m0 *1 155.1,81.9
X$15384 506 60 507 644 645 cell_1rw
* cell instance $15385 m0 *1 155.805,81.9
X$15385 508 60 509 644 645 cell_1rw
* cell instance $15386 m0 *1 156.51,81.9
X$15386 510 60 511 644 645 cell_1rw
* cell instance $15387 m0 *1 157.215,81.9
X$15387 512 60 513 644 645 cell_1rw
* cell instance $15388 m0 *1 157.92,81.9
X$15388 514 60 515 644 645 cell_1rw
* cell instance $15389 m0 *1 158.625,81.9
X$15389 516 60 517 644 645 cell_1rw
* cell instance $15390 m0 *1 159.33,81.9
X$15390 518 60 519 644 645 cell_1rw
* cell instance $15391 m0 *1 160.035,81.9
X$15391 520 60 521 644 645 cell_1rw
* cell instance $15392 m0 *1 160.74,81.9
X$15392 522 60 523 644 645 cell_1rw
* cell instance $15393 m0 *1 161.445,81.9
X$15393 524 60 525 644 645 cell_1rw
* cell instance $15394 m0 *1 162.15,81.9
X$15394 526 60 527 644 645 cell_1rw
* cell instance $15395 m0 *1 162.855,81.9
X$15395 528 60 529 644 645 cell_1rw
* cell instance $15396 m0 *1 163.56,81.9
X$15396 530 60 531 644 645 cell_1rw
* cell instance $15397 m0 *1 164.265,81.9
X$15397 532 60 533 644 645 cell_1rw
* cell instance $15398 m0 *1 164.97,81.9
X$15398 534 60 535 644 645 cell_1rw
* cell instance $15399 m0 *1 165.675,81.9
X$15399 536 60 537 644 645 cell_1rw
* cell instance $15400 m0 *1 166.38,81.9
X$15400 538 60 539 644 645 cell_1rw
* cell instance $15401 m0 *1 167.085,81.9
X$15401 540 60 541 644 645 cell_1rw
* cell instance $15402 m0 *1 167.79,81.9
X$15402 542 60 543 644 645 cell_1rw
* cell instance $15403 m0 *1 168.495,81.9
X$15403 544 60 545 644 645 cell_1rw
* cell instance $15404 m0 *1 169.2,81.9
X$15404 546 60 547 644 645 cell_1rw
* cell instance $15405 m0 *1 169.905,81.9
X$15405 548 60 549 644 645 cell_1rw
* cell instance $15406 m0 *1 170.61,81.9
X$15406 550 60 551 644 645 cell_1rw
* cell instance $15407 m0 *1 171.315,81.9
X$15407 552 60 553 644 645 cell_1rw
* cell instance $15408 m0 *1 172.02,81.9
X$15408 554 60 555 644 645 cell_1rw
* cell instance $15409 m0 *1 172.725,81.9
X$15409 556 60 557 644 645 cell_1rw
* cell instance $15410 m0 *1 173.43,81.9
X$15410 558 60 559 644 645 cell_1rw
* cell instance $15411 m0 *1 174.135,81.9
X$15411 560 60 561 644 645 cell_1rw
* cell instance $15412 m0 *1 174.84,81.9
X$15412 562 60 563 644 645 cell_1rw
* cell instance $15413 m0 *1 175.545,81.9
X$15413 564 60 565 644 645 cell_1rw
* cell instance $15414 m0 *1 176.25,81.9
X$15414 566 60 567 644 645 cell_1rw
* cell instance $15415 m0 *1 176.955,81.9
X$15415 568 60 569 644 645 cell_1rw
* cell instance $15416 m0 *1 177.66,81.9
X$15416 570 60 571 644 645 cell_1rw
* cell instance $15417 m0 *1 178.365,81.9
X$15417 572 60 573 644 645 cell_1rw
* cell instance $15418 m0 *1 179.07,81.9
X$15418 574 60 575 644 645 cell_1rw
* cell instance $15419 m0 *1 179.775,81.9
X$15419 576 60 577 644 645 cell_1rw
* cell instance $15420 m0 *1 180.48,81.9
X$15420 578 60 579 644 645 cell_1rw
* cell instance $15421 r0 *1 0.705,81.9
X$15421 67 61 68 644 645 cell_1rw
* cell instance $15422 r0 *1 0,81.9
X$15422 65 61 66 644 645 cell_1rw
* cell instance $15423 r0 *1 1.41,81.9
X$15423 69 61 70 644 645 cell_1rw
* cell instance $15424 r0 *1 2.115,81.9
X$15424 71 61 72 644 645 cell_1rw
* cell instance $15425 r0 *1 2.82,81.9
X$15425 73 61 74 644 645 cell_1rw
* cell instance $15426 r0 *1 3.525,81.9
X$15426 75 61 76 644 645 cell_1rw
* cell instance $15427 r0 *1 4.23,81.9
X$15427 77 61 78 644 645 cell_1rw
* cell instance $15428 r0 *1 4.935,81.9
X$15428 79 61 80 644 645 cell_1rw
* cell instance $15429 r0 *1 5.64,81.9
X$15429 81 61 82 644 645 cell_1rw
* cell instance $15430 r0 *1 6.345,81.9
X$15430 83 61 84 644 645 cell_1rw
* cell instance $15431 r0 *1 7.05,81.9
X$15431 85 61 86 644 645 cell_1rw
* cell instance $15432 r0 *1 7.755,81.9
X$15432 87 61 88 644 645 cell_1rw
* cell instance $15433 r0 *1 8.46,81.9
X$15433 89 61 90 644 645 cell_1rw
* cell instance $15434 r0 *1 9.165,81.9
X$15434 91 61 92 644 645 cell_1rw
* cell instance $15435 r0 *1 9.87,81.9
X$15435 93 61 94 644 645 cell_1rw
* cell instance $15436 r0 *1 10.575,81.9
X$15436 95 61 96 644 645 cell_1rw
* cell instance $15437 r0 *1 11.28,81.9
X$15437 97 61 98 644 645 cell_1rw
* cell instance $15438 r0 *1 11.985,81.9
X$15438 99 61 100 644 645 cell_1rw
* cell instance $15439 r0 *1 12.69,81.9
X$15439 101 61 102 644 645 cell_1rw
* cell instance $15440 r0 *1 13.395,81.9
X$15440 103 61 104 644 645 cell_1rw
* cell instance $15441 r0 *1 14.1,81.9
X$15441 105 61 106 644 645 cell_1rw
* cell instance $15442 r0 *1 14.805,81.9
X$15442 107 61 108 644 645 cell_1rw
* cell instance $15443 r0 *1 15.51,81.9
X$15443 109 61 110 644 645 cell_1rw
* cell instance $15444 r0 *1 16.215,81.9
X$15444 111 61 112 644 645 cell_1rw
* cell instance $15445 r0 *1 16.92,81.9
X$15445 113 61 114 644 645 cell_1rw
* cell instance $15446 r0 *1 17.625,81.9
X$15446 115 61 116 644 645 cell_1rw
* cell instance $15447 r0 *1 18.33,81.9
X$15447 117 61 118 644 645 cell_1rw
* cell instance $15448 r0 *1 19.035,81.9
X$15448 119 61 120 644 645 cell_1rw
* cell instance $15449 r0 *1 19.74,81.9
X$15449 121 61 122 644 645 cell_1rw
* cell instance $15450 r0 *1 20.445,81.9
X$15450 123 61 124 644 645 cell_1rw
* cell instance $15451 r0 *1 21.15,81.9
X$15451 125 61 126 644 645 cell_1rw
* cell instance $15452 r0 *1 21.855,81.9
X$15452 127 61 128 644 645 cell_1rw
* cell instance $15453 r0 *1 22.56,81.9
X$15453 129 61 130 644 645 cell_1rw
* cell instance $15454 r0 *1 23.265,81.9
X$15454 131 61 132 644 645 cell_1rw
* cell instance $15455 r0 *1 23.97,81.9
X$15455 133 61 134 644 645 cell_1rw
* cell instance $15456 r0 *1 24.675,81.9
X$15456 135 61 136 644 645 cell_1rw
* cell instance $15457 r0 *1 25.38,81.9
X$15457 137 61 138 644 645 cell_1rw
* cell instance $15458 r0 *1 26.085,81.9
X$15458 139 61 140 644 645 cell_1rw
* cell instance $15459 r0 *1 26.79,81.9
X$15459 141 61 142 644 645 cell_1rw
* cell instance $15460 r0 *1 27.495,81.9
X$15460 143 61 144 644 645 cell_1rw
* cell instance $15461 r0 *1 28.2,81.9
X$15461 145 61 146 644 645 cell_1rw
* cell instance $15462 r0 *1 28.905,81.9
X$15462 147 61 148 644 645 cell_1rw
* cell instance $15463 r0 *1 29.61,81.9
X$15463 149 61 150 644 645 cell_1rw
* cell instance $15464 r0 *1 30.315,81.9
X$15464 151 61 152 644 645 cell_1rw
* cell instance $15465 r0 *1 31.02,81.9
X$15465 153 61 154 644 645 cell_1rw
* cell instance $15466 r0 *1 31.725,81.9
X$15466 155 61 156 644 645 cell_1rw
* cell instance $15467 r0 *1 32.43,81.9
X$15467 157 61 158 644 645 cell_1rw
* cell instance $15468 r0 *1 33.135,81.9
X$15468 159 61 160 644 645 cell_1rw
* cell instance $15469 r0 *1 33.84,81.9
X$15469 161 61 162 644 645 cell_1rw
* cell instance $15470 r0 *1 34.545,81.9
X$15470 163 61 164 644 645 cell_1rw
* cell instance $15471 r0 *1 35.25,81.9
X$15471 165 61 166 644 645 cell_1rw
* cell instance $15472 r0 *1 35.955,81.9
X$15472 167 61 168 644 645 cell_1rw
* cell instance $15473 r0 *1 36.66,81.9
X$15473 169 61 170 644 645 cell_1rw
* cell instance $15474 r0 *1 37.365,81.9
X$15474 171 61 172 644 645 cell_1rw
* cell instance $15475 r0 *1 38.07,81.9
X$15475 173 61 174 644 645 cell_1rw
* cell instance $15476 r0 *1 38.775,81.9
X$15476 175 61 176 644 645 cell_1rw
* cell instance $15477 r0 *1 39.48,81.9
X$15477 177 61 178 644 645 cell_1rw
* cell instance $15478 r0 *1 40.185,81.9
X$15478 179 61 180 644 645 cell_1rw
* cell instance $15479 r0 *1 40.89,81.9
X$15479 181 61 182 644 645 cell_1rw
* cell instance $15480 r0 *1 41.595,81.9
X$15480 183 61 184 644 645 cell_1rw
* cell instance $15481 r0 *1 42.3,81.9
X$15481 185 61 186 644 645 cell_1rw
* cell instance $15482 r0 *1 43.005,81.9
X$15482 187 61 188 644 645 cell_1rw
* cell instance $15483 r0 *1 43.71,81.9
X$15483 189 61 190 644 645 cell_1rw
* cell instance $15484 r0 *1 44.415,81.9
X$15484 191 61 192 644 645 cell_1rw
* cell instance $15485 r0 *1 45.12,81.9
X$15485 193 61 194 644 645 cell_1rw
* cell instance $15486 r0 *1 45.825,81.9
X$15486 195 61 196 644 645 cell_1rw
* cell instance $15487 r0 *1 46.53,81.9
X$15487 197 61 198 644 645 cell_1rw
* cell instance $15488 r0 *1 47.235,81.9
X$15488 199 61 200 644 645 cell_1rw
* cell instance $15489 r0 *1 47.94,81.9
X$15489 201 61 202 644 645 cell_1rw
* cell instance $15490 r0 *1 48.645,81.9
X$15490 203 61 204 644 645 cell_1rw
* cell instance $15491 r0 *1 49.35,81.9
X$15491 205 61 206 644 645 cell_1rw
* cell instance $15492 r0 *1 50.055,81.9
X$15492 207 61 208 644 645 cell_1rw
* cell instance $15493 r0 *1 50.76,81.9
X$15493 209 61 210 644 645 cell_1rw
* cell instance $15494 r0 *1 51.465,81.9
X$15494 211 61 212 644 645 cell_1rw
* cell instance $15495 r0 *1 52.17,81.9
X$15495 213 61 214 644 645 cell_1rw
* cell instance $15496 r0 *1 52.875,81.9
X$15496 215 61 216 644 645 cell_1rw
* cell instance $15497 r0 *1 53.58,81.9
X$15497 217 61 218 644 645 cell_1rw
* cell instance $15498 r0 *1 54.285,81.9
X$15498 219 61 220 644 645 cell_1rw
* cell instance $15499 r0 *1 54.99,81.9
X$15499 221 61 222 644 645 cell_1rw
* cell instance $15500 r0 *1 55.695,81.9
X$15500 223 61 224 644 645 cell_1rw
* cell instance $15501 r0 *1 56.4,81.9
X$15501 225 61 226 644 645 cell_1rw
* cell instance $15502 r0 *1 57.105,81.9
X$15502 227 61 228 644 645 cell_1rw
* cell instance $15503 r0 *1 57.81,81.9
X$15503 229 61 230 644 645 cell_1rw
* cell instance $15504 r0 *1 58.515,81.9
X$15504 231 61 232 644 645 cell_1rw
* cell instance $15505 r0 *1 59.22,81.9
X$15505 233 61 234 644 645 cell_1rw
* cell instance $15506 r0 *1 59.925,81.9
X$15506 235 61 236 644 645 cell_1rw
* cell instance $15507 r0 *1 60.63,81.9
X$15507 237 61 238 644 645 cell_1rw
* cell instance $15508 r0 *1 61.335,81.9
X$15508 239 61 240 644 645 cell_1rw
* cell instance $15509 r0 *1 62.04,81.9
X$15509 241 61 242 644 645 cell_1rw
* cell instance $15510 r0 *1 62.745,81.9
X$15510 243 61 244 644 645 cell_1rw
* cell instance $15511 r0 *1 63.45,81.9
X$15511 245 61 246 644 645 cell_1rw
* cell instance $15512 r0 *1 64.155,81.9
X$15512 247 61 248 644 645 cell_1rw
* cell instance $15513 r0 *1 64.86,81.9
X$15513 249 61 250 644 645 cell_1rw
* cell instance $15514 r0 *1 65.565,81.9
X$15514 251 61 252 644 645 cell_1rw
* cell instance $15515 r0 *1 66.27,81.9
X$15515 253 61 254 644 645 cell_1rw
* cell instance $15516 r0 *1 66.975,81.9
X$15516 255 61 256 644 645 cell_1rw
* cell instance $15517 r0 *1 67.68,81.9
X$15517 257 61 258 644 645 cell_1rw
* cell instance $15518 r0 *1 68.385,81.9
X$15518 259 61 260 644 645 cell_1rw
* cell instance $15519 r0 *1 69.09,81.9
X$15519 261 61 262 644 645 cell_1rw
* cell instance $15520 r0 *1 69.795,81.9
X$15520 263 61 264 644 645 cell_1rw
* cell instance $15521 r0 *1 70.5,81.9
X$15521 265 61 266 644 645 cell_1rw
* cell instance $15522 r0 *1 71.205,81.9
X$15522 267 61 268 644 645 cell_1rw
* cell instance $15523 r0 *1 71.91,81.9
X$15523 269 61 270 644 645 cell_1rw
* cell instance $15524 r0 *1 72.615,81.9
X$15524 271 61 272 644 645 cell_1rw
* cell instance $15525 r0 *1 73.32,81.9
X$15525 273 61 274 644 645 cell_1rw
* cell instance $15526 r0 *1 74.025,81.9
X$15526 275 61 276 644 645 cell_1rw
* cell instance $15527 r0 *1 74.73,81.9
X$15527 277 61 278 644 645 cell_1rw
* cell instance $15528 r0 *1 75.435,81.9
X$15528 279 61 280 644 645 cell_1rw
* cell instance $15529 r0 *1 76.14,81.9
X$15529 281 61 282 644 645 cell_1rw
* cell instance $15530 r0 *1 76.845,81.9
X$15530 283 61 284 644 645 cell_1rw
* cell instance $15531 r0 *1 77.55,81.9
X$15531 285 61 286 644 645 cell_1rw
* cell instance $15532 r0 *1 78.255,81.9
X$15532 287 61 288 644 645 cell_1rw
* cell instance $15533 r0 *1 78.96,81.9
X$15533 289 61 290 644 645 cell_1rw
* cell instance $15534 r0 *1 79.665,81.9
X$15534 291 61 292 644 645 cell_1rw
* cell instance $15535 r0 *1 80.37,81.9
X$15535 293 61 294 644 645 cell_1rw
* cell instance $15536 r0 *1 81.075,81.9
X$15536 295 61 296 644 645 cell_1rw
* cell instance $15537 r0 *1 81.78,81.9
X$15537 297 61 298 644 645 cell_1rw
* cell instance $15538 r0 *1 82.485,81.9
X$15538 299 61 300 644 645 cell_1rw
* cell instance $15539 r0 *1 83.19,81.9
X$15539 301 61 302 644 645 cell_1rw
* cell instance $15540 r0 *1 83.895,81.9
X$15540 303 61 304 644 645 cell_1rw
* cell instance $15541 r0 *1 84.6,81.9
X$15541 305 61 306 644 645 cell_1rw
* cell instance $15542 r0 *1 85.305,81.9
X$15542 307 61 308 644 645 cell_1rw
* cell instance $15543 r0 *1 86.01,81.9
X$15543 309 61 310 644 645 cell_1rw
* cell instance $15544 r0 *1 86.715,81.9
X$15544 311 61 312 644 645 cell_1rw
* cell instance $15545 r0 *1 87.42,81.9
X$15545 313 61 314 644 645 cell_1rw
* cell instance $15546 r0 *1 88.125,81.9
X$15546 315 61 316 644 645 cell_1rw
* cell instance $15547 r0 *1 88.83,81.9
X$15547 317 61 318 644 645 cell_1rw
* cell instance $15548 r0 *1 89.535,81.9
X$15548 319 61 320 644 645 cell_1rw
* cell instance $15549 r0 *1 90.24,81.9
X$15549 321 61 323 644 645 cell_1rw
* cell instance $15550 r0 *1 90.945,81.9
X$15550 324 61 325 644 645 cell_1rw
* cell instance $15551 r0 *1 91.65,81.9
X$15551 326 61 327 644 645 cell_1rw
* cell instance $15552 r0 *1 92.355,81.9
X$15552 328 61 329 644 645 cell_1rw
* cell instance $15553 r0 *1 93.06,81.9
X$15553 330 61 331 644 645 cell_1rw
* cell instance $15554 r0 *1 93.765,81.9
X$15554 332 61 333 644 645 cell_1rw
* cell instance $15555 r0 *1 94.47,81.9
X$15555 334 61 335 644 645 cell_1rw
* cell instance $15556 r0 *1 95.175,81.9
X$15556 336 61 337 644 645 cell_1rw
* cell instance $15557 r0 *1 95.88,81.9
X$15557 338 61 339 644 645 cell_1rw
* cell instance $15558 r0 *1 96.585,81.9
X$15558 340 61 341 644 645 cell_1rw
* cell instance $15559 r0 *1 97.29,81.9
X$15559 342 61 343 644 645 cell_1rw
* cell instance $15560 r0 *1 97.995,81.9
X$15560 344 61 345 644 645 cell_1rw
* cell instance $15561 r0 *1 98.7,81.9
X$15561 346 61 347 644 645 cell_1rw
* cell instance $15562 r0 *1 99.405,81.9
X$15562 348 61 349 644 645 cell_1rw
* cell instance $15563 r0 *1 100.11,81.9
X$15563 350 61 351 644 645 cell_1rw
* cell instance $15564 r0 *1 100.815,81.9
X$15564 352 61 353 644 645 cell_1rw
* cell instance $15565 r0 *1 101.52,81.9
X$15565 354 61 355 644 645 cell_1rw
* cell instance $15566 r0 *1 102.225,81.9
X$15566 356 61 357 644 645 cell_1rw
* cell instance $15567 r0 *1 102.93,81.9
X$15567 358 61 359 644 645 cell_1rw
* cell instance $15568 r0 *1 103.635,81.9
X$15568 360 61 361 644 645 cell_1rw
* cell instance $15569 r0 *1 104.34,81.9
X$15569 362 61 363 644 645 cell_1rw
* cell instance $15570 r0 *1 105.045,81.9
X$15570 364 61 365 644 645 cell_1rw
* cell instance $15571 r0 *1 105.75,81.9
X$15571 366 61 367 644 645 cell_1rw
* cell instance $15572 r0 *1 106.455,81.9
X$15572 368 61 369 644 645 cell_1rw
* cell instance $15573 r0 *1 107.16,81.9
X$15573 370 61 371 644 645 cell_1rw
* cell instance $15574 r0 *1 107.865,81.9
X$15574 372 61 373 644 645 cell_1rw
* cell instance $15575 r0 *1 108.57,81.9
X$15575 374 61 375 644 645 cell_1rw
* cell instance $15576 r0 *1 109.275,81.9
X$15576 376 61 377 644 645 cell_1rw
* cell instance $15577 r0 *1 109.98,81.9
X$15577 378 61 379 644 645 cell_1rw
* cell instance $15578 r0 *1 110.685,81.9
X$15578 380 61 381 644 645 cell_1rw
* cell instance $15579 r0 *1 111.39,81.9
X$15579 382 61 383 644 645 cell_1rw
* cell instance $15580 r0 *1 112.095,81.9
X$15580 384 61 385 644 645 cell_1rw
* cell instance $15581 r0 *1 112.8,81.9
X$15581 386 61 387 644 645 cell_1rw
* cell instance $15582 r0 *1 113.505,81.9
X$15582 388 61 389 644 645 cell_1rw
* cell instance $15583 r0 *1 114.21,81.9
X$15583 390 61 391 644 645 cell_1rw
* cell instance $15584 r0 *1 114.915,81.9
X$15584 392 61 393 644 645 cell_1rw
* cell instance $15585 r0 *1 115.62,81.9
X$15585 394 61 395 644 645 cell_1rw
* cell instance $15586 r0 *1 116.325,81.9
X$15586 396 61 397 644 645 cell_1rw
* cell instance $15587 r0 *1 117.03,81.9
X$15587 398 61 399 644 645 cell_1rw
* cell instance $15588 r0 *1 117.735,81.9
X$15588 400 61 401 644 645 cell_1rw
* cell instance $15589 r0 *1 118.44,81.9
X$15589 402 61 403 644 645 cell_1rw
* cell instance $15590 r0 *1 119.145,81.9
X$15590 404 61 405 644 645 cell_1rw
* cell instance $15591 r0 *1 119.85,81.9
X$15591 406 61 407 644 645 cell_1rw
* cell instance $15592 r0 *1 120.555,81.9
X$15592 408 61 409 644 645 cell_1rw
* cell instance $15593 r0 *1 121.26,81.9
X$15593 410 61 411 644 645 cell_1rw
* cell instance $15594 r0 *1 121.965,81.9
X$15594 412 61 413 644 645 cell_1rw
* cell instance $15595 r0 *1 122.67,81.9
X$15595 414 61 415 644 645 cell_1rw
* cell instance $15596 r0 *1 123.375,81.9
X$15596 416 61 417 644 645 cell_1rw
* cell instance $15597 r0 *1 124.08,81.9
X$15597 418 61 419 644 645 cell_1rw
* cell instance $15598 r0 *1 124.785,81.9
X$15598 420 61 421 644 645 cell_1rw
* cell instance $15599 r0 *1 125.49,81.9
X$15599 422 61 423 644 645 cell_1rw
* cell instance $15600 r0 *1 126.195,81.9
X$15600 424 61 425 644 645 cell_1rw
* cell instance $15601 r0 *1 126.9,81.9
X$15601 426 61 427 644 645 cell_1rw
* cell instance $15602 r0 *1 127.605,81.9
X$15602 428 61 429 644 645 cell_1rw
* cell instance $15603 r0 *1 128.31,81.9
X$15603 430 61 431 644 645 cell_1rw
* cell instance $15604 r0 *1 129.015,81.9
X$15604 432 61 433 644 645 cell_1rw
* cell instance $15605 r0 *1 129.72,81.9
X$15605 434 61 435 644 645 cell_1rw
* cell instance $15606 r0 *1 130.425,81.9
X$15606 436 61 437 644 645 cell_1rw
* cell instance $15607 r0 *1 131.13,81.9
X$15607 438 61 439 644 645 cell_1rw
* cell instance $15608 r0 *1 131.835,81.9
X$15608 440 61 441 644 645 cell_1rw
* cell instance $15609 r0 *1 132.54,81.9
X$15609 442 61 443 644 645 cell_1rw
* cell instance $15610 r0 *1 133.245,81.9
X$15610 444 61 445 644 645 cell_1rw
* cell instance $15611 r0 *1 133.95,81.9
X$15611 446 61 447 644 645 cell_1rw
* cell instance $15612 r0 *1 134.655,81.9
X$15612 448 61 449 644 645 cell_1rw
* cell instance $15613 r0 *1 135.36,81.9
X$15613 450 61 451 644 645 cell_1rw
* cell instance $15614 r0 *1 136.065,81.9
X$15614 452 61 453 644 645 cell_1rw
* cell instance $15615 r0 *1 136.77,81.9
X$15615 454 61 455 644 645 cell_1rw
* cell instance $15616 r0 *1 137.475,81.9
X$15616 456 61 457 644 645 cell_1rw
* cell instance $15617 r0 *1 138.18,81.9
X$15617 458 61 459 644 645 cell_1rw
* cell instance $15618 r0 *1 138.885,81.9
X$15618 460 61 461 644 645 cell_1rw
* cell instance $15619 r0 *1 139.59,81.9
X$15619 462 61 463 644 645 cell_1rw
* cell instance $15620 r0 *1 140.295,81.9
X$15620 464 61 465 644 645 cell_1rw
* cell instance $15621 r0 *1 141,81.9
X$15621 466 61 467 644 645 cell_1rw
* cell instance $15622 r0 *1 141.705,81.9
X$15622 468 61 469 644 645 cell_1rw
* cell instance $15623 r0 *1 142.41,81.9
X$15623 470 61 471 644 645 cell_1rw
* cell instance $15624 r0 *1 143.115,81.9
X$15624 472 61 473 644 645 cell_1rw
* cell instance $15625 r0 *1 143.82,81.9
X$15625 474 61 475 644 645 cell_1rw
* cell instance $15626 r0 *1 144.525,81.9
X$15626 476 61 477 644 645 cell_1rw
* cell instance $15627 r0 *1 145.23,81.9
X$15627 478 61 479 644 645 cell_1rw
* cell instance $15628 r0 *1 145.935,81.9
X$15628 480 61 481 644 645 cell_1rw
* cell instance $15629 r0 *1 146.64,81.9
X$15629 482 61 483 644 645 cell_1rw
* cell instance $15630 r0 *1 147.345,81.9
X$15630 484 61 485 644 645 cell_1rw
* cell instance $15631 r0 *1 148.05,81.9
X$15631 486 61 487 644 645 cell_1rw
* cell instance $15632 r0 *1 148.755,81.9
X$15632 488 61 489 644 645 cell_1rw
* cell instance $15633 r0 *1 149.46,81.9
X$15633 490 61 491 644 645 cell_1rw
* cell instance $15634 r0 *1 150.165,81.9
X$15634 492 61 493 644 645 cell_1rw
* cell instance $15635 r0 *1 150.87,81.9
X$15635 494 61 495 644 645 cell_1rw
* cell instance $15636 r0 *1 151.575,81.9
X$15636 496 61 497 644 645 cell_1rw
* cell instance $15637 r0 *1 152.28,81.9
X$15637 498 61 499 644 645 cell_1rw
* cell instance $15638 r0 *1 152.985,81.9
X$15638 500 61 501 644 645 cell_1rw
* cell instance $15639 r0 *1 153.69,81.9
X$15639 502 61 503 644 645 cell_1rw
* cell instance $15640 r0 *1 154.395,81.9
X$15640 504 61 505 644 645 cell_1rw
* cell instance $15641 r0 *1 155.1,81.9
X$15641 506 61 507 644 645 cell_1rw
* cell instance $15642 r0 *1 155.805,81.9
X$15642 508 61 509 644 645 cell_1rw
* cell instance $15643 r0 *1 156.51,81.9
X$15643 510 61 511 644 645 cell_1rw
* cell instance $15644 r0 *1 157.215,81.9
X$15644 512 61 513 644 645 cell_1rw
* cell instance $15645 r0 *1 157.92,81.9
X$15645 514 61 515 644 645 cell_1rw
* cell instance $15646 r0 *1 158.625,81.9
X$15646 516 61 517 644 645 cell_1rw
* cell instance $15647 r0 *1 159.33,81.9
X$15647 518 61 519 644 645 cell_1rw
* cell instance $15648 r0 *1 160.035,81.9
X$15648 520 61 521 644 645 cell_1rw
* cell instance $15649 r0 *1 160.74,81.9
X$15649 522 61 523 644 645 cell_1rw
* cell instance $15650 r0 *1 161.445,81.9
X$15650 524 61 525 644 645 cell_1rw
* cell instance $15651 r0 *1 162.15,81.9
X$15651 526 61 527 644 645 cell_1rw
* cell instance $15652 r0 *1 162.855,81.9
X$15652 528 61 529 644 645 cell_1rw
* cell instance $15653 r0 *1 163.56,81.9
X$15653 530 61 531 644 645 cell_1rw
* cell instance $15654 r0 *1 164.265,81.9
X$15654 532 61 533 644 645 cell_1rw
* cell instance $15655 r0 *1 164.97,81.9
X$15655 534 61 535 644 645 cell_1rw
* cell instance $15656 r0 *1 165.675,81.9
X$15656 536 61 537 644 645 cell_1rw
* cell instance $15657 r0 *1 166.38,81.9
X$15657 538 61 539 644 645 cell_1rw
* cell instance $15658 r0 *1 167.085,81.9
X$15658 540 61 541 644 645 cell_1rw
* cell instance $15659 r0 *1 167.79,81.9
X$15659 542 61 543 644 645 cell_1rw
* cell instance $15660 r0 *1 168.495,81.9
X$15660 544 61 545 644 645 cell_1rw
* cell instance $15661 r0 *1 169.2,81.9
X$15661 546 61 547 644 645 cell_1rw
* cell instance $15662 r0 *1 169.905,81.9
X$15662 548 61 549 644 645 cell_1rw
* cell instance $15663 r0 *1 170.61,81.9
X$15663 550 61 551 644 645 cell_1rw
* cell instance $15664 r0 *1 171.315,81.9
X$15664 552 61 553 644 645 cell_1rw
* cell instance $15665 r0 *1 172.02,81.9
X$15665 554 61 555 644 645 cell_1rw
* cell instance $15666 r0 *1 172.725,81.9
X$15666 556 61 557 644 645 cell_1rw
* cell instance $15667 r0 *1 173.43,81.9
X$15667 558 61 559 644 645 cell_1rw
* cell instance $15668 r0 *1 174.135,81.9
X$15668 560 61 561 644 645 cell_1rw
* cell instance $15669 r0 *1 174.84,81.9
X$15669 562 61 563 644 645 cell_1rw
* cell instance $15670 r0 *1 175.545,81.9
X$15670 564 61 565 644 645 cell_1rw
* cell instance $15671 r0 *1 176.25,81.9
X$15671 566 61 567 644 645 cell_1rw
* cell instance $15672 r0 *1 176.955,81.9
X$15672 568 61 569 644 645 cell_1rw
* cell instance $15673 r0 *1 177.66,81.9
X$15673 570 61 571 644 645 cell_1rw
* cell instance $15674 r0 *1 178.365,81.9
X$15674 572 61 573 644 645 cell_1rw
* cell instance $15675 r0 *1 179.07,81.9
X$15675 574 61 575 644 645 cell_1rw
* cell instance $15676 r0 *1 179.775,81.9
X$15676 576 61 577 644 645 cell_1rw
* cell instance $15677 r0 *1 180.48,81.9
X$15677 578 61 579 644 645 cell_1rw
* cell instance $15678 m0 *1 0.705,84.63
X$15678 67 62 68 644 645 cell_1rw
* cell instance $15679 m0 *1 0,84.63
X$15679 65 62 66 644 645 cell_1rw
* cell instance $15680 m0 *1 1.41,84.63
X$15680 69 62 70 644 645 cell_1rw
* cell instance $15681 m0 *1 2.115,84.63
X$15681 71 62 72 644 645 cell_1rw
* cell instance $15682 m0 *1 2.82,84.63
X$15682 73 62 74 644 645 cell_1rw
* cell instance $15683 m0 *1 3.525,84.63
X$15683 75 62 76 644 645 cell_1rw
* cell instance $15684 m0 *1 4.23,84.63
X$15684 77 62 78 644 645 cell_1rw
* cell instance $15685 m0 *1 4.935,84.63
X$15685 79 62 80 644 645 cell_1rw
* cell instance $15686 m0 *1 5.64,84.63
X$15686 81 62 82 644 645 cell_1rw
* cell instance $15687 m0 *1 6.345,84.63
X$15687 83 62 84 644 645 cell_1rw
* cell instance $15688 m0 *1 7.05,84.63
X$15688 85 62 86 644 645 cell_1rw
* cell instance $15689 m0 *1 7.755,84.63
X$15689 87 62 88 644 645 cell_1rw
* cell instance $15690 m0 *1 8.46,84.63
X$15690 89 62 90 644 645 cell_1rw
* cell instance $15691 m0 *1 9.165,84.63
X$15691 91 62 92 644 645 cell_1rw
* cell instance $15692 m0 *1 9.87,84.63
X$15692 93 62 94 644 645 cell_1rw
* cell instance $15693 m0 *1 10.575,84.63
X$15693 95 62 96 644 645 cell_1rw
* cell instance $15694 m0 *1 11.28,84.63
X$15694 97 62 98 644 645 cell_1rw
* cell instance $15695 m0 *1 11.985,84.63
X$15695 99 62 100 644 645 cell_1rw
* cell instance $15696 m0 *1 12.69,84.63
X$15696 101 62 102 644 645 cell_1rw
* cell instance $15697 m0 *1 13.395,84.63
X$15697 103 62 104 644 645 cell_1rw
* cell instance $15698 m0 *1 14.1,84.63
X$15698 105 62 106 644 645 cell_1rw
* cell instance $15699 m0 *1 14.805,84.63
X$15699 107 62 108 644 645 cell_1rw
* cell instance $15700 m0 *1 15.51,84.63
X$15700 109 62 110 644 645 cell_1rw
* cell instance $15701 m0 *1 16.215,84.63
X$15701 111 62 112 644 645 cell_1rw
* cell instance $15702 m0 *1 16.92,84.63
X$15702 113 62 114 644 645 cell_1rw
* cell instance $15703 m0 *1 17.625,84.63
X$15703 115 62 116 644 645 cell_1rw
* cell instance $15704 m0 *1 18.33,84.63
X$15704 117 62 118 644 645 cell_1rw
* cell instance $15705 m0 *1 19.035,84.63
X$15705 119 62 120 644 645 cell_1rw
* cell instance $15706 m0 *1 19.74,84.63
X$15706 121 62 122 644 645 cell_1rw
* cell instance $15707 m0 *1 20.445,84.63
X$15707 123 62 124 644 645 cell_1rw
* cell instance $15708 m0 *1 21.15,84.63
X$15708 125 62 126 644 645 cell_1rw
* cell instance $15709 m0 *1 21.855,84.63
X$15709 127 62 128 644 645 cell_1rw
* cell instance $15710 m0 *1 22.56,84.63
X$15710 129 62 130 644 645 cell_1rw
* cell instance $15711 m0 *1 23.265,84.63
X$15711 131 62 132 644 645 cell_1rw
* cell instance $15712 m0 *1 23.97,84.63
X$15712 133 62 134 644 645 cell_1rw
* cell instance $15713 m0 *1 24.675,84.63
X$15713 135 62 136 644 645 cell_1rw
* cell instance $15714 m0 *1 25.38,84.63
X$15714 137 62 138 644 645 cell_1rw
* cell instance $15715 m0 *1 26.085,84.63
X$15715 139 62 140 644 645 cell_1rw
* cell instance $15716 m0 *1 26.79,84.63
X$15716 141 62 142 644 645 cell_1rw
* cell instance $15717 m0 *1 27.495,84.63
X$15717 143 62 144 644 645 cell_1rw
* cell instance $15718 m0 *1 28.2,84.63
X$15718 145 62 146 644 645 cell_1rw
* cell instance $15719 m0 *1 28.905,84.63
X$15719 147 62 148 644 645 cell_1rw
* cell instance $15720 m0 *1 29.61,84.63
X$15720 149 62 150 644 645 cell_1rw
* cell instance $15721 m0 *1 30.315,84.63
X$15721 151 62 152 644 645 cell_1rw
* cell instance $15722 m0 *1 31.02,84.63
X$15722 153 62 154 644 645 cell_1rw
* cell instance $15723 m0 *1 31.725,84.63
X$15723 155 62 156 644 645 cell_1rw
* cell instance $15724 m0 *1 32.43,84.63
X$15724 157 62 158 644 645 cell_1rw
* cell instance $15725 m0 *1 33.135,84.63
X$15725 159 62 160 644 645 cell_1rw
* cell instance $15726 m0 *1 33.84,84.63
X$15726 161 62 162 644 645 cell_1rw
* cell instance $15727 m0 *1 34.545,84.63
X$15727 163 62 164 644 645 cell_1rw
* cell instance $15728 m0 *1 35.25,84.63
X$15728 165 62 166 644 645 cell_1rw
* cell instance $15729 m0 *1 35.955,84.63
X$15729 167 62 168 644 645 cell_1rw
* cell instance $15730 m0 *1 36.66,84.63
X$15730 169 62 170 644 645 cell_1rw
* cell instance $15731 m0 *1 37.365,84.63
X$15731 171 62 172 644 645 cell_1rw
* cell instance $15732 m0 *1 38.07,84.63
X$15732 173 62 174 644 645 cell_1rw
* cell instance $15733 m0 *1 38.775,84.63
X$15733 175 62 176 644 645 cell_1rw
* cell instance $15734 m0 *1 39.48,84.63
X$15734 177 62 178 644 645 cell_1rw
* cell instance $15735 m0 *1 40.185,84.63
X$15735 179 62 180 644 645 cell_1rw
* cell instance $15736 m0 *1 40.89,84.63
X$15736 181 62 182 644 645 cell_1rw
* cell instance $15737 m0 *1 41.595,84.63
X$15737 183 62 184 644 645 cell_1rw
* cell instance $15738 m0 *1 42.3,84.63
X$15738 185 62 186 644 645 cell_1rw
* cell instance $15739 m0 *1 43.005,84.63
X$15739 187 62 188 644 645 cell_1rw
* cell instance $15740 m0 *1 43.71,84.63
X$15740 189 62 190 644 645 cell_1rw
* cell instance $15741 m0 *1 44.415,84.63
X$15741 191 62 192 644 645 cell_1rw
* cell instance $15742 m0 *1 45.12,84.63
X$15742 193 62 194 644 645 cell_1rw
* cell instance $15743 m0 *1 45.825,84.63
X$15743 195 62 196 644 645 cell_1rw
* cell instance $15744 m0 *1 46.53,84.63
X$15744 197 62 198 644 645 cell_1rw
* cell instance $15745 m0 *1 47.235,84.63
X$15745 199 62 200 644 645 cell_1rw
* cell instance $15746 m0 *1 47.94,84.63
X$15746 201 62 202 644 645 cell_1rw
* cell instance $15747 m0 *1 48.645,84.63
X$15747 203 62 204 644 645 cell_1rw
* cell instance $15748 m0 *1 49.35,84.63
X$15748 205 62 206 644 645 cell_1rw
* cell instance $15749 m0 *1 50.055,84.63
X$15749 207 62 208 644 645 cell_1rw
* cell instance $15750 m0 *1 50.76,84.63
X$15750 209 62 210 644 645 cell_1rw
* cell instance $15751 m0 *1 51.465,84.63
X$15751 211 62 212 644 645 cell_1rw
* cell instance $15752 m0 *1 52.17,84.63
X$15752 213 62 214 644 645 cell_1rw
* cell instance $15753 m0 *1 52.875,84.63
X$15753 215 62 216 644 645 cell_1rw
* cell instance $15754 m0 *1 53.58,84.63
X$15754 217 62 218 644 645 cell_1rw
* cell instance $15755 m0 *1 54.285,84.63
X$15755 219 62 220 644 645 cell_1rw
* cell instance $15756 m0 *1 54.99,84.63
X$15756 221 62 222 644 645 cell_1rw
* cell instance $15757 m0 *1 55.695,84.63
X$15757 223 62 224 644 645 cell_1rw
* cell instance $15758 m0 *1 56.4,84.63
X$15758 225 62 226 644 645 cell_1rw
* cell instance $15759 m0 *1 57.105,84.63
X$15759 227 62 228 644 645 cell_1rw
* cell instance $15760 m0 *1 57.81,84.63
X$15760 229 62 230 644 645 cell_1rw
* cell instance $15761 m0 *1 58.515,84.63
X$15761 231 62 232 644 645 cell_1rw
* cell instance $15762 m0 *1 59.22,84.63
X$15762 233 62 234 644 645 cell_1rw
* cell instance $15763 m0 *1 59.925,84.63
X$15763 235 62 236 644 645 cell_1rw
* cell instance $15764 m0 *1 60.63,84.63
X$15764 237 62 238 644 645 cell_1rw
* cell instance $15765 m0 *1 61.335,84.63
X$15765 239 62 240 644 645 cell_1rw
* cell instance $15766 m0 *1 62.04,84.63
X$15766 241 62 242 644 645 cell_1rw
* cell instance $15767 m0 *1 62.745,84.63
X$15767 243 62 244 644 645 cell_1rw
* cell instance $15768 m0 *1 63.45,84.63
X$15768 245 62 246 644 645 cell_1rw
* cell instance $15769 m0 *1 64.155,84.63
X$15769 247 62 248 644 645 cell_1rw
* cell instance $15770 m0 *1 64.86,84.63
X$15770 249 62 250 644 645 cell_1rw
* cell instance $15771 m0 *1 65.565,84.63
X$15771 251 62 252 644 645 cell_1rw
* cell instance $15772 m0 *1 66.27,84.63
X$15772 253 62 254 644 645 cell_1rw
* cell instance $15773 m0 *1 66.975,84.63
X$15773 255 62 256 644 645 cell_1rw
* cell instance $15774 m0 *1 67.68,84.63
X$15774 257 62 258 644 645 cell_1rw
* cell instance $15775 m0 *1 68.385,84.63
X$15775 259 62 260 644 645 cell_1rw
* cell instance $15776 m0 *1 69.09,84.63
X$15776 261 62 262 644 645 cell_1rw
* cell instance $15777 m0 *1 69.795,84.63
X$15777 263 62 264 644 645 cell_1rw
* cell instance $15778 m0 *1 70.5,84.63
X$15778 265 62 266 644 645 cell_1rw
* cell instance $15779 m0 *1 71.205,84.63
X$15779 267 62 268 644 645 cell_1rw
* cell instance $15780 m0 *1 71.91,84.63
X$15780 269 62 270 644 645 cell_1rw
* cell instance $15781 m0 *1 72.615,84.63
X$15781 271 62 272 644 645 cell_1rw
* cell instance $15782 m0 *1 73.32,84.63
X$15782 273 62 274 644 645 cell_1rw
* cell instance $15783 m0 *1 74.025,84.63
X$15783 275 62 276 644 645 cell_1rw
* cell instance $15784 m0 *1 74.73,84.63
X$15784 277 62 278 644 645 cell_1rw
* cell instance $15785 m0 *1 75.435,84.63
X$15785 279 62 280 644 645 cell_1rw
* cell instance $15786 m0 *1 76.14,84.63
X$15786 281 62 282 644 645 cell_1rw
* cell instance $15787 m0 *1 76.845,84.63
X$15787 283 62 284 644 645 cell_1rw
* cell instance $15788 m0 *1 77.55,84.63
X$15788 285 62 286 644 645 cell_1rw
* cell instance $15789 m0 *1 78.255,84.63
X$15789 287 62 288 644 645 cell_1rw
* cell instance $15790 m0 *1 78.96,84.63
X$15790 289 62 290 644 645 cell_1rw
* cell instance $15791 m0 *1 79.665,84.63
X$15791 291 62 292 644 645 cell_1rw
* cell instance $15792 m0 *1 80.37,84.63
X$15792 293 62 294 644 645 cell_1rw
* cell instance $15793 m0 *1 81.075,84.63
X$15793 295 62 296 644 645 cell_1rw
* cell instance $15794 m0 *1 81.78,84.63
X$15794 297 62 298 644 645 cell_1rw
* cell instance $15795 m0 *1 82.485,84.63
X$15795 299 62 300 644 645 cell_1rw
* cell instance $15796 m0 *1 83.19,84.63
X$15796 301 62 302 644 645 cell_1rw
* cell instance $15797 m0 *1 83.895,84.63
X$15797 303 62 304 644 645 cell_1rw
* cell instance $15798 m0 *1 84.6,84.63
X$15798 305 62 306 644 645 cell_1rw
* cell instance $15799 m0 *1 85.305,84.63
X$15799 307 62 308 644 645 cell_1rw
* cell instance $15800 m0 *1 86.01,84.63
X$15800 309 62 310 644 645 cell_1rw
* cell instance $15801 m0 *1 86.715,84.63
X$15801 311 62 312 644 645 cell_1rw
* cell instance $15802 m0 *1 87.42,84.63
X$15802 313 62 314 644 645 cell_1rw
* cell instance $15803 m0 *1 88.125,84.63
X$15803 315 62 316 644 645 cell_1rw
* cell instance $15804 m0 *1 88.83,84.63
X$15804 317 62 318 644 645 cell_1rw
* cell instance $15805 m0 *1 89.535,84.63
X$15805 319 62 320 644 645 cell_1rw
* cell instance $15806 m0 *1 90.24,84.63
X$15806 321 62 323 644 645 cell_1rw
* cell instance $15807 m0 *1 90.945,84.63
X$15807 324 62 325 644 645 cell_1rw
* cell instance $15808 m0 *1 91.65,84.63
X$15808 326 62 327 644 645 cell_1rw
* cell instance $15809 m0 *1 92.355,84.63
X$15809 328 62 329 644 645 cell_1rw
* cell instance $15810 m0 *1 93.06,84.63
X$15810 330 62 331 644 645 cell_1rw
* cell instance $15811 m0 *1 93.765,84.63
X$15811 332 62 333 644 645 cell_1rw
* cell instance $15812 m0 *1 94.47,84.63
X$15812 334 62 335 644 645 cell_1rw
* cell instance $15813 m0 *1 95.175,84.63
X$15813 336 62 337 644 645 cell_1rw
* cell instance $15814 m0 *1 95.88,84.63
X$15814 338 62 339 644 645 cell_1rw
* cell instance $15815 m0 *1 96.585,84.63
X$15815 340 62 341 644 645 cell_1rw
* cell instance $15816 m0 *1 97.29,84.63
X$15816 342 62 343 644 645 cell_1rw
* cell instance $15817 m0 *1 97.995,84.63
X$15817 344 62 345 644 645 cell_1rw
* cell instance $15818 m0 *1 98.7,84.63
X$15818 346 62 347 644 645 cell_1rw
* cell instance $15819 m0 *1 99.405,84.63
X$15819 348 62 349 644 645 cell_1rw
* cell instance $15820 m0 *1 100.11,84.63
X$15820 350 62 351 644 645 cell_1rw
* cell instance $15821 m0 *1 100.815,84.63
X$15821 352 62 353 644 645 cell_1rw
* cell instance $15822 m0 *1 101.52,84.63
X$15822 354 62 355 644 645 cell_1rw
* cell instance $15823 m0 *1 102.225,84.63
X$15823 356 62 357 644 645 cell_1rw
* cell instance $15824 m0 *1 102.93,84.63
X$15824 358 62 359 644 645 cell_1rw
* cell instance $15825 m0 *1 103.635,84.63
X$15825 360 62 361 644 645 cell_1rw
* cell instance $15826 m0 *1 104.34,84.63
X$15826 362 62 363 644 645 cell_1rw
* cell instance $15827 m0 *1 105.045,84.63
X$15827 364 62 365 644 645 cell_1rw
* cell instance $15828 m0 *1 105.75,84.63
X$15828 366 62 367 644 645 cell_1rw
* cell instance $15829 m0 *1 106.455,84.63
X$15829 368 62 369 644 645 cell_1rw
* cell instance $15830 m0 *1 107.16,84.63
X$15830 370 62 371 644 645 cell_1rw
* cell instance $15831 m0 *1 107.865,84.63
X$15831 372 62 373 644 645 cell_1rw
* cell instance $15832 m0 *1 108.57,84.63
X$15832 374 62 375 644 645 cell_1rw
* cell instance $15833 m0 *1 109.275,84.63
X$15833 376 62 377 644 645 cell_1rw
* cell instance $15834 m0 *1 109.98,84.63
X$15834 378 62 379 644 645 cell_1rw
* cell instance $15835 m0 *1 110.685,84.63
X$15835 380 62 381 644 645 cell_1rw
* cell instance $15836 m0 *1 111.39,84.63
X$15836 382 62 383 644 645 cell_1rw
* cell instance $15837 m0 *1 112.095,84.63
X$15837 384 62 385 644 645 cell_1rw
* cell instance $15838 m0 *1 112.8,84.63
X$15838 386 62 387 644 645 cell_1rw
* cell instance $15839 m0 *1 113.505,84.63
X$15839 388 62 389 644 645 cell_1rw
* cell instance $15840 m0 *1 114.21,84.63
X$15840 390 62 391 644 645 cell_1rw
* cell instance $15841 m0 *1 114.915,84.63
X$15841 392 62 393 644 645 cell_1rw
* cell instance $15842 m0 *1 115.62,84.63
X$15842 394 62 395 644 645 cell_1rw
* cell instance $15843 m0 *1 116.325,84.63
X$15843 396 62 397 644 645 cell_1rw
* cell instance $15844 m0 *1 117.03,84.63
X$15844 398 62 399 644 645 cell_1rw
* cell instance $15845 m0 *1 117.735,84.63
X$15845 400 62 401 644 645 cell_1rw
* cell instance $15846 m0 *1 118.44,84.63
X$15846 402 62 403 644 645 cell_1rw
* cell instance $15847 m0 *1 119.145,84.63
X$15847 404 62 405 644 645 cell_1rw
* cell instance $15848 m0 *1 119.85,84.63
X$15848 406 62 407 644 645 cell_1rw
* cell instance $15849 m0 *1 120.555,84.63
X$15849 408 62 409 644 645 cell_1rw
* cell instance $15850 m0 *1 121.26,84.63
X$15850 410 62 411 644 645 cell_1rw
* cell instance $15851 m0 *1 121.965,84.63
X$15851 412 62 413 644 645 cell_1rw
* cell instance $15852 m0 *1 122.67,84.63
X$15852 414 62 415 644 645 cell_1rw
* cell instance $15853 m0 *1 123.375,84.63
X$15853 416 62 417 644 645 cell_1rw
* cell instance $15854 m0 *1 124.08,84.63
X$15854 418 62 419 644 645 cell_1rw
* cell instance $15855 m0 *1 124.785,84.63
X$15855 420 62 421 644 645 cell_1rw
* cell instance $15856 m0 *1 125.49,84.63
X$15856 422 62 423 644 645 cell_1rw
* cell instance $15857 m0 *1 126.195,84.63
X$15857 424 62 425 644 645 cell_1rw
* cell instance $15858 m0 *1 126.9,84.63
X$15858 426 62 427 644 645 cell_1rw
* cell instance $15859 m0 *1 127.605,84.63
X$15859 428 62 429 644 645 cell_1rw
* cell instance $15860 m0 *1 128.31,84.63
X$15860 430 62 431 644 645 cell_1rw
* cell instance $15861 m0 *1 129.015,84.63
X$15861 432 62 433 644 645 cell_1rw
* cell instance $15862 m0 *1 129.72,84.63
X$15862 434 62 435 644 645 cell_1rw
* cell instance $15863 m0 *1 130.425,84.63
X$15863 436 62 437 644 645 cell_1rw
* cell instance $15864 m0 *1 131.13,84.63
X$15864 438 62 439 644 645 cell_1rw
* cell instance $15865 m0 *1 131.835,84.63
X$15865 440 62 441 644 645 cell_1rw
* cell instance $15866 m0 *1 132.54,84.63
X$15866 442 62 443 644 645 cell_1rw
* cell instance $15867 m0 *1 133.245,84.63
X$15867 444 62 445 644 645 cell_1rw
* cell instance $15868 m0 *1 133.95,84.63
X$15868 446 62 447 644 645 cell_1rw
* cell instance $15869 m0 *1 134.655,84.63
X$15869 448 62 449 644 645 cell_1rw
* cell instance $15870 m0 *1 135.36,84.63
X$15870 450 62 451 644 645 cell_1rw
* cell instance $15871 m0 *1 136.065,84.63
X$15871 452 62 453 644 645 cell_1rw
* cell instance $15872 m0 *1 136.77,84.63
X$15872 454 62 455 644 645 cell_1rw
* cell instance $15873 m0 *1 137.475,84.63
X$15873 456 62 457 644 645 cell_1rw
* cell instance $15874 m0 *1 138.18,84.63
X$15874 458 62 459 644 645 cell_1rw
* cell instance $15875 m0 *1 138.885,84.63
X$15875 460 62 461 644 645 cell_1rw
* cell instance $15876 m0 *1 139.59,84.63
X$15876 462 62 463 644 645 cell_1rw
* cell instance $15877 m0 *1 140.295,84.63
X$15877 464 62 465 644 645 cell_1rw
* cell instance $15878 m0 *1 141,84.63
X$15878 466 62 467 644 645 cell_1rw
* cell instance $15879 m0 *1 141.705,84.63
X$15879 468 62 469 644 645 cell_1rw
* cell instance $15880 m0 *1 142.41,84.63
X$15880 470 62 471 644 645 cell_1rw
* cell instance $15881 m0 *1 143.115,84.63
X$15881 472 62 473 644 645 cell_1rw
* cell instance $15882 m0 *1 143.82,84.63
X$15882 474 62 475 644 645 cell_1rw
* cell instance $15883 m0 *1 144.525,84.63
X$15883 476 62 477 644 645 cell_1rw
* cell instance $15884 m0 *1 145.23,84.63
X$15884 478 62 479 644 645 cell_1rw
* cell instance $15885 m0 *1 145.935,84.63
X$15885 480 62 481 644 645 cell_1rw
* cell instance $15886 m0 *1 146.64,84.63
X$15886 482 62 483 644 645 cell_1rw
* cell instance $15887 m0 *1 147.345,84.63
X$15887 484 62 485 644 645 cell_1rw
* cell instance $15888 m0 *1 148.05,84.63
X$15888 486 62 487 644 645 cell_1rw
* cell instance $15889 m0 *1 148.755,84.63
X$15889 488 62 489 644 645 cell_1rw
* cell instance $15890 m0 *1 149.46,84.63
X$15890 490 62 491 644 645 cell_1rw
* cell instance $15891 m0 *1 150.165,84.63
X$15891 492 62 493 644 645 cell_1rw
* cell instance $15892 m0 *1 150.87,84.63
X$15892 494 62 495 644 645 cell_1rw
* cell instance $15893 m0 *1 151.575,84.63
X$15893 496 62 497 644 645 cell_1rw
* cell instance $15894 m0 *1 152.28,84.63
X$15894 498 62 499 644 645 cell_1rw
* cell instance $15895 m0 *1 152.985,84.63
X$15895 500 62 501 644 645 cell_1rw
* cell instance $15896 m0 *1 153.69,84.63
X$15896 502 62 503 644 645 cell_1rw
* cell instance $15897 m0 *1 154.395,84.63
X$15897 504 62 505 644 645 cell_1rw
* cell instance $15898 m0 *1 155.1,84.63
X$15898 506 62 507 644 645 cell_1rw
* cell instance $15899 m0 *1 155.805,84.63
X$15899 508 62 509 644 645 cell_1rw
* cell instance $15900 m0 *1 156.51,84.63
X$15900 510 62 511 644 645 cell_1rw
* cell instance $15901 m0 *1 157.215,84.63
X$15901 512 62 513 644 645 cell_1rw
* cell instance $15902 m0 *1 157.92,84.63
X$15902 514 62 515 644 645 cell_1rw
* cell instance $15903 m0 *1 158.625,84.63
X$15903 516 62 517 644 645 cell_1rw
* cell instance $15904 m0 *1 159.33,84.63
X$15904 518 62 519 644 645 cell_1rw
* cell instance $15905 m0 *1 160.035,84.63
X$15905 520 62 521 644 645 cell_1rw
* cell instance $15906 m0 *1 160.74,84.63
X$15906 522 62 523 644 645 cell_1rw
* cell instance $15907 m0 *1 161.445,84.63
X$15907 524 62 525 644 645 cell_1rw
* cell instance $15908 m0 *1 162.15,84.63
X$15908 526 62 527 644 645 cell_1rw
* cell instance $15909 m0 *1 162.855,84.63
X$15909 528 62 529 644 645 cell_1rw
* cell instance $15910 m0 *1 163.56,84.63
X$15910 530 62 531 644 645 cell_1rw
* cell instance $15911 m0 *1 164.265,84.63
X$15911 532 62 533 644 645 cell_1rw
* cell instance $15912 m0 *1 164.97,84.63
X$15912 534 62 535 644 645 cell_1rw
* cell instance $15913 m0 *1 165.675,84.63
X$15913 536 62 537 644 645 cell_1rw
* cell instance $15914 m0 *1 166.38,84.63
X$15914 538 62 539 644 645 cell_1rw
* cell instance $15915 m0 *1 167.085,84.63
X$15915 540 62 541 644 645 cell_1rw
* cell instance $15916 m0 *1 167.79,84.63
X$15916 542 62 543 644 645 cell_1rw
* cell instance $15917 m0 *1 168.495,84.63
X$15917 544 62 545 644 645 cell_1rw
* cell instance $15918 m0 *1 169.2,84.63
X$15918 546 62 547 644 645 cell_1rw
* cell instance $15919 m0 *1 169.905,84.63
X$15919 548 62 549 644 645 cell_1rw
* cell instance $15920 m0 *1 170.61,84.63
X$15920 550 62 551 644 645 cell_1rw
* cell instance $15921 m0 *1 171.315,84.63
X$15921 552 62 553 644 645 cell_1rw
* cell instance $15922 m0 *1 172.02,84.63
X$15922 554 62 555 644 645 cell_1rw
* cell instance $15923 m0 *1 172.725,84.63
X$15923 556 62 557 644 645 cell_1rw
* cell instance $15924 m0 *1 173.43,84.63
X$15924 558 62 559 644 645 cell_1rw
* cell instance $15925 m0 *1 174.135,84.63
X$15925 560 62 561 644 645 cell_1rw
* cell instance $15926 m0 *1 174.84,84.63
X$15926 562 62 563 644 645 cell_1rw
* cell instance $15927 m0 *1 175.545,84.63
X$15927 564 62 565 644 645 cell_1rw
* cell instance $15928 m0 *1 176.25,84.63
X$15928 566 62 567 644 645 cell_1rw
* cell instance $15929 m0 *1 176.955,84.63
X$15929 568 62 569 644 645 cell_1rw
* cell instance $15930 m0 *1 177.66,84.63
X$15930 570 62 571 644 645 cell_1rw
* cell instance $15931 m0 *1 178.365,84.63
X$15931 572 62 573 644 645 cell_1rw
* cell instance $15932 m0 *1 179.07,84.63
X$15932 574 62 575 644 645 cell_1rw
* cell instance $15933 m0 *1 179.775,84.63
X$15933 576 62 577 644 645 cell_1rw
* cell instance $15934 m0 *1 180.48,84.63
X$15934 578 62 579 644 645 cell_1rw
* cell instance $15935 r0 *1 0.705,84.63
X$15935 67 63 68 644 645 cell_1rw
* cell instance $15936 r0 *1 0,84.63
X$15936 65 63 66 644 645 cell_1rw
* cell instance $15937 r0 *1 1.41,84.63
X$15937 69 63 70 644 645 cell_1rw
* cell instance $15938 r0 *1 2.115,84.63
X$15938 71 63 72 644 645 cell_1rw
* cell instance $15939 r0 *1 2.82,84.63
X$15939 73 63 74 644 645 cell_1rw
* cell instance $15940 r0 *1 3.525,84.63
X$15940 75 63 76 644 645 cell_1rw
* cell instance $15941 r0 *1 4.23,84.63
X$15941 77 63 78 644 645 cell_1rw
* cell instance $15942 r0 *1 4.935,84.63
X$15942 79 63 80 644 645 cell_1rw
* cell instance $15943 r0 *1 5.64,84.63
X$15943 81 63 82 644 645 cell_1rw
* cell instance $15944 r0 *1 6.345,84.63
X$15944 83 63 84 644 645 cell_1rw
* cell instance $15945 r0 *1 7.05,84.63
X$15945 85 63 86 644 645 cell_1rw
* cell instance $15946 r0 *1 7.755,84.63
X$15946 87 63 88 644 645 cell_1rw
* cell instance $15947 r0 *1 8.46,84.63
X$15947 89 63 90 644 645 cell_1rw
* cell instance $15948 r0 *1 9.165,84.63
X$15948 91 63 92 644 645 cell_1rw
* cell instance $15949 r0 *1 9.87,84.63
X$15949 93 63 94 644 645 cell_1rw
* cell instance $15950 r0 *1 10.575,84.63
X$15950 95 63 96 644 645 cell_1rw
* cell instance $15951 r0 *1 11.28,84.63
X$15951 97 63 98 644 645 cell_1rw
* cell instance $15952 r0 *1 11.985,84.63
X$15952 99 63 100 644 645 cell_1rw
* cell instance $15953 r0 *1 12.69,84.63
X$15953 101 63 102 644 645 cell_1rw
* cell instance $15954 r0 *1 13.395,84.63
X$15954 103 63 104 644 645 cell_1rw
* cell instance $15955 r0 *1 14.1,84.63
X$15955 105 63 106 644 645 cell_1rw
* cell instance $15956 r0 *1 14.805,84.63
X$15956 107 63 108 644 645 cell_1rw
* cell instance $15957 r0 *1 15.51,84.63
X$15957 109 63 110 644 645 cell_1rw
* cell instance $15958 r0 *1 16.215,84.63
X$15958 111 63 112 644 645 cell_1rw
* cell instance $15959 r0 *1 16.92,84.63
X$15959 113 63 114 644 645 cell_1rw
* cell instance $15960 r0 *1 17.625,84.63
X$15960 115 63 116 644 645 cell_1rw
* cell instance $15961 r0 *1 18.33,84.63
X$15961 117 63 118 644 645 cell_1rw
* cell instance $15962 r0 *1 19.035,84.63
X$15962 119 63 120 644 645 cell_1rw
* cell instance $15963 r0 *1 19.74,84.63
X$15963 121 63 122 644 645 cell_1rw
* cell instance $15964 r0 *1 20.445,84.63
X$15964 123 63 124 644 645 cell_1rw
* cell instance $15965 r0 *1 21.15,84.63
X$15965 125 63 126 644 645 cell_1rw
* cell instance $15966 r0 *1 21.855,84.63
X$15966 127 63 128 644 645 cell_1rw
* cell instance $15967 r0 *1 22.56,84.63
X$15967 129 63 130 644 645 cell_1rw
* cell instance $15968 r0 *1 23.265,84.63
X$15968 131 63 132 644 645 cell_1rw
* cell instance $15969 r0 *1 23.97,84.63
X$15969 133 63 134 644 645 cell_1rw
* cell instance $15970 r0 *1 24.675,84.63
X$15970 135 63 136 644 645 cell_1rw
* cell instance $15971 r0 *1 25.38,84.63
X$15971 137 63 138 644 645 cell_1rw
* cell instance $15972 r0 *1 26.085,84.63
X$15972 139 63 140 644 645 cell_1rw
* cell instance $15973 r0 *1 26.79,84.63
X$15973 141 63 142 644 645 cell_1rw
* cell instance $15974 r0 *1 27.495,84.63
X$15974 143 63 144 644 645 cell_1rw
* cell instance $15975 r0 *1 28.2,84.63
X$15975 145 63 146 644 645 cell_1rw
* cell instance $15976 r0 *1 28.905,84.63
X$15976 147 63 148 644 645 cell_1rw
* cell instance $15977 r0 *1 29.61,84.63
X$15977 149 63 150 644 645 cell_1rw
* cell instance $15978 r0 *1 30.315,84.63
X$15978 151 63 152 644 645 cell_1rw
* cell instance $15979 r0 *1 31.02,84.63
X$15979 153 63 154 644 645 cell_1rw
* cell instance $15980 r0 *1 31.725,84.63
X$15980 155 63 156 644 645 cell_1rw
* cell instance $15981 r0 *1 32.43,84.63
X$15981 157 63 158 644 645 cell_1rw
* cell instance $15982 r0 *1 33.135,84.63
X$15982 159 63 160 644 645 cell_1rw
* cell instance $15983 r0 *1 33.84,84.63
X$15983 161 63 162 644 645 cell_1rw
* cell instance $15984 r0 *1 34.545,84.63
X$15984 163 63 164 644 645 cell_1rw
* cell instance $15985 r0 *1 35.25,84.63
X$15985 165 63 166 644 645 cell_1rw
* cell instance $15986 r0 *1 35.955,84.63
X$15986 167 63 168 644 645 cell_1rw
* cell instance $15987 r0 *1 36.66,84.63
X$15987 169 63 170 644 645 cell_1rw
* cell instance $15988 r0 *1 37.365,84.63
X$15988 171 63 172 644 645 cell_1rw
* cell instance $15989 r0 *1 38.07,84.63
X$15989 173 63 174 644 645 cell_1rw
* cell instance $15990 r0 *1 38.775,84.63
X$15990 175 63 176 644 645 cell_1rw
* cell instance $15991 r0 *1 39.48,84.63
X$15991 177 63 178 644 645 cell_1rw
* cell instance $15992 r0 *1 40.185,84.63
X$15992 179 63 180 644 645 cell_1rw
* cell instance $15993 r0 *1 40.89,84.63
X$15993 181 63 182 644 645 cell_1rw
* cell instance $15994 r0 *1 41.595,84.63
X$15994 183 63 184 644 645 cell_1rw
* cell instance $15995 r0 *1 42.3,84.63
X$15995 185 63 186 644 645 cell_1rw
* cell instance $15996 r0 *1 43.005,84.63
X$15996 187 63 188 644 645 cell_1rw
* cell instance $15997 r0 *1 43.71,84.63
X$15997 189 63 190 644 645 cell_1rw
* cell instance $15998 r0 *1 44.415,84.63
X$15998 191 63 192 644 645 cell_1rw
* cell instance $15999 r0 *1 45.12,84.63
X$15999 193 63 194 644 645 cell_1rw
* cell instance $16000 r0 *1 45.825,84.63
X$16000 195 63 196 644 645 cell_1rw
* cell instance $16001 r0 *1 46.53,84.63
X$16001 197 63 198 644 645 cell_1rw
* cell instance $16002 r0 *1 47.235,84.63
X$16002 199 63 200 644 645 cell_1rw
* cell instance $16003 r0 *1 47.94,84.63
X$16003 201 63 202 644 645 cell_1rw
* cell instance $16004 r0 *1 48.645,84.63
X$16004 203 63 204 644 645 cell_1rw
* cell instance $16005 r0 *1 49.35,84.63
X$16005 205 63 206 644 645 cell_1rw
* cell instance $16006 r0 *1 50.055,84.63
X$16006 207 63 208 644 645 cell_1rw
* cell instance $16007 r0 *1 50.76,84.63
X$16007 209 63 210 644 645 cell_1rw
* cell instance $16008 r0 *1 51.465,84.63
X$16008 211 63 212 644 645 cell_1rw
* cell instance $16009 r0 *1 52.17,84.63
X$16009 213 63 214 644 645 cell_1rw
* cell instance $16010 r0 *1 52.875,84.63
X$16010 215 63 216 644 645 cell_1rw
* cell instance $16011 r0 *1 53.58,84.63
X$16011 217 63 218 644 645 cell_1rw
* cell instance $16012 r0 *1 54.285,84.63
X$16012 219 63 220 644 645 cell_1rw
* cell instance $16013 r0 *1 54.99,84.63
X$16013 221 63 222 644 645 cell_1rw
* cell instance $16014 r0 *1 55.695,84.63
X$16014 223 63 224 644 645 cell_1rw
* cell instance $16015 r0 *1 56.4,84.63
X$16015 225 63 226 644 645 cell_1rw
* cell instance $16016 r0 *1 57.105,84.63
X$16016 227 63 228 644 645 cell_1rw
* cell instance $16017 r0 *1 57.81,84.63
X$16017 229 63 230 644 645 cell_1rw
* cell instance $16018 r0 *1 58.515,84.63
X$16018 231 63 232 644 645 cell_1rw
* cell instance $16019 r0 *1 59.22,84.63
X$16019 233 63 234 644 645 cell_1rw
* cell instance $16020 r0 *1 59.925,84.63
X$16020 235 63 236 644 645 cell_1rw
* cell instance $16021 r0 *1 60.63,84.63
X$16021 237 63 238 644 645 cell_1rw
* cell instance $16022 r0 *1 61.335,84.63
X$16022 239 63 240 644 645 cell_1rw
* cell instance $16023 r0 *1 62.04,84.63
X$16023 241 63 242 644 645 cell_1rw
* cell instance $16024 r0 *1 62.745,84.63
X$16024 243 63 244 644 645 cell_1rw
* cell instance $16025 r0 *1 63.45,84.63
X$16025 245 63 246 644 645 cell_1rw
* cell instance $16026 r0 *1 64.155,84.63
X$16026 247 63 248 644 645 cell_1rw
* cell instance $16027 r0 *1 64.86,84.63
X$16027 249 63 250 644 645 cell_1rw
* cell instance $16028 r0 *1 65.565,84.63
X$16028 251 63 252 644 645 cell_1rw
* cell instance $16029 r0 *1 66.27,84.63
X$16029 253 63 254 644 645 cell_1rw
* cell instance $16030 r0 *1 66.975,84.63
X$16030 255 63 256 644 645 cell_1rw
* cell instance $16031 r0 *1 67.68,84.63
X$16031 257 63 258 644 645 cell_1rw
* cell instance $16032 r0 *1 68.385,84.63
X$16032 259 63 260 644 645 cell_1rw
* cell instance $16033 r0 *1 69.09,84.63
X$16033 261 63 262 644 645 cell_1rw
* cell instance $16034 r0 *1 69.795,84.63
X$16034 263 63 264 644 645 cell_1rw
* cell instance $16035 r0 *1 70.5,84.63
X$16035 265 63 266 644 645 cell_1rw
* cell instance $16036 r0 *1 71.205,84.63
X$16036 267 63 268 644 645 cell_1rw
* cell instance $16037 r0 *1 71.91,84.63
X$16037 269 63 270 644 645 cell_1rw
* cell instance $16038 r0 *1 72.615,84.63
X$16038 271 63 272 644 645 cell_1rw
* cell instance $16039 r0 *1 73.32,84.63
X$16039 273 63 274 644 645 cell_1rw
* cell instance $16040 r0 *1 74.025,84.63
X$16040 275 63 276 644 645 cell_1rw
* cell instance $16041 r0 *1 74.73,84.63
X$16041 277 63 278 644 645 cell_1rw
* cell instance $16042 r0 *1 75.435,84.63
X$16042 279 63 280 644 645 cell_1rw
* cell instance $16043 r0 *1 76.14,84.63
X$16043 281 63 282 644 645 cell_1rw
* cell instance $16044 r0 *1 76.845,84.63
X$16044 283 63 284 644 645 cell_1rw
* cell instance $16045 r0 *1 77.55,84.63
X$16045 285 63 286 644 645 cell_1rw
* cell instance $16046 r0 *1 78.255,84.63
X$16046 287 63 288 644 645 cell_1rw
* cell instance $16047 r0 *1 78.96,84.63
X$16047 289 63 290 644 645 cell_1rw
* cell instance $16048 r0 *1 79.665,84.63
X$16048 291 63 292 644 645 cell_1rw
* cell instance $16049 r0 *1 80.37,84.63
X$16049 293 63 294 644 645 cell_1rw
* cell instance $16050 r0 *1 81.075,84.63
X$16050 295 63 296 644 645 cell_1rw
* cell instance $16051 r0 *1 81.78,84.63
X$16051 297 63 298 644 645 cell_1rw
* cell instance $16052 r0 *1 82.485,84.63
X$16052 299 63 300 644 645 cell_1rw
* cell instance $16053 r0 *1 83.19,84.63
X$16053 301 63 302 644 645 cell_1rw
* cell instance $16054 r0 *1 83.895,84.63
X$16054 303 63 304 644 645 cell_1rw
* cell instance $16055 r0 *1 84.6,84.63
X$16055 305 63 306 644 645 cell_1rw
* cell instance $16056 r0 *1 85.305,84.63
X$16056 307 63 308 644 645 cell_1rw
* cell instance $16057 r0 *1 86.01,84.63
X$16057 309 63 310 644 645 cell_1rw
* cell instance $16058 r0 *1 86.715,84.63
X$16058 311 63 312 644 645 cell_1rw
* cell instance $16059 r0 *1 87.42,84.63
X$16059 313 63 314 644 645 cell_1rw
* cell instance $16060 r0 *1 88.125,84.63
X$16060 315 63 316 644 645 cell_1rw
* cell instance $16061 r0 *1 88.83,84.63
X$16061 317 63 318 644 645 cell_1rw
* cell instance $16062 r0 *1 89.535,84.63
X$16062 319 63 320 644 645 cell_1rw
* cell instance $16063 r0 *1 90.24,84.63
X$16063 321 63 323 644 645 cell_1rw
* cell instance $16064 r0 *1 90.945,84.63
X$16064 324 63 325 644 645 cell_1rw
* cell instance $16065 r0 *1 91.65,84.63
X$16065 326 63 327 644 645 cell_1rw
* cell instance $16066 r0 *1 92.355,84.63
X$16066 328 63 329 644 645 cell_1rw
* cell instance $16067 r0 *1 93.06,84.63
X$16067 330 63 331 644 645 cell_1rw
* cell instance $16068 r0 *1 93.765,84.63
X$16068 332 63 333 644 645 cell_1rw
* cell instance $16069 r0 *1 94.47,84.63
X$16069 334 63 335 644 645 cell_1rw
* cell instance $16070 r0 *1 95.175,84.63
X$16070 336 63 337 644 645 cell_1rw
* cell instance $16071 r0 *1 95.88,84.63
X$16071 338 63 339 644 645 cell_1rw
* cell instance $16072 r0 *1 96.585,84.63
X$16072 340 63 341 644 645 cell_1rw
* cell instance $16073 r0 *1 97.29,84.63
X$16073 342 63 343 644 645 cell_1rw
* cell instance $16074 r0 *1 97.995,84.63
X$16074 344 63 345 644 645 cell_1rw
* cell instance $16075 r0 *1 98.7,84.63
X$16075 346 63 347 644 645 cell_1rw
* cell instance $16076 r0 *1 99.405,84.63
X$16076 348 63 349 644 645 cell_1rw
* cell instance $16077 r0 *1 100.11,84.63
X$16077 350 63 351 644 645 cell_1rw
* cell instance $16078 r0 *1 100.815,84.63
X$16078 352 63 353 644 645 cell_1rw
* cell instance $16079 r0 *1 101.52,84.63
X$16079 354 63 355 644 645 cell_1rw
* cell instance $16080 r0 *1 102.225,84.63
X$16080 356 63 357 644 645 cell_1rw
* cell instance $16081 r0 *1 102.93,84.63
X$16081 358 63 359 644 645 cell_1rw
* cell instance $16082 r0 *1 103.635,84.63
X$16082 360 63 361 644 645 cell_1rw
* cell instance $16083 r0 *1 104.34,84.63
X$16083 362 63 363 644 645 cell_1rw
* cell instance $16084 r0 *1 105.045,84.63
X$16084 364 63 365 644 645 cell_1rw
* cell instance $16085 r0 *1 105.75,84.63
X$16085 366 63 367 644 645 cell_1rw
* cell instance $16086 r0 *1 106.455,84.63
X$16086 368 63 369 644 645 cell_1rw
* cell instance $16087 r0 *1 107.16,84.63
X$16087 370 63 371 644 645 cell_1rw
* cell instance $16088 r0 *1 107.865,84.63
X$16088 372 63 373 644 645 cell_1rw
* cell instance $16089 r0 *1 108.57,84.63
X$16089 374 63 375 644 645 cell_1rw
* cell instance $16090 r0 *1 109.275,84.63
X$16090 376 63 377 644 645 cell_1rw
* cell instance $16091 r0 *1 109.98,84.63
X$16091 378 63 379 644 645 cell_1rw
* cell instance $16092 r0 *1 110.685,84.63
X$16092 380 63 381 644 645 cell_1rw
* cell instance $16093 r0 *1 111.39,84.63
X$16093 382 63 383 644 645 cell_1rw
* cell instance $16094 r0 *1 112.095,84.63
X$16094 384 63 385 644 645 cell_1rw
* cell instance $16095 r0 *1 112.8,84.63
X$16095 386 63 387 644 645 cell_1rw
* cell instance $16096 r0 *1 113.505,84.63
X$16096 388 63 389 644 645 cell_1rw
* cell instance $16097 r0 *1 114.21,84.63
X$16097 390 63 391 644 645 cell_1rw
* cell instance $16098 r0 *1 114.915,84.63
X$16098 392 63 393 644 645 cell_1rw
* cell instance $16099 r0 *1 115.62,84.63
X$16099 394 63 395 644 645 cell_1rw
* cell instance $16100 r0 *1 116.325,84.63
X$16100 396 63 397 644 645 cell_1rw
* cell instance $16101 r0 *1 117.03,84.63
X$16101 398 63 399 644 645 cell_1rw
* cell instance $16102 r0 *1 117.735,84.63
X$16102 400 63 401 644 645 cell_1rw
* cell instance $16103 r0 *1 118.44,84.63
X$16103 402 63 403 644 645 cell_1rw
* cell instance $16104 r0 *1 119.145,84.63
X$16104 404 63 405 644 645 cell_1rw
* cell instance $16105 r0 *1 119.85,84.63
X$16105 406 63 407 644 645 cell_1rw
* cell instance $16106 r0 *1 120.555,84.63
X$16106 408 63 409 644 645 cell_1rw
* cell instance $16107 r0 *1 121.26,84.63
X$16107 410 63 411 644 645 cell_1rw
* cell instance $16108 r0 *1 121.965,84.63
X$16108 412 63 413 644 645 cell_1rw
* cell instance $16109 r0 *1 122.67,84.63
X$16109 414 63 415 644 645 cell_1rw
* cell instance $16110 r0 *1 123.375,84.63
X$16110 416 63 417 644 645 cell_1rw
* cell instance $16111 r0 *1 124.08,84.63
X$16111 418 63 419 644 645 cell_1rw
* cell instance $16112 r0 *1 124.785,84.63
X$16112 420 63 421 644 645 cell_1rw
* cell instance $16113 r0 *1 125.49,84.63
X$16113 422 63 423 644 645 cell_1rw
* cell instance $16114 r0 *1 126.195,84.63
X$16114 424 63 425 644 645 cell_1rw
* cell instance $16115 r0 *1 126.9,84.63
X$16115 426 63 427 644 645 cell_1rw
* cell instance $16116 r0 *1 127.605,84.63
X$16116 428 63 429 644 645 cell_1rw
* cell instance $16117 r0 *1 128.31,84.63
X$16117 430 63 431 644 645 cell_1rw
* cell instance $16118 r0 *1 129.015,84.63
X$16118 432 63 433 644 645 cell_1rw
* cell instance $16119 r0 *1 129.72,84.63
X$16119 434 63 435 644 645 cell_1rw
* cell instance $16120 r0 *1 130.425,84.63
X$16120 436 63 437 644 645 cell_1rw
* cell instance $16121 r0 *1 131.13,84.63
X$16121 438 63 439 644 645 cell_1rw
* cell instance $16122 r0 *1 131.835,84.63
X$16122 440 63 441 644 645 cell_1rw
* cell instance $16123 r0 *1 132.54,84.63
X$16123 442 63 443 644 645 cell_1rw
* cell instance $16124 r0 *1 133.245,84.63
X$16124 444 63 445 644 645 cell_1rw
* cell instance $16125 r0 *1 133.95,84.63
X$16125 446 63 447 644 645 cell_1rw
* cell instance $16126 r0 *1 134.655,84.63
X$16126 448 63 449 644 645 cell_1rw
* cell instance $16127 r0 *1 135.36,84.63
X$16127 450 63 451 644 645 cell_1rw
* cell instance $16128 r0 *1 136.065,84.63
X$16128 452 63 453 644 645 cell_1rw
* cell instance $16129 r0 *1 136.77,84.63
X$16129 454 63 455 644 645 cell_1rw
* cell instance $16130 r0 *1 137.475,84.63
X$16130 456 63 457 644 645 cell_1rw
* cell instance $16131 r0 *1 138.18,84.63
X$16131 458 63 459 644 645 cell_1rw
* cell instance $16132 r0 *1 138.885,84.63
X$16132 460 63 461 644 645 cell_1rw
* cell instance $16133 r0 *1 139.59,84.63
X$16133 462 63 463 644 645 cell_1rw
* cell instance $16134 r0 *1 140.295,84.63
X$16134 464 63 465 644 645 cell_1rw
* cell instance $16135 r0 *1 141,84.63
X$16135 466 63 467 644 645 cell_1rw
* cell instance $16136 r0 *1 141.705,84.63
X$16136 468 63 469 644 645 cell_1rw
* cell instance $16137 r0 *1 142.41,84.63
X$16137 470 63 471 644 645 cell_1rw
* cell instance $16138 r0 *1 143.115,84.63
X$16138 472 63 473 644 645 cell_1rw
* cell instance $16139 r0 *1 143.82,84.63
X$16139 474 63 475 644 645 cell_1rw
* cell instance $16140 r0 *1 144.525,84.63
X$16140 476 63 477 644 645 cell_1rw
* cell instance $16141 r0 *1 145.23,84.63
X$16141 478 63 479 644 645 cell_1rw
* cell instance $16142 r0 *1 145.935,84.63
X$16142 480 63 481 644 645 cell_1rw
* cell instance $16143 r0 *1 146.64,84.63
X$16143 482 63 483 644 645 cell_1rw
* cell instance $16144 r0 *1 147.345,84.63
X$16144 484 63 485 644 645 cell_1rw
* cell instance $16145 r0 *1 148.05,84.63
X$16145 486 63 487 644 645 cell_1rw
* cell instance $16146 r0 *1 148.755,84.63
X$16146 488 63 489 644 645 cell_1rw
* cell instance $16147 r0 *1 149.46,84.63
X$16147 490 63 491 644 645 cell_1rw
* cell instance $16148 r0 *1 150.165,84.63
X$16148 492 63 493 644 645 cell_1rw
* cell instance $16149 r0 *1 150.87,84.63
X$16149 494 63 495 644 645 cell_1rw
* cell instance $16150 r0 *1 151.575,84.63
X$16150 496 63 497 644 645 cell_1rw
* cell instance $16151 r0 *1 152.28,84.63
X$16151 498 63 499 644 645 cell_1rw
* cell instance $16152 r0 *1 152.985,84.63
X$16152 500 63 501 644 645 cell_1rw
* cell instance $16153 r0 *1 153.69,84.63
X$16153 502 63 503 644 645 cell_1rw
* cell instance $16154 r0 *1 154.395,84.63
X$16154 504 63 505 644 645 cell_1rw
* cell instance $16155 r0 *1 155.1,84.63
X$16155 506 63 507 644 645 cell_1rw
* cell instance $16156 r0 *1 155.805,84.63
X$16156 508 63 509 644 645 cell_1rw
* cell instance $16157 r0 *1 156.51,84.63
X$16157 510 63 511 644 645 cell_1rw
* cell instance $16158 r0 *1 157.215,84.63
X$16158 512 63 513 644 645 cell_1rw
* cell instance $16159 r0 *1 157.92,84.63
X$16159 514 63 515 644 645 cell_1rw
* cell instance $16160 r0 *1 158.625,84.63
X$16160 516 63 517 644 645 cell_1rw
* cell instance $16161 r0 *1 159.33,84.63
X$16161 518 63 519 644 645 cell_1rw
* cell instance $16162 r0 *1 160.035,84.63
X$16162 520 63 521 644 645 cell_1rw
* cell instance $16163 r0 *1 160.74,84.63
X$16163 522 63 523 644 645 cell_1rw
* cell instance $16164 r0 *1 161.445,84.63
X$16164 524 63 525 644 645 cell_1rw
* cell instance $16165 r0 *1 162.15,84.63
X$16165 526 63 527 644 645 cell_1rw
* cell instance $16166 r0 *1 162.855,84.63
X$16166 528 63 529 644 645 cell_1rw
* cell instance $16167 r0 *1 163.56,84.63
X$16167 530 63 531 644 645 cell_1rw
* cell instance $16168 r0 *1 164.265,84.63
X$16168 532 63 533 644 645 cell_1rw
* cell instance $16169 r0 *1 164.97,84.63
X$16169 534 63 535 644 645 cell_1rw
* cell instance $16170 r0 *1 165.675,84.63
X$16170 536 63 537 644 645 cell_1rw
* cell instance $16171 r0 *1 166.38,84.63
X$16171 538 63 539 644 645 cell_1rw
* cell instance $16172 r0 *1 167.085,84.63
X$16172 540 63 541 644 645 cell_1rw
* cell instance $16173 r0 *1 167.79,84.63
X$16173 542 63 543 644 645 cell_1rw
* cell instance $16174 r0 *1 168.495,84.63
X$16174 544 63 545 644 645 cell_1rw
* cell instance $16175 r0 *1 169.2,84.63
X$16175 546 63 547 644 645 cell_1rw
* cell instance $16176 r0 *1 169.905,84.63
X$16176 548 63 549 644 645 cell_1rw
* cell instance $16177 r0 *1 170.61,84.63
X$16177 550 63 551 644 645 cell_1rw
* cell instance $16178 r0 *1 171.315,84.63
X$16178 552 63 553 644 645 cell_1rw
* cell instance $16179 r0 *1 172.02,84.63
X$16179 554 63 555 644 645 cell_1rw
* cell instance $16180 r0 *1 172.725,84.63
X$16180 556 63 557 644 645 cell_1rw
* cell instance $16181 r0 *1 173.43,84.63
X$16181 558 63 559 644 645 cell_1rw
* cell instance $16182 r0 *1 174.135,84.63
X$16182 560 63 561 644 645 cell_1rw
* cell instance $16183 r0 *1 174.84,84.63
X$16183 562 63 563 644 645 cell_1rw
* cell instance $16184 r0 *1 175.545,84.63
X$16184 564 63 565 644 645 cell_1rw
* cell instance $16185 r0 *1 176.25,84.63
X$16185 566 63 567 644 645 cell_1rw
* cell instance $16186 r0 *1 176.955,84.63
X$16186 568 63 569 644 645 cell_1rw
* cell instance $16187 r0 *1 177.66,84.63
X$16187 570 63 571 644 645 cell_1rw
* cell instance $16188 r0 *1 178.365,84.63
X$16188 572 63 573 644 645 cell_1rw
* cell instance $16189 r0 *1 179.07,84.63
X$16189 574 63 575 644 645 cell_1rw
* cell instance $16190 r0 *1 179.775,84.63
X$16190 576 63 577 644 645 cell_1rw
* cell instance $16191 r0 *1 180.48,84.63
X$16191 578 63 579 644 645 cell_1rw
* cell instance $16192 m0 *1 0.705,87.36
X$16192 67 64 68 644 645 cell_1rw
* cell instance $16193 m0 *1 0,87.36
X$16193 65 64 66 644 645 cell_1rw
* cell instance $16194 m0 *1 1.41,87.36
X$16194 69 64 70 644 645 cell_1rw
* cell instance $16195 m0 *1 2.115,87.36
X$16195 71 64 72 644 645 cell_1rw
* cell instance $16196 m0 *1 2.82,87.36
X$16196 73 64 74 644 645 cell_1rw
* cell instance $16197 m0 *1 3.525,87.36
X$16197 75 64 76 644 645 cell_1rw
* cell instance $16198 m0 *1 4.23,87.36
X$16198 77 64 78 644 645 cell_1rw
* cell instance $16199 m0 *1 4.935,87.36
X$16199 79 64 80 644 645 cell_1rw
* cell instance $16200 m0 *1 5.64,87.36
X$16200 81 64 82 644 645 cell_1rw
* cell instance $16201 m0 *1 6.345,87.36
X$16201 83 64 84 644 645 cell_1rw
* cell instance $16202 m0 *1 7.05,87.36
X$16202 85 64 86 644 645 cell_1rw
* cell instance $16203 m0 *1 7.755,87.36
X$16203 87 64 88 644 645 cell_1rw
* cell instance $16204 m0 *1 8.46,87.36
X$16204 89 64 90 644 645 cell_1rw
* cell instance $16205 m0 *1 9.165,87.36
X$16205 91 64 92 644 645 cell_1rw
* cell instance $16206 m0 *1 9.87,87.36
X$16206 93 64 94 644 645 cell_1rw
* cell instance $16207 m0 *1 10.575,87.36
X$16207 95 64 96 644 645 cell_1rw
* cell instance $16208 m0 *1 11.28,87.36
X$16208 97 64 98 644 645 cell_1rw
* cell instance $16209 m0 *1 11.985,87.36
X$16209 99 64 100 644 645 cell_1rw
* cell instance $16210 m0 *1 12.69,87.36
X$16210 101 64 102 644 645 cell_1rw
* cell instance $16211 m0 *1 13.395,87.36
X$16211 103 64 104 644 645 cell_1rw
* cell instance $16212 m0 *1 14.1,87.36
X$16212 105 64 106 644 645 cell_1rw
* cell instance $16213 m0 *1 14.805,87.36
X$16213 107 64 108 644 645 cell_1rw
* cell instance $16214 m0 *1 15.51,87.36
X$16214 109 64 110 644 645 cell_1rw
* cell instance $16215 m0 *1 16.215,87.36
X$16215 111 64 112 644 645 cell_1rw
* cell instance $16216 m0 *1 16.92,87.36
X$16216 113 64 114 644 645 cell_1rw
* cell instance $16217 m0 *1 17.625,87.36
X$16217 115 64 116 644 645 cell_1rw
* cell instance $16218 m0 *1 18.33,87.36
X$16218 117 64 118 644 645 cell_1rw
* cell instance $16219 m0 *1 19.035,87.36
X$16219 119 64 120 644 645 cell_1rw
* cell instance $16220 m0 *1 19.74,87.36
X$16220 121 64 122 644 645 cell_1rw
* cell instance $16221 m0 *1 20.445,87.36
X$16221 123 64 124 644 645 cell_1rw
* cell instance $16222 m0 *1 21.15,87.36
X$16222 125 64 126 644 645 cell_1rw
* cell instance $16223 m0 *1 21.855,87.36
X$16223 127 64 128 644 645 cell_1rw
* cell instance $16224 m0 *1 22.56,87.36
X$16224 129 64 130 644 645 cell_1rw
* cell instance $16225 m0 *1 23.265,87.36
X$16225 131 64 132 644 645 cell_1rw
* cell instance $16226 m0 *1 23.97,87.36
X$16226 133 64 134 644 645 cell_1rw
* cell instance $16227 m0 *1 24.675,87.36
X$16227 135 64 136 644 645 cell_1rw
* cell instance $16228 m0 *1 25.38,87.36
X$16228 137 64 138 644 645 cell_1rw
* cell instance $16229 m0 *1 26.085,87.36
X$16229 139 64 140 644 645 cell_1rw
* cell instance $16230 m0 *1 26.79,87.36
X$16230 141 64 142 644 645 cell_1rw
* cell instance $16231 m0 *1 27.495,87.36
X$16231 143 64 144 644 645 cell_1rw
* cell instance $16232 m0 *1 28.2,87.36
X$16232 145 64 146 644 645 cell_1rw
* cell instance $16233 m0 *1 28.905,87.36
X$16233 147 64 148 644 645 cell_1rw
* cell instance $16234 m0 *1 29.61,87.36
X$16234 149 64 150 644 645 cell_1rw
* cell instance $16235 m0 *1 30.315,87.36
X$16235 151 64 152 644 645 cell_1rw
* cell instance $16236 m0 *1 31.02,87.36
X$16236 153 64 154 644 645 cell_1rw
* cell instance $16237 m0 *1 31.725,87.36
X$16237 155 64 156 644 645 cell_1rw
* cell instance $16238 m0 *1 32.43,87.36
X$16238 157 64 158 644 645 cell_1rw
* cell instance $16239 m0 *1 33.135,87.36
X$16239 159 64 160 644 645 cell_1rw
* cell instance $16240 m0 *1 33.84,87.36
X$16240 161 64 162 644 645 cell_1rw
* cell instance $16241 m0 *1 34.545,87.36
X$16241 163 64 164 644 645 cell_1rw
* cell instance $16242 m0 *1 35.25,87.36
X$16242 165 64 166 644 645 cell_1rw
* cell instance $16243 m0 *1 35.955,87.36
X$16243 167 64 168 644 645 cell_1rw
* cell instance $16244 m0 *1 36.66,87.36
X$16244 169 64 170 644 645 cell_1rw
* cell instance $16245 m0 *1 37.365,87.36
X$16245 171 64 172 644 645 cell_1rw
* cell instance $16246 m0 *1 38.07,87.36
X$16246 173 64 174 644 645 cell_1rw
* cell instance $16247 m0 *1 38.775,87.36
X$16247 175 64 176 644 645 cell_1rw
* cell instance $16248 m0 *1 39.48,87.36
X$16248 177 64 178 644 645 cell_1rw
* cell instance $16249 m0 *1 40.185,87.36
X$16249 179 64 180 644 645 cell_1rw
* cell instance $16250 m0 *1 40.89,87.36
X$16250 181 64 182 644 645 cell_1rw
* cell instance $16251 m0 *1 41.595,87.36
X$16251 183 64 184 644 645 cell_1rw
* cell instance $16252 m0 *1 42.3,87.36
X$16252 185 64 186 644 645 cell_1rw
* cell instance $16253 m0 *1 43.005,87.36
X$16253 187 64 188 644 645 cell_1rw
* cell instance $16254 m0 *1 43.71,87.36
X$16254 189 64 190 644 645 cell_1rw
* cell instance $16255 m0 *1 44.415,87.36
X$16255 191 64 192 644 645 cell_1rw
* cell instance $16256 m0 *1 45.12,87.36
X$16256 193 64 194 644 645 cell_1rw
* cell instance $16257 m0 *1 45.825,87.36
X$16257 195 64 196 644 645 cell_1rw
* cell instance $16258 m0 *1 46.53,87.36
X$16258 197 64 198 644 645 cell_1rw
* cell instance $16259 m0 *1 47.235,87.36
X$16259 199 64 200 644 645 cell_1rw
* cell instance $16260 m0 *1 47.94,87.36
X$16260 201 64 202 644 645 cell_1rw
* cell instance $16261 m0 *1 48.645,87.36
X$16261 203 64 204 644 645 cell_1rw
* cell instance $16262 m0 *1 49.35,87.36
X$16262 205 64 206 644 645 cell_1rw
* cell instance $16263 m0 *1 50.055,87.36
X$16263 207 64 208 644 645 cell_1rw
* cell instance $16264 m0 *1 50.76,87.36
X$16264 209 64 210 644 645 cell_1rw
* cell instance $16265 m0 *1 51.465,87.36
X$16265 211 64 212 644 645 cell_1rw
* cell instance $16266 m0 *1 52.17,87.36
X$16266 213 64 214 644 645 cell_1rw
* cell instance $16267 m0 *1 52.875,87.36
X$16267 215 64 216 644 645 cell_1rw
* cell instance $16268 m0 *1 53.58,87.36
X$16268 217 64 218 644 645 cell_1rw
* cell instance $16269 m0 *1 54.285,87.36
X$16269 219 64 220 644 645 cell_1rw
* cell instance $16270 m0 *1 54.99,87.36
X$16270 221 64 222 644 645 cell_1rw
* cell instance $16271 m0 *1 55.695,87.36
X$16271 223 64 224 644 645 cell_1rw
* cell instance $16272 m0 *1 56.4,87.36
X$16272 225 64 226 644 645 cell_1rw
* cell instance $16273 m0 *1 57.105,87.36
X$16273 227 64 228 644 645 cell_1rw
* cell instance $16274 m0 *1 57.81,87.36
X$16274 229 64 230 644 645 cell_1rw
* cell instance $16275 m0 *1 58.515,87.36
X$16275 231 64 232 644 645 cell_1rw
* cell instance $16276 m0 *1 59.22,87.36
X$16276 233 64 234 644 645 cell_1rw
* cell instance $16277 m0 *1 59.925,87.36
X$16277 235 64 236 644 645 cell_1rw
* cell instance $16278 m0 *1 60.63,87.36
X$16278 237 64 238 644 645 cell_1rw
* cell instance $16279 m0 *1 61.335,87.36
X$16279 239 64 240 644 645 cell_1rw
* cell instance $16280 m0 *1 62.04,87.36
X$16280 241 64 242 644 645 cell_1rw
* cell instance $16281 m0 *1 62.745,87.36
X$16281 243 64 244 644 645 cell_1rw
* cell instance $16282 m0 *1 63.45,87.36
X$16282 245 64 246 644 645 cell_1rw
* cell instance $16283 m0 *1 64.155,87.36
X$16283 247 64 248 644 645 cell_1rw
* cell instance $16284 m0 *1 64.86,87.36
X$16284 249 64 250 644 645 cell_1rw
* cell instance $16285 m0 *1 65.565,87.36
X$16285 251 64 252 644 645 cell_1rw
* cell instance $16286 m0 *1 66.27,87.36
X$16286 253 64 254 644 645 cell_1rw
* cell instance $16287 m0 *1 66.975,87.36
X$16287 255 64 256 644 645 cell_1rw
* cell instance $16288 m0 *1 67.68,87.36
X$16288 257 64 258 644 645 cell_1rw
* cell instance $16289 m0 *1 68.385,87.36
X$16289 259 64 260 644 645 cell_1rw
* cell instance $16290 m0 *1 69.09,87.36
X$16290 261 64 262 644 645 cell_1rw
* cell instance $16291 m0 *1 69.795,87.36
X$16291 263 64 264 644 645 cell_1rw
* cell instance $16292 m0 *1 70.5,87.36
X$16292 265 64 266 644 645 cell_1rw
* cell instance $16293 m0 *1 71.205,87.36
X$16293 267 64 268 644 645 cell_1rw
* cell instance $16294 m0 *1 71.91,87.36
X$16294 269 64 270 644 645 cell_1rw
* cell instance $16295 m0 *1 72.615,87.36
X$16295 271 64 272 644 645 cell_1rw
* cell instance $16296 m0 *1 73.32,87.36
X$16296 273 64 274 644 645 cell_1rw
* cell instance $16297 m0 *1 74.025,87.36
X$16297 275 64 276 644 645 cell_1rw
* cell instance $16298 m0 *1 74.73,87.36
X$16298 277 64 278 644 645 cell_1rw
* cell instance $16299 m0 *1 75.435,87.36
X$16299 279 64 280 644 645 cell_1rw
* cell instance $16300 m0 *1 76.14,87.36
X$16300 281 64 282 644 645 cell_1rw
* cell instance $16301 m0 *1 76.845,87.36
X$16301 283 64 284 644 645 cell_1rw
* cell instance $16302 m0 *1 77.55,87.36
X$16302 285 64 286 644 645 cell_1rw
* cell instance $16303 m0 *1 78.255,87.36
X$16303 287 64 288 644 645 cell_1rw
* cell instance $16304 m0 *1 78.96,87.36
X$16304 289 64 290 644 645 cell_1rw
* cell instance $16305 m0 *1 79.665,87.36
X$16305 291 64 292 644 645 cell_1rw
* cell instance $16306 m0 *1 80.37,87.36
X$16306 293 64 294 644 645 cell_1rw
* cell instance $16307 m0 *1 81.075,87.36
X$16307 295 64 296 644 645 cell_1rw
* cell instance $16308 m0 *1 81.78,87.36
X$16308 297 64 298 644 645 cell_1rw
* cell instance $16309 m0 *1 82.485,87.36
X$16309 299 64 300 644 645 cell_1rw
* cell instance $16310 m0 *1 83.19,87.36
X$16310 301 64 302 644 645 cell_1rw
* cell instance $16311 m0 *1 83.895,87.36
X$16311 303 64 304 644 645 cell_1rw
* cell instance $16312 m0 *1 84.6,87.36
X$16312 305 64 306 644 645 cell_1rw
* cell instance $16313 m0 *1 85.305,87.36
X$16313 307 64 308 644 645 cell_1rw
* cell instance $16314 m0 *1 86.01,87.36
X$16314 309 64 310 644 645 cell_1rw
* cell instance $16315 m0 *1 86.715,87.36
X$16315 311 64 312 644 645 cell_1rw
* cell instance $16316 m0 *1 87.42,87.36
X$16316 313 64 314 644 645 cell_1rw
* cell instance $16317 m0 *1 88.125,87.36
X$16317 315 64 316 644 645 cell_1rw
* cell instance $16318 m0 *1 88.83,87.36
X$16318 317 64 318 644 645 cell_1rw
* cell instance $16319 m0 *1 89.535,87.36
X$16319 319 64 320 644 645 cell_1rw
* cell instance $16320 m0 *1 90.24,87.36
X$16320 321 64 323 644 645 cell_1rw
* cell instance $16321 m0 *1 90.945,87.36
X$16321 324 64 325 644 645 cell_1rw
* cell instance $16322 m0 *1 91.65,87.36
X$16322 326 64 327 644 645 cell_1rw
* cell instance $16323 m0 *1 92.355,87.36
X$16323 328 64 329 644 645 cell_1rw
* cell instance $16324 m0 *1 93.06,87.36
X$16324 330 64 331 644 645 cell_1rw
* cell instance $16325 m0 *1 93.765,87.36
X$16325 332 64 333 644 645 cell_1rw
* cell instance $16326 m0 *1 94.47,87.36
X$16326 334 64 335 644 645 cell_1rw
* cell instance $16327 m0 *1 95.175,87.36
X$16327 336 64 337 644 645 cell_1rw
* cell instance $16328 m0 *1 95.88,87.36
X$16328 338 64 339 644 645 cell_1rw
* cell instance $16329 m0 *1 96.585,87.36
X$16329 340 64 341 644 645 cell_1rw
* cell instance $16330 m0 *1 97.29,87.36
X$16330 342 64 343 644 645 cell_1rw
* cell instance $16331 m0 *1 97.995,87.36
X$16331 344 64 345 644 645 cell_1rw
* cell instance $16332 m0 *1 98.7,87.36
X$16332 346 64 347 644 645 cell_1rw
* cell instance $16333 m0 *1 99.405,87.36
X$16333 348 64 349 644 645 cell_1rw
* cell instance $16334 m0 *1 100.11,87.36
X$16334 350 64 351 644 645 cell_1rw
* cell instance $16335 m0 *1 100.815,87.36
X$16335 352 64 353 644 645 cell_1rw
* cell instance $16336 m0 *1 101.52,87.36
X$16336 354 64 355 644 645 cell_1rw
* cell instance $16337 m0 *1 102.225,87.36
X$16337 356 64 357 644 645 cell_1rw
* cell instance $16338 m0 *1 102.93,87.36
X$16338 358 64 359 644 645 cell_1rw
* cell instance $16339 m0 *1 103.635,87.36
X$16339 360 64 361 644 645 cell_1rw
* cell instance $16340 m0 *1 104.34,87.36
X$16340 362 64 363 644 645 cell_1rw
* cell instance $16341 m0 *1 105.045,87.36
X$16341 364 64 365 644 645 cell_1rw
* cell instance $16342 m0 *1 105.75,87.36
X$16342 366 64 367 644 645 cell_1rw
* cell instance $16343 m0 *1 106.455,87.36
X$16343 368 64 369 644 645 cell_1rw
* cell instance $16344 m0 *1 107.16,87.36
X$16344 370 64 371 644 645 cell_1rw
* cell instance $16345 m0 *1 107.865,87.36
X$16345 372 64 373 644 645 cell_1rw
* cell instance $16346 m0 *1 108.57,87.36
X$16346 374 64 375 644 645 cell_1rw
* cell instance $16347 m0 *1 109.275,87.36
X$16347 376 64 377 644 645 cell_1rw
* cell instance $16348 m0 *1 109.98,87.36
X$16348 378 64 379 644 645 cell_1rw
* cell instance $16349 m0 *1 110.685,87.36
X$16349 380 64 381 644 645 cell_1rw
* cell instance $16350 m0 *1 111.39,87.36
X$16350 382 64 383 644 645 cell_1rw
* cell instance $16351 m0 *1 112.095,87.36
X$16351 384 64 385 644 645 cell_1rw
* cell instance $16352 m0 *1 112.8,87.36
X$16352 386 64 387 644 645 cell_1rw
* cell instance $16353 m0 *1 113.505,87.36
X$16353 388 64 389 644 645 cell_1rw
* cell instance $16354 m0 *1 114.21,87.36
X$16354 390 64 391 644 645 cell_1rw
* cell instance $16355 m0 *1 114.915,87.36
X$16355 392 64 393 644 645 cell_1rw
* cell instance $16356 m0 *1 115.62,87.36
X$16356 394 64 395 644 645 cell_1rw
* cell instance $16357 m0 *1 116.325,87.36
X$16357 396 64 397 644 645 cell_1rw
* cell instance $16358 m0 *1 117.03,87.36
X$16358 398 64 399 644 645 cell_1rw
* cell instance $16359 m0 *1 117.735,87.36
X$16359 400 64 401 644 645 cell_1rw
* cell instance $16360 m0 *1 118.44,87.36
X$16360 402 64 403 644 645 cell_1rw
* cell instance $16361 m0 *1 119.145,87.36
X$16361 404 64 405 644 645 cell_1rw
* cell instance $16362 m0 *1 119.85,87.36
X$16362 406 64 407 644 645 cell_1rw
* cell instance $16363 m0 *1 120.555,87.36
X$16363 408 64 409 644 645 cell_1rw
* cell instance $16364 m0 *1 121.26,87.36
X$16364 410 64 411 644 645 cell_1rw
* cell instance $16365 m0 *1 121.965,87.36
X$16365 412 64 413 644 645 cell_1rw
* cell instance $16366 m0 *1 122.67,87.36
X$16366 414 64 415 644 645 cell_1rw
* cell instance $16367 m0 *1 123.375,87.36
X$16367 416 64 417 644 645 cell_1rw
* cell instance $16368 m0 *1 124.08,87.36
X$16368 418 64 419 644 645 cell_1rw
* cell instance $16369 m0 *1 124.785,87.36
X$16369 420 64 421 644 645 cell_1rw
* cell instance $16370 m0 *1 125.49,87.36
X$16370 422 64 423 644 645 cell_1rw
* cell instance $16371 m0 *1 126.195,87.36
X$16371 424 64 425 644 645 cell_1rw
* cell instance $16372 m0 *1 126.9,87.36
X$16372 426 64 427 644 645 cell_1rw
* cell instance $16373 m0 *1 127.605,87.36
X$16373 428 64 429 644 645 cell_1rw
* cell instance $16374 m0 *1 128.31,87.36
X$16374 430 64 431 644 645 cell_1rw
* cell instance $16375 m0 *1 129.015,87.36
X$16375 432 64 433 644 645 cell_1rw
* cell instance $16376 m0 *1 129.72,87.36
X$16376 434 64 435 644 645 cell_1rw
* cell instance $16377 m0 *1 130.425,87.36
X$16377 436 64 437 644 645 cell_1rw
* cell instance $16378 m0 *1 131.13,87.36
X$16378 438 64 439 644 645 cell_1rw
* cell instance $16379 m0 *1 131.835,87.36
X$16379 440 64 441 644 645 cell_1rw
* cell instance $16380 m0 *1 132.54,87.36
X$16380 442 64 443 644 645 cell_1rw
* cell instance $16381 m0 *1 133.245,87.36
X$16381 444 64 445 644 645 cell_1rw
* cell instance $16382 m0 *1 133.95,87.36
X$16382 446 64 447 644 645 cell_1rw
* cell instance $16383 m0 *1 134.655,87.36
X$16383 448 64 449 644 645 cell_1rw
* cell instance $16384 m0 *1 135.36,87.36
X$16384 450 64 451 644 645 cell_1rw
* cell instance $16385 m0 *1 136.065,87.36
X$16385 452 64 453 644 645 cell_1rw
* cell instance $16386 m0 *1 136.77,87.36
X$16386 454 64 455 644 645 cell_1rw
* cell instance $16387 m0 *1 137.475,87.36
X$16387 456 64 457 644 645 cell_1rw
* cell instance $16388 m0 *1 138.18,87.36
X$16388 458 64 459 644 645 cell_1rw
* cell instance $16389 m0 *1 138.885,87.36
X$16389 460 64 461 644 645 cell_1rw
* cell instance $16390 m0 *1 139.59,87.36
X$16390 462 64 463 644 645 cell_1rw
* cell instance $16391 m0 *1 140.295,87.36
X$16391 464 64 465 644 645 cell_1rw
* cell instance $16392 m0 *1 141,87.36
X$16392 466 64 467 644 645 cell_1rw
* cell instance $16393 m0 *1 141.705,87.36
X$16393 468 64 469 644 645 cell_1rw
* cell instance $16394 m0 *1 142.41,87.36
X$16394 470 64 471 644 645 cell_1rw
* cell instance $16395 m0 *1 143.115,87.36
X$16395 472 64 473 644 645 cell_1rw
* cell instance $16396 m0 *1 143.82,87.36
X$16396 474 64 475 644 645 cell_1rw
* cell instance $16397 m0 *1 144.525,87.36
X$16397 476 64 477 644 645 cell_1rw
* cell instance $16398 m0 *1 145.23,87.36
X$16398 478 64 479 644 645 cell_1rw
* cell instance $16399 m0 *1 145.935,87.36
X$16399 480 64 481 644 645 cell_1rw
* cell instance $16400 m0 *1 146.64,87.36
X$16400 482 64 483 644 645 cell_1rw
* cell instance $16401 m0 *1 147.345,87.36
X$16401 484 64 485 644 645 cell_1rw
* cell instance $16402 m0 *1 148.05,87.36
X$16402 486 64 487 644 645 cell_1rw
* cell instance $16403 m0 *1 148.755,87.36
X$16403 488 64 489 644 645 cell_1rw
* cell instance $16404 m0 *1 149.46,87.36
X$16404 490 64 491 644 645 cell_1rw
* cell instance $16405 m0 *1 150.165,87.36
X$16405 492 64 493 644 645 cell_1rw
* cell instance $16406 m0 *1 150.87,87.36
X$16406 494 64 495 644 645 cell_1rw
* cell instance $16407 m0 *1 151.575,87.36
X$16407 496 64 497 644 645 cell_1rw
* cell instance $16408 m0 *1 152.28,87.36
X$16408 498 64 499 644 645 cell_1rw
* cell instance $16409 m0 *1 152.985,87.36
X$16409 500 64 501 644 645 cell_1rw
* cell instance $16410 m0 *1 153.69,87.36
X$16410 502 64 503 644 645 cell_1rw
* cell instance $16411 m0 *1 154.395,87.36
X$16411 504 64 505 644 645 cell_1rw
* cell instance $16412 m0 *1 155.1,87.36
X$16412 506 64 507 644 645 cell_1rw
* cell instance $16413 m0 *1 155.805,87.36
X$16413 508 64 509 644 645 cell_1rw
* cell instance $16414 m0 *1 156.51,87.36
X$16414 510 64 511 644 645 cell_1rw
* cell instance $16415 m0 *1 157.215,87.36
X$16415 512 64 513 644 645 cell_1rw
* cell instance $16416 m0 *1 157.92,87.36
X$16416 514 64 515 644 645 cell_1rw
* cell instance $16417 m0 *1 158.625,87.36
X$16417 516 64 517 644 645 cell_1rw
* cell instance $16418 m0 *1 159.33,87.36
X$16418 518 64 519 644 645 cell_1rw
* cell instance $16419 m0 *1 160.035,87.36
X$16419 520 64 521 644 645 cell_1rw
* cell instance $16420 m0 *1 160.74,87.36
X$16420 522 64 523 644 645 cell_1rw
* cell instance $16421 m0 *1 161.445,87.36
X$16421 524 64 525 644 645 cell_1rw
* cell instance $16422 m0 *1 162.15,87.36
X$16422 526 64 527 644 645 cell_1rw
* cell instance $16423 m0 *1 162.855,87.36
X$16423 528 64 529 644 645 cell_1rw
* cell instance $16424 m0 *1 163.56,87.36
X$16424 530 64 531 644 645 cell_1rw
* cell instance $16425 m0 *1 164.265,87.36
X$16425 532 64 533 644 645 cell_1rw
* cell instance $16426 m0 *1 164.97,87.36
X$16426 534 64 535 644 645 cell_1rw
* cell instance $16427 m0 *1 165.675,87.36
X$16427 536 64 537 644 645 cell_1rw
* cell instance $16428 m0 *1 166.38,87.36
X$16428 538 64 539 644 645 cell_1rw
* cell instance $16429 m0 *1 167.085,87.36
X$16429 540 64 541 644 645 cell_1rw
* cell instance $16430 m0 *1 167.79,87.36
X$16430 542 64 543 644 645 cell_1rw
* cell instance $16431 m0 *1 168.495,87.36
X$16431 544 64 545 644 645 cell_1rw
* cell instance $16432 m0 *1 169.2,87.36
X$16432 546 64 547 644 645 cell_1rw
* cell instance $16433 m0 *1 169.905,87.36
X$16433 548 64 549 644 645 cell_1rw
* cell instance $16434 m0 *1 170.61,87.36
X$16434 550 64 551 644 645 cell_1rw
* cell instance $16435 m0 *1 171.315,87.36
X$16435 552 64 553 644 645 cell_1rw
* cell instance $16436 m0 *1 172.02,87.36
X$16436 554 64 555 644 645 cell_1rw
* cell instance $16437 m0 *1 172.725,87.36
X$16437 556 64 557 644 645 cell_1rw
* cell instance $16438 m0 *1 173.43,87.36
X$16438 558 64 559 644 645 cell_1rw
* cell instance $16439 m0 *1 174.135,87.36
X$16439 560 64 561 644 645 cell_1rw
* cell instance $16440 m0 *1 174.84,87.36
X$16440 562 64 563 644 645 cell_1rw
* cell instance $16441 m0 *1 175.545,87.36
X$16441 564 64 565 644 645 cell_1rw
* cell instance $16442 m0 *1 176.25,87.36
X$16442 566 64 567 644 645 cell_1rw
* cell instance $16443 m0 *1 176.955,87.36
X$16443 568 64 569 644 645 cell_1rw
* cell instance $16444 m0 *1 177.66,87.36
X$16444 570 64 571 644 645 cell_1rw
* cell instance $16445 m0 *1 178.365,87.36
X$16445 572 64 573 644 645 cell_1rw
* cell instance $16446 m0 *1 179.07,87.36
X$16446 574 64 575 644 645 cell_1rw
* cell instance $16447 m0 *1 179.775,87.36
X$16447 576 64 577 644 645 cell_1rw
* cell instance $16448 m0 *1 180.48,87.36
X$16448 578 64 579 644 645 cell_1rw
* cell instance $16449 m0 *1 0,90.09
X$16449 65 581 66 644 645 cell_1rw
* cell instance $16450 r0 *1 0,87.36
X$16450 65 322 66 644 645 cell_1rw
* cell instance $16451 m0 *1 0,92.82
X$16451 65 583 66 644 645 cell_1rw
* cell instance $16452 r0 *1 0,90.09
X$16452 65 580 66 644 645 cell_1rw
* cell instance $16453 m0 *1 0,95.55
X$16453 65 584 66 644 645 cell_1rw
* cell instance $16454 r0 *1 0,92.82
X$16454 65 582 66 644 645 cell_1rw
* cell instance $16455 r0 *1 0,95.55
X$16455 65 585 66 644 645 cell_1rw
* cell instance $16456 m0 *1 0,98.28
X$16456 65 586 66 644 645 cell_1rw
* cell instance $16457 r0 *1 0,98.28
X$16457 65 587 66 644 645 cell_1rw
* cell instance $16458 m0 *1 0,101.01
X$16458 65 588 66 644 645 cell_1rw
* cell instance $16459 r0 *1 0,101.01
X$16459 65 589 66 644 645 cell_1rw
* cell instance $16460 m0 *1 0,103.74
X$16460 65 590 66 644 645 cell_1rw
* cell instance $16461 r0 *1 0,103.74
X$16461 65 591 66 644 645 cell_1rw
* cell instance $16462 m0 *1 0,106.47
X$16462 65 593 66 644 645 cell_1rw
* cell instance $16463 r0 *1 0,106.47
X$16463 65 592 66 644 645 cell_1rw
* cell instance $16464 m0 *1 0,109.2
X$16464 65 594 66 644 645 cell_1rw
* cell instance $16465 r0 *1 0,109.2
X$16465 65 595 66 644 645 cell_1rw
* cell instance $16466 m0 *1 0,111.93
X$16466 65 597 66 644 645 cell_1rw
* cell instance $16467 r0 *1 0,111.93
X$16467 65 596 66 644 645 cell_1rw
* cell instance $16468 m0 *1 0,114.66
X$16468 65 598 66 644 645 cell_1rw
* cell instance $16469 r0 *1 0,114.66
X$16469 65 599 66 644 645 cell_1rw
* cell instance $16470 m0 *1 0,117.39
X$16470 65 600 66 644 645 cell_1rw
* cell instance $16471 r0 *1 0,117.39
X$16471 65 601 66 644 645 cell_1rw
* cell instance $16472 m0 *1 0,120.12
X$16472 65 602 66 644 645 cell_1rw
* cell instance $16473 r0 *1 0,120.12
X$16473 65 603 66 644 645 cell_1rw
* cell instance $16474 m0 *1 0,122.85
X$16474 65 604 66 644 645 cell_1rw
* cell instance $16475 r0 *1 0,122.85
X$16475 65 605 66 644 645 cell_1rw
* cell instance $16476 m0 *1 0,125.58
X$16476 65 606 66 644 645 cell_1rw
* cell instance $16477 r0 *1 0,125.58
X$16477 65 607 66 644 645 cell_1rw
* cell instance $16478 m0 *1 0,128.31
X$16478 65 609 66 644 645 cell_1rw
* cell instance $16479 r0 *1 0,128.31
X$16479 65 608 66 644 645 cell_1rw
* cell instance $16480 m0 *1 0,131.04
X$16480 65 610 66 644 645 cell_1rw
* cell instance $16481 r0 *1 0,131.04
X$16481 65 611 66 644 645 cell_1rw
* cell instance $16482 m0 *1 0,133.77
X$16482 65 612 66 644 645 cell_1rw
* cell instance $16483 r0 *1 0,133.77
X$16483 65 613 66 644 645 cell_1rw
* cell instance $16484 m0 *1 0,136.5
X$16484 65 615 66 644 645 cell_1rw
* cell instance $16485 r0 *1 0,136.5
X$16485 65 614 66 644 645 cell_1rw
* cell instance $16486 m0 *1 0,139.23
X$16486 65 617 66 644 645 cell_1rw
* cell instance $16487 r0 *1 0,139.23
X$16487 65 616 66 644 645 cell_1rw
* cell instance $16488 m0 *1 0,141.96
X$16488 65 618 66 644 645 cell_1rw
* cell instance $16489 r0 *1 0,141.96
X$16489 65 619 66 644 645 cell_1rw
* cell instance $16490 m0 *1 0,144.69
X$16490 65 620 66 644 645 cell_1rw
* cell instance $16491 m0 *1 0,147.42
X$16491 65 622 66 644 645 cell_1rw
* cell instance $16492 r0 *1 0,144.69
X$16492 65 621 66 644 645 cell_1rw
* cell instance $16493 r0 *1 0,147.42
X$16493 65 623 66 644 645 cell_1rw
* cell instance $16494 m0 *1 0,150.15
X$16494 65 624 66 644 645 cell_1rw
* cell instance $16495 r0 *1 0,150.15
X$16495 65 625 66 644 645 cell_1rw
* cell instance $16496 m0 *1 0,152.88
X$16496 65 626 66 644 645 cell_1rw
* cell instance $16497 m0 *1 0,155.61
X$16497 65 628 66 644 645 cell_1rw
* cell instance $16498 r0 *1 0,152.88
X$16498 65 627 66 644 645 cell_1rw
* cell instance $16499 r0 *1 0,155.61
X$16499 65 629 66 644 645 cell_1rw
* cell instance $16500 m0 *1 0,158.34
X$16500 65 630 66 644 645 cell_1rw
* cell instance $16501 r0 *1 0,158.34
X$16501 65 631 66 644 645 cell_1rw
* cell instance $16502 m0 *1 0,161.07
X$16502 65 632 66 644 645 cell_1rw
* cell instance $16503 m0 *1 0,163.8
X$16503 65 634 66 644 645 cell_1rw
* cell instance $16504 r0 *1 0,161.07
X$16504 65 633 66 644 645 cell_1rw
* cell instance $16505 r0 *1 0,163.8
X$16505 65 635 66 644 645 cell_1rw
* cell instance $16506 m0 *1 0,166.53
X$16506 65 637 66 644 645 cell_1rw
* cell instance $16507 r0 *1 0,166.53
X$16507 65 636 66 644 645 cell_1rw
* cell instance $16508 m0 *1 0,169.26
X$16508 65 639 66 644 645 cell_1rw
* cell instance $16509 r0 *1 0,169.26
X$16509 65 638 66 644 645 cell_1rw
* cell instance $16510 m0 *1 0,171.99
X$16510 65 640 66 644 645 cell_1rw
* cell instance $16511 r0 *1 0,171.99
X$16511 65 641 66 644 645 cell_1rw
* cell instance $16512 m0 *1 0,174.72
X$16512 65 642 66 644 645 cell_1rw
* cell instance $16513 r0 *1 0,174.72
X$16513 65 643 66 644 645 cell_1rw
* cell instance $16514 m0 *1 0.705,90.09
X$16514 67 581 68 644 645 cell_1rw
* cell instance $16515 r0 *1 0.705,87.36
X$16515 67 322 68 644 645 cell_1rw
* cell instance $16516 r0 *1 0.705,90.09
X$16516 67 580 68 644 645 cell_1rw
* cell instance $16517 m0 *1 0.705,92.82
X$16517 67 583 68 644 645 cell_1rw
* cell instance $16518 m0 *1 0.705,95.55
X$16518 67 584 68 644 645 cell_1rw
* cell instance $16519 r0 *1 0.705,92.82
X$16519 67 582 68 644 645 cell_1rw
* cell instance $16520 r0 *1 0.705,95.55
X$16520 67 585 68 644 645 cell_1rw
* cell instance $16521 m0 *1 0.705,98.28
X$16521 67 586 68 644 645 cell_1rw
* cell instance $16522 r0 *1 0.705,98.28
X$16522 67 587 68 644 645 cell_1rw
* cell instance $16523 m0 *1 0.705,101.01
X$16523 67 588 68 644 645 cell_1rw
* cell instance $16524 r0 *1 0.705,101.01
X$16524 67 589 68 644 645 cell_1rw
* cell instance $16525 m0 *1 0.705,103.74
X$16525 67 590 68 644 645 cell_1rw
* cell instance $16526 r0 *1 0.705,103.74
X$16526 67 591 68 644 645 cell_1rw
* cell instance $16527 m0 *1 0.705,106.47
X$16527 67 593 68 644 645 cell_1rw
* cell instance $16528 m0 *1 0.705,109.2
X$16528 67 594 68 644 645 cell_1rw
* cell instance $16529 r0 *1 0.705,106.47
X$16529 67 592 68 644 645 cell_1rw
* cell instance $16530 r0 *1 0.705,109.2
X$16530 67 595 68 644 645 cell_1rw
* cell instance $16531 m0 *1 0.705,111.93
X$16531 67 597 68 644 645 cell_1rw
* cell instance $16532 r0 *1 0.705,111.93
X$16532 67 596 68 644 645 cell_1rw
* cell instance $16533 m0 *1 0.705,114.66
X$16533 67 598 68 644 645 cell_1rw
* cell instance $16534 r0 *1 0.705,114.66
X$16534 67 599 68 644 645 cell_1rw
* cell instance $16535 m0 *1 0.705,117.39
X$16535 67 600 68 644 645 cell_1rw
* cell instance $16536 r0 *1 0.705,117.39
X$16536 67 601 68 644 645 cell_1rw
* cell instance $16537 m0 *1 0.705,120.12
X$16537 67 602 68 644 645 cell_1rw
* cell instance $16538 r0 *1 0.705,120.12
X$16538 67 603 68 644 645 cell_1rw
* cell instance $16539 m0 *1 0.705,122.85
X$16539 67 604 68 644 645 cell_1rw
* cell instance $16540 r0 *1 0.705,122.85
X$16540 67 605 68 644 645 cell_1rw
* cell instance $16541 m0 *1 0.705,125.58
X$16541 67 606 68 644 645 cell_1rw
* cell instance $16542 r0 *1 0.705,125.58
X$16542 67 607 68 644 645 cell_1rw
* cell instance $16543 m0 *1 0.705,128.31
X$16543 67 609 68 644 645 cell_1rw
* cell instance $16544 r0 *1 0.705,128.31
X$16544 67 608 68 644 645 cell_1rw
* cell instance $16545 m0 *1 0.705,131.04
X$16545 67 610 68 644 645 cell_1rw
* cell instance $16546 r0 *1 0.705,131.04
X$16546 67 611 68 644 645 cell_1rw
* cell instance $16547 m0 *1 0.705,133.77
X$16547 67 612 68 644 645 cell_1rw
* cell instance $16548 r0 *1 0.705,133.77
X$16548 67 613 68 644 645 cell_1rw
* cell instance $16549 m0 *1 0.705,136.5
X$16549 67 615 68 644 645 cell_1rw
* cell instance $16550 r0 *1 0.705,136.5
X$16550 67 614 68 644 645 cell_1rw
* cell instance $16551 m0 *1 0.705,139.23
X$16551 67 617 68 644 645 cell_1rw
* cell instance $16552 r0 *1 0.705,139.23
X$16552 67 616 68 644 645 cell_1rw
* cell instance $16553 m0 *1 0.705,141.96
X$16553 67 618 68 644 645 cell_1rw
* cell instance $16554 r0 *1 0.705,141.96
X$16554 67 619 68 644 645 cell_1rw
* cell instance $16555 m0 *1 0.705,144.69
X$16555 67 620 68 644 645 cell_1rw
* cell instance $16556 m0 *1 0.705,147.42
X$16556 67 622 68 644 645 cell_1rw
* cell instance $16557 r0 *1 0.705,144.69
X$16557 67 621 68 644 645 cell_1rw
* cell instance $16558 r0 *1 0.705,147.42
X$16558 67 623 68 644 645 cell_1rw
* cell instance $16559 m0 *1 0.705,150.15
X$16559 67 624 68 644 645 cell_1rw
* cell instance $16560 r0 *1 0.705,150.15
X$16560 67 625 68 644 645 cell_1rw
* cell instance $16561 m0 *1 0.705,152.88
X$16561 67 626 68 644 645 cell_1rw
* cell instance $16562 r0 *1 0.705,152.88
X$16562 67 627 68 644 645 cell_1rw
* cell instance $16563 m0 *1 0.705,155.61
X$16563 67 628 68 644 645 cell_1rw
* cell instance $16564 r0 *1 0.705,155.61
X$16564 67 629 68 644 645 cell_1rw
* cell instance $16565 m0 *1 0.705,158.34
X$16565 67 630 68 644 645 cell_1rw
* cell instance $16566 r0 *1 0.705,158.34
X$16566 67 631 68 644 645 cell_1rw
* cell instance $16567 m0 *1 0.705,161.07
X$16567 67 632 68 644 645 cell_1rw
* cell instance $16568 r0 *1 0.705,161.07
X$16568 67 633 68 644 645 cell_1rw
* cell instance $16569 m0 *1 0.705,163.8
X$16569 67 634 68 644 645 cell_1rw
* cell instance $16570 m0 *1 0.705,166.53
X$16570 67 637 68 644 645 cell_1rw
* cell instance $16571 r0 *1 0.705,163.8
X$16571 67 635 68 644 645 cell_1rw
* cell instance $16572 r0 *1 0.705,166.53
X$16572 67 636 68 644 645 cell_1rw
* cell instance $16573 m0 *1 0.705,169.26
X$16573 67 639 68 644 645 cell_1rw
* cell instance $16574 r0 *1 0.705,169.26
X$16574 67 638 68 644 645 cell_1rw
* cell instance $16575 m0 *1 0.705,171.99
X$16575 67 640 68 644 645 cell_1rw
* cell instance $16576 r0 *1 0.705,171.99
X$16576 67 641 68 644 645 cell_1rw
* cell instance $16577 m0 *1 0.705,174.72
X$16577 67 642 68 644 645 cell_1rw
* cell instance $16578 r0 *1 0.705,174.72
X$16578 67 643 68 644 645 cell_1rw
* cell instance $16579 r0 *1 1.41,87.36
X$16579 69 322 70 644 645 cell_1rw
* cell instance $16580 m0 *1 1.41,90.09
X$16580 69 581 70 644 645 cell_1rw
* cell instance $16581 r0 *1 1.41,90.09
X$16581 69 580 70 644 645 cell_1rw
* cell instance $16582 m0 *1 1.41,92.82
X$16582 69 583 70 644 645 cell_1rw
* cell instance $16583 r0 *1 1.41,92.82
X$16583 69 582 70 644 645 cell_1rw
* cell instance $16584 m0 *1 1.41,95.55
X$16584 69 584 70 644 645 cell_1rw
* cell instance $16585 r0 *1 1.41,95.55
X$16585 69 585 70 644 645 cell_1rw
* cell instance $16586 m0 *1 1.41,98.28
X$16586 69 586 70 644 645 cell_1rw
* cell instance $16587 r0 *1 1.41,98.28
X$16587 69 587 70 644 645 cell_1rw
* cell instance $16588 m0 *1 1.41,101.01
X$16588 69 588 70 644 645 cell_1rw
* cell instance $16589 m0 *1 1.41,103.74
X$16589 69 590 70 644 645 cell_1rw
* cell instance $16590 r0 *1 1.41,101.01
X$16590 69 589 70 644 645 cell_1rw
* cell instance $16591 r0 *1 1.41,103.74
X$16591 69 591 70 644 645 cell_1rw
* cell instance $16592 m0 *1 1.41,106.47
X$16592 69 593 70 644 645 cell_1rw
* cell instance $16593 m0 *1 1.41,109.2
X$16593 69 594 70 644 645 cell_1rw
* cell instance $16594 r0 *1 1.41,106.47
X$16594 69 592 70 644 645 cell_1rw
* cell instance $16595 r0 *1 1.41,109.2
X$16595 69 595 70 644 645 cell_1rw
* cell instance $16596 m0 *1 1.41,111.93
X$16596 69 597 70 644 645 cell_1rw
* cell instance $16597 r0 *1 1.41,111.93
X$16597 69 596 70 644 645 cell_1rw
* cell instance $16598 m0 *1 1.41,114.66
X$16598 69 598 70 644 645 cell_1rw
* cell instance $16599 m0 *1 1.41,117.39
X$16599 69 600 70 644 645 cell_1rw
* cell instance $16600 r0 *1 1.41,114.66
X$16600 69 599 70 644 645 cell_1rw
* cell instance $16601 r0 *1 1.41,117.39
X$16601 69 601 70 644 645 cell_1rw
* cell instance $16602 m0 *1 1.41,120.12
X$16602 69 602 70 644 645 cell_1rw
* cell instance $16603 r0 *1 1.41,120.12
X$16603 69 603 70 644 645 cell_1rw
* cell instance $16604 m0 *1 1.41,122.85
X$16604 69 604 70 644 645 cell_1rw
* cell instance $16605 r0 *1 1.41,122.85
X$16605 69 605 70 644 645 cell_1rw
* cell instance $16606 m0 *1 1.41,125.58
X$16606 69 606 70 644 645 cell_1rw
* cell instance $16607 r0 *1 1.41,125.58
X$16607 69 607 70 644 645 cell_1rw
* cell instance $16608 m0 *1 1.41,128.31
X$16608 69 609 70 644 645 cell_1rw
* cell instance $16609 m0 *1 1.41,131.04
X$16609 69 610 70 644 645 cell_1rw
* cell instance $16610 r0 *1 1.41,128.31
X$16610 69 608 70 644 645 cell_1rw
* cell instance $16611 r0 *1 1.41,131.04
X$16611 69 611 70 644 645 cell_1rw
* cell instance $16612 m0 *1 1.41,133.77
X$16612 69 612 70 644 645 cell_1rw
* cell instance $16613 r0 *1 1.41,133.77
X$16613 69 613 70 644 645 cell_1rw
* cell instance $16614 m0 *1 1.41,136.5
X$16614 69 615 70 644 645 cell_1rw
* cell instance $16615 r0 *1 1.41,136.5
X$16615 69 614 70 644 645 cell_1rw
* cell instance $16616 m0 *1 1.41,139.23
X$16616 69 617 70 644 645 cell_1rw
* cell instance $16617 r0 *1 1.41,139.23
X$16617 69 616 70 644 645 cell_1rw
* cell instance $16618 m0 *1 1.41,141.96
X$16618 69 618 70 644 645 cell_1rw
* cell instance $16619 r0 *1 1.41,141.96
X$16619 69 619 70 644 645 cell_1rw
* cell instance $16620 m0 *1 1.41,144.69
X$16620 69 620 70 644 645 cell_1rw
* cell instance $16621 m0 *1 1.41,147.42
X$16621 69 622 70 644 645 cell_1rw
* cell instance $16622 r0 *1 1.41,144.69
X$16622 69 621 70 644 645 cell_1rw
* cell instance $16623 r0 *1 1.41,147.42
X$16623 69 623 70 644 645 cell_1rw
* cell instance $16624 m0 *1 1.41,150.15
X$16624 69 624 70 644 645 cell_1rw
* cell instance $16625 m0 *1 1.41,152.88
X$16625 69 626 70 644 645 cell_1rw
* cell instance $16626 r0 *1 1.41,150.15
X$16626 69 625 70 644 645 cell_1rw
* cell instance $16627 r0 *1 1.41,152.88
X$16627 69 627 70 644 645 cell_1rw
* cell instance $16628 m0 *1 1.41,155.61
X$16628 69 628 70 644 645 cell_1rw
* cell instance $16629 r0 *1 1.41,155.61
X$16629 69 629 70 644 645 cell_1rw
* cell instance $16630 m0 *1 1.41,158.34
X$16630 69 630 70 644 645 cell_1rw
* cell instance $16631 r0 *1 1.41,158.34
X$16631 69 631 70 644 645 cell_1rw
* cell instance $16632 m0 *1 1.41,161.07
X$16632 69 632 70 644 645 cell_1rw
* cell instance $16633 r0 *1 1.41,161.07
X$16633 69 633 70 644 645 cell_1rw
* cell instance $16634 m0 *1 1.41,163.8
X$16634 69 634 70 644 645 cell_1rw
* cell instance $16635 m0 *1 1.41,166.53
X$16635 69 637 70 644 645 cell_1rw
* cell instance $16636 r0 *1 1.41,163.8
X$16636 69 635 70 644 645 cell_1rw
* cell instance $16637 r0 *1 1.41,166.53
X$16637 69 636 70 644 645 cell_1rw
* cell instance $16638 m0 *1 1.41,169.26
X$16638 69 639 70 644 645 cell_1rw
* cell instance $16639 r0 *1 1.41,169.26
X$16639 69 638 70 644 645 cell_1rw
* cell instance $16640 m0 *1 1.41,171.99
X$16640 69 640 70 644 645 cell_1rw
* cell instance $16641 r0 *1 1.41,171.99
X$16641 69 641 70 644 645 cell_1rw
* cell instance $16642 m0 *1 1.41,174.72
X$16642 69 642 70 644 645 cell_1rw
* cell instance $16643 r0 *1 1.41,174.72
X$16643 69 643 70 644 645 cell_1rw
* cell instance $16644 r0 *1 2.115,87.36
X$16644 71 322 72 644 645 cell_1rw
* cell instance $16645 m0 *1 2.115,90.09
X$16645 71 581 72 644 645 cell_1rw
* cell instance $16646 r0 *1 2.115,90.09
X$16646 71 580 72 644 645 cell_1rw
* cell instance $16647 m0 *1 2.115,92.82
X$16647 71 583 72 644 645 cell_1rw
* cell instance $16648 r0 *1 2.115,92.82
X$16648 71 582 72 644 645 cell_1rw
* cell instance $16649 m0 *1 2.115,95.55
X$16649 71 584 72 644 645 cell_1rw
* cell instance $16650 m0 *1 2.115,98.28
X$16650 71 586 72 644 645 cell_1rw
* cell instance $16651 r0 *1 2.115,95.55
X$16651 71 585 72 644 645 cell_1rw
* cell instance $16652 m0 *1 2.115,101.01
X$16652 71 588 72 644 645 cell_1rw
* cell instance $16653 r0 *1 2.115,98.28
X$16653 71 587 72 644 645 cell_1rw
* cell instance $16654 r0 *1 2.115,101.01
X$16654 71 589 72 644 645 cell_1rw
* cell instance $16655 m0 *1 2.115,103.74
X$16655 71 590 72 644 645 cell_1rw
* cell instance $16656 r0 *1 2.115,103.74
X$16656 71 591 72 644 645 cell_1rw
* cell instance $16657 m0 *1 2.115,106.47
X$16657 71 593 72 644 645 cell_1rw
* cell instance $16658 r0 *1 2.115,106.47
X$16658 71 592 72 644 645 cell_1rw
* cell instance $16659 m0 *1 2.115,109.2
X$16659 71 594 72 644 645 cell_1rw
* cell instance $16660 r0 *1 2.115,109.2
X$16660 71 595 72 644 645 cell_1rw
* cell instance $16661 m0 *1 2.115,111.93
X$16661 71 597 72 644 645 cell_1rw
* cell instance $16662 r0 *1 2.115,111.93
X$16662 71 596 72 644 645 cell_1rw
* cell instance $16663 m0 *1 2.115,114.66
X$16663 71 598 72 644 645 cell_1rw
* cell instance $16664 r0 *1 2.115,114.66
X$16664 71 599 72 644 645 cell_1rw
* cell instance $16665 m0 *1 2.115,117.39
X$16665 71 600 72 644 645 cell_1rw
* cell instance $16666 r0 *1 2.115,117.39
X$16666 71 601 72 644 645 cell_1rw
* cell instance $16667 m0 *1 2.115,120.12
X$16667 71 602 72 644 645 cell_1rw
* cell instance $16668 r0 *1 2.115,120.12
X$16668 71 603 72 644 645 cell_1rw
* cell instance $16669 m0 *1 2.115,122.85
X$16669 71 604 72 644 645 cell_1rw
* cell instance $16670 m0 *1 2.115,125.58
X$16670 71 606 72 644 645 cell_1rw
* cell instance $16671 r0 *1 2.115,122.85
X$16671 71 605 72 644 645 cell_1rw
* cell instance $16672 r0 *1 2.115,125.58
X$16672 71 607 72 644 645 cell_1rw
* cell instance $16673 m0 *1 2.115,128.31
X$16673 71 609 72 644 645 cell_1rw
* cell instance $16674 r0 *1 2.115,128.31
X$16674 71 608 72 644 645 cell_1rw
* cell instance $16675 m0 *1 2.115,131.04
X$16675 71 610 72 644 645 cell_1rw
* cell instance $16676 r0 *1 2.115,131.04
X$16676 71 611 72 644 645 cell_1rw
* cell instance $16677 m0 *1 2.115,133.77
X$16677 71 612 72 644 645 cell_1rw
* cell instance $16678 m0 *1 2.115,136.5
X$16678 71 615 72 644 645 cell_1rw
* cell instance $16679 r0 *1 2.115,133.77
X$16679 71 613 72 644 645 cell_1rw
* cell instance $16680 r0 *1 2.115,136.5
X$16680 71 614 72 644 645 cell_1rw
* cell instance $16681 m0 *1 2.115,139.23
X$16681 71 617 72 644 645 cell_1rw
* cell instance $16682 r0 *1 2.115,139.23
X$16682 71 616 72 644 645 cell_1rw
* cell instance $16683 m0 *1 2.115,141.96
X$16683 71 618 72 644 645 cell_1rw
* cell instance $16684 r0 *1 2.115,141.96
X$16684 71 619 72 644 645 cell_1rw
* cell instance $16685 m0 *1 2.115,144.69
X$16685 71 620 72 644 645 cell_1rw
* cell instance $16686 r0 *1 2.115,144.69
X$16686 71 621 72 644 645 cell_1rw
* cell instance $16687 m0 *1 2.115,147.42
X$16687 71 622 72 644 645 cell_1rw
* cell instance $16688 m0 *1 2.115,150.15
X$16688 71 624 72 644 645 cell_1rw
* cell instance $16689 r0 *1 2.115,147.42
X$16689 71 623 72 644 645 cell_1rw
* cell instance $16690 r0 *1 2.115,150.15
X$16690 71 625 72 644 645 cell_1rw
* cell instance $16691 m0 *1 2.115,152.88
X$16691 71 626 72 644 645 cell_1rw
* cell instance $16692 m0 *1 2.115,155.61
X$16692 71 628 72 644 645 cell_1rw
* cell instance $16693 r0 *1 2.115,152.88
X$16693 71 627 72 644 645 cell_1rw
* cell instance $16694 r0 *1 2.115,155.61
X$16694 71 629 72 644 645 cell_1rw
* cell instance $16695 m0 *1 2.115,158.34
X$16695 71 630 72 644 645 cell_1rw
* cell instance $16696 r0 *1 2.115,158.34
X$16696 71 631 72 644 645 cell_1rw
* cell instance $16697 m0 *1 2.115,161.07
X$16697 71 632 72 644 645 cell_1rw
* cell instance $16698 r0 *1 2.115,161.07
X$16698 71 633 72 644 645 cell_1rw
* cell instance $16699 m0 *1 2.115,163.8
X$16699 71 634 72 644 645 cell_1rw
* cell instance $16700 r0 *1 2.115,163.8
X$16700 71 635 72 644 645 cell_1rw
* cell instance $16701 m0 *1 2.115,166.53
X$16701 71 637 72 644 645 cell_1rw
* cell instance $16702 r0 *1 2.115,166.53
X$16702 71 636 72 644 645 cell_1rw
* cell instance $16703 m0 *1 2.115,169.26
X$16703 71 639 72 644 645 cell_1rw
* cell instance $16704 r0 *1 2.115,169.26
X$16704 71 638 72 644 645 cell_1rw
* cell instance $16705 m0 *1 2.115,171.99
X$16705 71 640 72 644 645 cell_1rw
* cell instance $16706 r0 *1 2.115,171.99
X$16706 71 641 72 644 645 cell_1rw
* cell instance $16707 m0 *1 2.115,174.72
X$16707 71 642 72 644 645 cell_1rw
* cell instance $16708 r0 *1 2.115,174.72
X$16708 71 643 72 644 645 cell_1rw
* cell instance $16709 r0 *1 2.82,87.36
X$16709 73 322 74 644 645 cell_1rw
* cell instance $16710 m0 *1 2.82,90.09
X$16710 73 581 74 644 645 cell_1rw
* cell instance $16711 r0 *1 2.82,90.09
X$16711 73 580 74 644 645 cell_1rw
* cell instance $16712 m0 *1 2.82,92.82
X$16712 73 583 74 644 645 cell_1rw
* cell instance $16713 r0 *1 2.82,92.82
X$16713 73 582 74 644 645 cell_1rw
* cell instance $16714 m0 *1 2.82,95.55
X$16714 73 584 74 644 645 cell_1rw
* cell instance $16715 r0 *1 2.82,95.55
X$16715 73 585 74 644 645 cell_1rw
* cell instance $16716 m0 *1 2.82,98.28
X$16716 73 586 74 644 645 cell_1rw
* cell instance $16717 r0 *1 2.82,98.28
X$16717 73 587 74 644 645 cell_1rw
* cell instance $16718 m0 *1 2.82,101.01
X$16718 73 588 74 644 645 cell_1rw
* cell instance $16719 r0 *1 2.82,101.01
X$16719 73 589 74 644 645 cell_1rw
* cell instance $16720 m0 *1 2.82,103.74
X$16720 73 590 74 644 645 cell_1rw
* cell instance $16721 m0 *1 2.82,106.47
X$16721 73 593 74 644 645 cell_1rw
* cell instance $16722 r0 *1 2.82,103.74
X$16722 73 591 74 644 645 cell_1rw
* cell instance $16723 m0 *1 2.82,109.2
X$16723 73 594 74 644 645 cell_1rw
* cell instance $16724 r0 *1 2.82,106.47
X$16724 73 592 74 644 645 cell_1rw
* cell instance $16725 m0 *1 2.82,111.93
X$16725 73 597 74 644 645 cell_1rw
* cell instance $16726 r0 *1 2.82,109.2
X$16726 73 595 74 644 645 cell_1rw
* cell instance $16727 r0 *1 2.82,111.93
X$16727 73 596 74 644 645 cell_1rw
* cell instance $16728 m0 *1 2.82,114.66
X$16728 73 598 74 644 645 cell_1rw
* cell instance $16729 r0 *1 2.82,114.66
X$16729 73 599 74 644 645 cell_1rw
* cell instance $16730 m0 *1 2.82,117.39
X$16730 73 600 74 644 645 cell_1rw
* cell instance $16731 r0 *1 2.82,117.39
X$16731 73 601 74 644 645 cell_1rw
* cell instance $16732 m0 *1 2.82,120.12
X$16732 73 602 74 644 645 cell_1rw
* cell instance $16733 r0 *1 2.82,120.12
X$16733 73 603 74 644 645 cell_1rw
* cell instance $16734 m0 *1 2.82,122.85
X$16734 73 604 74 644 645 cell_1rw
* cell instance $16735 r0 *1 2.82,122.85
X$16735 73 605 74 644 645 cell_1rw
* cell instance $16736 m0 *1 2.82,125.58
X$16736 73 606 74 644 645 cell_1rw
* cell instance $16737 r0 *1 2.82,125.58
X$16737 73 607 74 644 645 cell_1rw
* cell instance $16738 m0 *1 2.82,128.31
X$16738 73 609 74 644 645 cell_1rw
* cell instance $16739 r0 *1 2.82,128.31
X$16739 73 608 74 644 645 cell_1rw
* cell instance $16740 m0 *1 2.82,131.04
X$16740 73 610 74 644 645 cell_1rw
* cell instance $16741 m0 *1 2.82,133.77
X$16741 73 612 74 644 645 cell_1rw
* cell instance $16742 r0 *1 2.82,131.04
X$16742 73 611 74 644 645 cell_1rw
* cell instance $16743 r0 *1 2.82,133.77
X$16743 73 613 74 644 645 cell_1rw
* cell instance $16744 m0 *1 2.82,136.5
X$16744 73 615 74 644 645 cell_1rw
* cell instance $16745 m0 *1 2.82,139.23
X$16745 73 617 74 644 645 cell_1rw
* cell instance $16746 r0 *1 2.82,136.5
X$16746 73 614 74 644 645 cell_1rw
* cell instance $16747 r0 *1 2.82,139.23
X$16747 73 616 74 644 645 cell_1rw
* cell instance $16748 m0 *1 2.82,141.96
X$16748 73 618 74 644 645 cell_1rw
* cell instance $16749 m0 *1 2.82,144.69
X$16749 73 620 74 644 645 cell_1rw
* cell instance $16750 r0 *1 2.82,141.96
X$16750 73 619 74 644 645 cell_1rw
* cell instance $16751 r0 *1 2.82,144.69
X$16751 73 621 74 644 645 cell_1rw
* cell instance $16752 m0 *1 2.82,147.42
X$16752 73 622 74 644 645 cell_1rw
* cell instance $16753 r0 *1 2.82,147.42
X$16753 73 623 74 644 645 cell_1rw
* cell instance $16754 m0 *1 2.82,150.15
X$16754 73 624 74 644 645 cell_1rw
* cell instance $16755 r0 *1 2.82,150.15
X$16755 73 625 74 644 645 cell_1rw
* cell instance $16756 m0 *1 2.82,152.88
X$16756 73 626 74 644 645 cell_1rw
* cell instance $16757 r0 *1 2.82,152.88
X$16757 73 627 74 644 645 cell_1rw
* cell instance $16758 m0 *1 2.82,155.61
X$16758 73 628 74 644 645 cell_1rw
* cell instance $16759 r0 *1 2.82,155.61
X$16759 73 629 74 644 645 cell_1rw
* cell instance $16760 m0 *1 2.82,158.34
X$16760 73 630 74 644 645 cell_1rw
* cell instance $16761 r0 *1 2.82,158.34
X$16761 73 631 74 644 645 cell_1rw
* cell instance $16762 m0 *1 2.82,161.07
X$16762 73 632 74 644 645 cell_1rw
* cell instance $16763 r0 *1 2.82,161.07
X$16763 73 633 74 644 645 cell_1rw
* cell instance $16764 m0 *1 2.82,163.8
X$16764 73 634 74 644 645 cell_1rw
* cell instance $16765 r0 *1 2.82,163.8
X$16765 73 635 74 644 645 cell_1rw
* cell instance $16766 m0 *1 2.82,166.53
X$16766 73 637 74 644 645 cell_1rw
* cell instance $16767 r0 *1 2.82,166.53
X$16767 73 636 74 644 645 cell_1rw
* cell instance $16768 m0 *1 2.82,169.26
X$16768 73 639 74 644 645 cell_1rw
* cell instance $16769 r0 *1 2.82,169.26
X$16769 73 638 74 644 645 cell_1rw
* cell instance $16770 m0 *1 2.82,171.99
X$16770 73 640 74 644 645 cell_1rw
* cell instance $16771 r0 *1 2.82,171.99
X$16771 73 641 74 644 645 cell_1rw
* cell instance $16772 m0 *1 2.82,174.72
X$16772 73 642 74 644 645 cell_1rw
* cell instance $16773 r0 *1 2.82,174.72
X$16773 73 643 74 644 645 cell_1rw
* cell instance $16774 m0 *1 3.525,90.09
X$16774 75 581 76 644 645 cell_1rw
* cell instance $16775 r0 *1 3.525,87.36
X$16775 75 322 76 644 645 cell_1rw
* cell instance $16776 r0 *1 3.525,90.09
X$16776 75 580 76 644 645 cell_1rw
* cell instance $16777 m0 *1 3.525,92.82
X$16777 75 583 76 644 645 cell_1rw
* cell instance $16778 r0 *1 3.525,92.82
X$16778 75 582 76 644 645 cell_1rw
* cell instance $16779 m0 *1 3.525,95.55
X$16779 75 584 76 644 645 cell_1rw
* cell instance $16780 r0 *1 3.525,95.55
X$16780 75 585 76 644 645 cell_1rw
* cell instance $16781 m0 *1 3.525,98.28
X$16781 75 586 76 644 645 cell_1rw
* cell instance $16782 m0 *1 3.525,101.01
X$16782 75 588 76 644 645 cell_1rw
* cell instance $16783 r0 *1 3.525,98.28
X$16783 75 587 76 644 645 cell_1rw
* cell instance $16784 r0 *1 3.525,101.01
X$16784 75 589 76 644 645 cell_1rw
* cell instance $16785 m0 *1 3.525,103.74
X$16785 75 590 76 644 645 cell_1rw
* cell instance $16786 m0 *1 3.525,106.47
X$16786 75 593 76 644 645 cell_1rw
* cell instance $16787 r0 *1 3.525,103.74
X$16787 75 591 76 644 645 cell_1rw
* cell instance $16788 r0 *1 3.525,106.47
X$16788 75 592 76 644 645 cell_1rw
* cell instance $16789 m0 *1 3.525,109.2
X$16789 75 594 76 644 645 cell_1rw
* cell instance $16790 r0 *1 3.525,109.2
X$16790 75 595 76 644 645 cell_1rw
* cell instance $16791 m0 *1 3.525,111.93
X$16791 75 597 76 644 645 cell_1rw
* cell instance $16792 r0 *1 3.525,111.93
X$16792 75 596 76 644 645 cell_1rw
* cell instance $16793 m0 *1 3.525,114.66
X$16793 75 598 76 644 645 cell_1rw
* cell instance $16794 r0 *1 3.525,114.66
X$16794 75 599 76 644 645 cell_1rw
* cell instance $16795 m0 *1 3.525,117.39
X$16795 75 600 76 644 645 cell_1rw
* cell instance $16796 r0 *1 3.525,117.39
X$16796 75 601 76 644 645 cell_1rw
* cell instance $16797 m0 *1 3.525,120.12
X$16797 75 602 76 644 645 cell_1rw
* cell instance $16798 r0 *1 3.525,120.12
X$16798 75 603 76 644 645 cell_1rw
* cell instance $16799 m0 *1 3.525,122.85
X$16799 75 604 76 644 645 cell_1rw
* cell instance $16800 r0 *1 3.525,122.85
X$16800 75 605 76 644 645 cell_1rw
* cell instance $16801 m0 *1 3.525,125.58
X$16801 75 606 76 644 645 cell_1rw
* cell instance $16802 m0 *1 3.525,128.31
X$16802 75 609 76 644 645 cell_1rw
* cell instance $16803 r0 *1 3.525,125.58
X$16803 75 607 76 644 645 cell_1rw
* cell instance $16804 m0 *1 3.525,131.04
X$16804 75 610 76 644 645 cell_1rw
* cell instance $16805 r0 *1 3.525,128.31
X$16805 75 608 76 644 645 cell_1rw
* cell instance $16806 r0 *1 3.525,131.04
X$16806 75 611 76 644 645 cell_1rw
* cell instance $16807 m0 *1 3.525,133.77
X$16807 75 612 76 644 645 cell_1rw
* cell instance $16808 r0 *1 3.525,133.77
X$16808 75 613 76 644 645 cell_1rw
* cell instance $16809 m0 *1 3.525,136.5
X$16809 75 615 76 644 645 cell_1rw
* cell instance $16810 r0 *1 3.525,136.5
X$16810 75 614 76 644 645 cell_1rw
* cell instance $16811 m0 *1 3.525,139.23
X$16811 75 617 76 644 645 cell_1rw
* cell instance $16812 m0 *1 3.525,141.96
X$16812 75 618 76 644 645 cell_1rw
* cell instance $16813 r0 *1 3.525,139.23
X$16813 75 616 76 644 645 cell_1rw
* cell instance $16814 r0 *1 3.525,141.96
X$16814 75 619 76 644 645 cell_1rw
* cell instance $16815 m0 *1 3.525,144.69
X$16815 75 620 76 644 645 cell_1rw
* cell instance $16816 r0 *1 3.525,144.69
X$16816 75 621 76 644 645 cell_1rw
* cell instance $16817 m0 *1 3.525,147.42
X$16817 75 622 76 644 645 cell_1rw
* cell instance $16818 r0 *1 3.525,147.42
X$16818 75 623 76 644 645 cell_1rw
* cell instance $16819 m0 *1 3.525,150.15
X$16819 75 624 76 644 645 cell_1rw
* cell instance $16820 r0 *1 3.525,150.15
X$16820 75 625 76 644 645 cell_1rw
* cell instance $16821 m0 *1 3.525,152.88
X$16821 75 626 76 644 645 cell_1rw
* cell instance $16822 r0 *1 3.525,152.88
X$16822 75 627 76 644 645 cell_1rw
* cell instance $16823 m0 *1 3.525,155.61
X$16823 75 628 76 644 645 cell_1rw
* cell instance $16824 m0 *1 3.525,158.34
X$16824 75 630 76 644 645 cell_1rw
* cell instance $16825 r0 *1 3.525,155.61
X$16825 75 629 76 644 645 cell_1rw
* cell instance $16826 r0 *1 3.525,158.34
X$16826 75 631 76 644 645 cell_1rw
* cell instance $16827 m0 *1 3.525,161.07
X$16827 75 632 76 644 645 cell_1rw
* cell instance $16828 r0 *1 3.525,161.07
X$16828 75 633 76 644 645 cell_1rw
* cell instance $16829 m0 *1 3.525,163.8
X$16829 75 634 76 644 645 cell_1rw
* cell instance $16830 r0 *1 3.525,163.8
X$16830 75 635 76 644 645 cell_1rw
* cell instance $16831 m0 *1 3.525,166.53
X$16831 75 637 76 644 645 cell_1rw
* cell instance $16832 r0 *1 3.525,166.53
X$16832 75 636 76 644 645 cell_1rw
* cell instance $16833 m0 *1 3.525,169.26
X$16833 75 639 76 644 645 cell_1rw
* cell instance $16834 r0 *1 3.525,169.26
X$16834 75 638 76 644 645 cell_1rw
* cell instance $16835 m0 *1 3.525,171.99
X$16835 75 640 76 644 645 cell_1rw
* cell instance $16836 r0 *1 3.525,171.99
X$16836 75 641 76 644 645 cell_1rw
* cell instance $16837 m0 *1 3.525,174.72
X$16837 75 642 76 644 645 cell_1rw
* cell instance $16838 r0 *1 3.525,174.72
X$16838 75 643 76 644 645 cell_1rw
* cell instance $16839 r0 *1 4.23,87.36
X$16839 77 322 78 644 645 cell_1rw
* cell instance $16840 m0 *1 4.23,90.09
X$16840 77 581 78 644 645 cell_1rw
* cell instance $16841 r0 *1 4.23,90.09
X$16841 77 580 78 644 645 cell_1rw
* cell instance $16842 m0 *1 4.23,92.82
X$16842 77 583 78 644 645 cell_1rw
* cell instance $16843 r0 *1 4.23,92.82
X$16843 77 582 78 644 645 cell_1rw
* cell instance $16844 m0 *1 4.23,95.55
X$16844 77 584 78 644 645 cell_1rw
* cell instance $16845 r0 *1 4.23,95.55
X$16845 77 585 78 644 645 cell_1rw
* cell instance $16846 m0 *1 4.23,98.28
X$16846 77 586 78 644 645 cell_1rw
* cell instance $16847 r0 *1 4.23,98.28
X$16847 77 587 78 644 645 cell_1rw
* cell instance $16848 m0 *1 4.23,101.01
X$16848 77 588 78 644 645 cell_1rw
* cell instance $16849 r0 *1 4.23,101.01
X$16849 77 589 78 644 645 cell_1rw
* cell instance $16850 m0 *1 4.23,103.74
X$16850 77 590 78 644 645 cell_1rw
* cell instance $16851 r0 *1 4.23,103.74
X$16851 77 591 78 644 645 cell_1rw
* cell instance $16852 m0 *1 4.23,106.47
X$16852 77 593 78 644 645 cell_1rw
* cell instance $16853 r0 *1 4.23,106.47
X$16853 77 592 78 644 645 cell_1rw
* cell instance $16854 m0 *1 4.23,109.2
X$16854 77 594 78 644 645 cell_1rw
* cell instance $16855 r0 *1 4.23,109.2
X$16855 77 595 78 644 645 cell_1rw
* cell instance $16856 m0 *1 4.23,111.93
X$16856 77 597 78 644 645 cell_1rw
* cell instance $16857 r0 *1 4.23,111.93
X$16857 77 596 78 644 645 cell_1rw
* cell instance $16858 m0 *1 4.23,114.66
X$16858 77 598 78 644 645 cell_1rw
* cell instance $16859 r0 *1 4.23,114.66
X$16859 77 599 78 644 645 cell_1rw
* cell instance $16860 m0 *1 4.23,117.39
X$16860 77 600 78 644 645 cell_1rw
* cell instance $16861 r0 *1 4.23,117.39
X$16861 77 601 78 644 645 cell_1rw
* cell instance $16862 m0 *1 4.23,120.12
X$16862 77 602 78 644 645 cell_1rw
* cell instance $16863 r0 *1 4.23,120.12
X$16863 77 603 78 644 645 cell_1rw
* cell instance $16864 m0 *1 4.23,122.85
X$16864 77 604 78 644 645 cell_1rw
* cell instance $16865 r0 *1 4.23,122.85
X$16865 77 605 78 644 645 cell_1rw
* cell instance $16866 m0 *1 4.23,125.58
X$16866 77 606 78 644 645 cell_1rw
* cell instance $16867 r0 *1 4.23,125.58
X$16867 77 607 78 644 645 cell_1rw
* cell instance $16868 m0 *1 4.23,128.31
X$16868 77 609 78 644 645 cell_1rw
* cell instance $16869 r0 *1 4.23,128.31
X$16869 77 608 78 644 645 cell_1rw
* cell instance $16870 m0 *1 4.23,131.04
X$16870 77 610 78 644 645 cell_1rw
* cell instance $16871 m0 *1 4.23,133.77
X$16871 77 612 78 644 645 cell_1rw
* cell instance $16872 r0 *1 4.23,131.04
X$16872 77 611 78 644 645 cell_1rw
* cell instance $16873 r0 *1 4.23,133.77
X$16873 77 613 78 644 645 cell_1rw
* cell instance $16874 m0 *1 4.23,136.5
X$16874 77 615 78 644 645 cell_1rw
* cell instance $16875 m0 *1 4.23,139.23
X$16875 77 617 78 644 645 cell_1rw
* cell instance $16876 r0 *1 4.23,136.5
X$16876 77 614 78 644 645 cell_1rw
* cell instance $16877 r0 *1 4.23,139.23
X$16877 77 616 78 644 645 cell_1rw
* cell instance $16878 m0 *1 4.23,141.96
X$16878 77 618 78 644 645 cell_1rw
* cell instance $16879 r0 *1 4.23,141.96
X$16879 77 619 78 644 645 cell_1rw
* cell instance $16880 m0 *1 4.23,144.69
X$16880 77 620 78 644 645 cell_1rw
* cell instance $16881 r0 *1 4.23,144.69
X$16881 77 621 78 644 645 cell_1rw
* cell instance $16882 m0 *1 4.23,147.42
X$16882 77 622 78 644 645 cell_1rw
* cell instance $16883 r0 *1 4.23,147.42
X$16883 77 623 78 644 645 cell_1rw
* cell instance $16884 m0 *1 4.23,150.15
X$16884 77 624 78 644 645 cell_1rw
* cell instance $16885 r0 *1 4.23,150.15
X$16885 77 625 78 644 645 cell_1rw
* cell instance $16886 m0 *1 4.23,152.88
X$16886 77 626 78 644 645 cell_1rw
* cell instance $16887 r0 *1 4.23,152.88
X$16887 77 627 78 644 645 cell_1rw
* cell instance $16888 m0 *1 4.23,155.61
X$16888 77 628 78 644 645 cell_1rw
* cell instance $16889 r0 *1 4.23,155.61
X$16889 77 629 78 644 645 cell_1rw
* cell instance $16890 m0 *1 4.23,158.34
X$16890 77 630 78 644 645 cell_1rw
* cell instance $16891 r0 *1 4.23,158.34
X$16891 77 631 78 644 645 cell_1rw
* cell instance $16892 m0 *1 4.23,161.07
X$16892 77 632 78 644 645 cell_1rw
* cell instance $16893 r0 *1 4.23,161.07
X$16893 77 633 78 644 645 cell_1rw
* cell instance $16894 m0 *1 4.23,163.8
X$16894 77 634 78 644 645 cell_1rw
* cell instance $16895 r0 *1 4.23,163.8
X$16895 77 635 78 644 645 cell_1rw
* cell instance $16896 m0 *1 4.23,166.53
X$16896 77 637 78 644 645 cell_1rw
* cell instance $16897 m0 *1 4.23,169.26
X$16897 77 639 78 644 645 cell_1rw
* cell instance $16898 r0 *1 4.23,166.53
X$16898 77 636 78 644 645 cell_1rw
* cell instance $16899 r0 *1 4.23,169.26
X$16899 77 638 78 644 645 cell_1rw
* cell instance $16900 m0 *1 4.23,171.99
X$16900 77 640 78 644 645 cell_1rw
* cell instance $16901 r0 *1 4.23,171.99
X$16901 77 641 78 644 645 cell_1rw
* cell instance $16902 m0 *1 4.23,174.72
X$16902 77 642 78 644 645 cell_1rw
* cell instance $16903 r0 *1 4.23,174.72
X$16903 77 643 78 644 645 cell_1rw
* cell instance $16904 r0 *1 4.935,87.36
X$16904 79 322 80 644 645 cell_1rw
* cell instance $16905 m0 *1 4.935,90.09
X$16905 79 581 80 644 645 cell_1rw
* cell instance $16906 r0 *1 4.935,90.09
X$16906 79 580 80 644 645 cell_1rw
* cell instance $16907 m0 *1 4.935,92.82
X$16907 79 583 80 644 645 cell_1rw
* cell instance $16908 r0 *1 4.935,92.82
X$16908 79 582 80 644 645 cell_1rw
* cell instance $16909 m0 *1 4.935,95.55
X$16909 79 584 80 644 645 cell_1rw
* cell instance $16910 r0 *1 4.935,95.55
X$16910 79 585 80 644 645 cell_1rw
* cell instance $16911 m0 *1 4.935,98.28
X$16911 79 586 80 644 645 cell_1rw
* cell instance $16912 r0 *1 4.935,98.28
X$16912 79 587 80 644 645 cell_1rw
* cell instance $16913 m0 *1 4.935,101.01
X$16913 79 588 80 644 645 cell_1rw
* cell instance $16914 r0 *1 4.935,101.01
X$16914 79 589 80 644 645 cell_1rw
* cell instance $16915 m0 *1 4.935,103.74
X$16915 79 590 80 644 645 cell_1rw
* cell instance $16916 r0 *1 4.935,103.74
X$16916 79 591 80 644 645 cell_1rw
* cell instance $16917 m0 *1 4.935,106.47
X$16917 79 593 80 644 645 cell_1rw
* cell instance $16918 r0 *1 4.935,106.47
X$16918 79 592 80 644 645 cell_1rw
* cell instance $16919 m0 *1 4.935,109.2
X$16919 79 594 80 644 645 cell_1rw
* cell instance $16920 r0 *1 4.935,109.2
X$16920 79 595 80 644 645 cell_1rw
* cell instance $16921 m0 *1 4.935,111.93
X$16921 79 597 80 644 645 cell_1rw
* cell instance $16922 r0 *1 4.935,111.93
X$16922 79 596 80 644 645 cell_1rw
* cell instance $16923 m0 *1 4.935,114.66
X$16923 79 598 80 644 645 cell_1rw
* cell instance $16924 r0 *1 4.935,114.66
X$16924 79 599 80 644 645 cell_1rw
* cell instance $16925 m0 *1 4.935,117.39
X$16925 79 600 80 644 645 cell_1rw
* cell instance $16926 r0 *1 4.935,117.39
X$16926 79 601 80 644 645 cell_1rw
* cell instance $16927 m0 *1 4.935,120.12
X$16927 79 602 80 644 645 cell_1rw
* cell instance $16928 m0 *1 4.935,122.85
X$16928 79 604 80 644 645 cell_1rw
* cell instance $16929 r0 *1 4.935,120.12
X$16929 79 603 80 644 645 cell_1rw
* cell instance $16930 r0 *1 4.935,122.85
X$16930 79 605 80 644 645 cell_1rw
* cell instance $16931 m0 *1 4.935,125.58
X$16931 79 606 80 644 645 cell_1rw
* cell instance $16932 r0 *1 4.935,125.58
X$16932 79 607 80 644 645 cell_1rw
* cell instance $16933 m0 *1 4.935,128.31
X$16933 79 609 80 644 645 cell_1rw
* cell instance $16934 r0 *1 4.935,128.31
X$16934 79 608 80 644 645 cell_1rw
* cell instance $16935 m0 *1 4.935,131.04
X$16935 79 610 80 644 645 cell_1rw
* cell instance $16936 r0 *1 4.935,131.04
X$16936 79 611 80 644 645 cell_1rw
* cell instance $16937 m0 *1 4.935,133.77
X$16937 79 612 80 644 645 cell_1rw
* cell instance $16938 r0 *1 4.935,133.77
X$16938 79 613 80 644 645 cell_1rw
* cell instance $16939 m0 *1 4.935,136.5
X$16939 79 615 80 644 645 cell_1rw
* cell instance $16940 r0 *1 4.935,136.5
X$16940 79 614 80 644 645 cell_1rw
* cell instance $16941 m0 *1 4.935,139.23
X$16941 79 617 80 644 645 cell_1rw
* cell instance $16942 r0 *1 4.935,139.23
X$16942 79 616 80 644 645 cell_1rw
* cell instance $16943 m0 *1 4.935,141.96
X$16943 79 618 80 644 645 cell_1rw
* cell instance $16944 r0 *1 4.935,141.96
X$16944 79 619 80 644 645 cell_1rw
* cell instance $16945 m0 *1 4.935,144.69
X$16945 79 620 80 644 645 cell_1rw
* cell instance $16946 r0 *1 4.935,144.69
X$16946 79 621 80 644 645 cell_1rw
* cell instance $16947 m0 *1 4.935,147.42
X$16947 79 622 80 644 645 cell_1rw
* cell instance $16948 r0 *1 4.935,147.42
X$16948 79 623 80 644 645 cell_1rw
* cell instance $16949 m0 *1 4.935,150.15
X$16949 79 624 80 644 645 cell_1rw
* cell instance $16950 r0 *1 4.935,150.15
X$16950 79 625 80 644 645 cell_1rw
* cell instance $16951 m0 *1 4.935,152.88
X$16951 79 626 80 644 645 cell_1rw
* cell instance $16952 r0 *1 4.935,152.88
X$16952 79 627 80 644 645 cell_1rw
* cell instance $16953 m0 *1 4.935,155.61
X$16953 79 628 80 644 645 cell_1rw
* cell instance $16954 r0 *1 4.935,155.61
X$16954 79 629 80 644 645 cell_1rw
* cell instance $16955 m0 *1 4.935,158.34
X$16955 79 630 80 644 645 cell_1rw
* cell instance $16956 r0 *1 4.935,158.34
X$16956 79 631 80 644 645 cell_1rw
* cell instance $16957 m0 *1 4.935,161.07
X$16957 79 632 80 644 645 cell_1rw
* cell instance $16958 r0 *1 4.935,161.07
X$16958 79 633 80 644 645 cell_1rw
* cell instance $16959 m0 *1 4.935,163.8
X$16959 79 634 80 644 645 cell_1rw
* cell instance $16960 r0 *1 4.935,163.8
X$16960 79 635 80 644 645 cell_1rw
* cell instance $16961 m0 *1 4.935,166.53
X$16961 79 637 80 644 645 cell_1rw
* cell instance $16962 r0 *1 4.935,166.53
X$16962 79 636 80 644 645 cell_1rw
* cell instance $16963 m0 *1 4.935,169.26
X$16963 79 639 80 644 645 cell_1rw
* cell instance $16964 r0 *1 4.935,169.26
X$16964 79 638 80 644 645 cell_1rw
* cell instance $16965 m0 *1 4.935,171.99
X$16965 79 640 80 644 645 cell_1rw
* cell instance $16966 r0 *1 4.935,171.99
X$16966 79 641 80 644 645 cell_1rw
* cell instance $16967 m0 *1 4.935,174.72
X$16967 79 642 80 644 645 cell_1rw
* cell instance $16968 r0 *1 4.935,174.72
X$16968 79 643 80 644 645 cell_1rw
* cell instance $16969 r0 *1 5.64,87.36
X$16969 81 322 82 644 645 cell_1rw
* cell instance $16970 m0 *1 5.64,90.09
X$16970 81 581 82 644 645 cell_1rw
* cell instance $16971 m0 *1 5.64,92.82
X$16971 81 583 82 644 645 cell_1rw
* cell instance $16972 r0 *1 5.64,90.09
X$16972 81 580 82 644 645 cell_1rw
* cell instance $16973 r0 *1 5.64,92.82
X$16973 81 582 82 644 645 cell_1rw
* cell instance $16974 m0 *1 5.64,95.55
X$16974 81 584 82 644 645 cell_1rw
* cell instance $16975 r0 *1 5.64,95.55
X$16975 81 585 82 644 645 cell_1rw
* cell instance $16976 m0 *1 5.64,98.28
X$16976 81 586 82 644 645 cell_1rw
* cell instance $16977 r0 *1 5.64,98.28
X$16977 81 587 82 644 645 cell_1rw
* cell instance $16978 m0 *1 5.64,101.01
X$16978 81 588 82 644 645 cell_1rw
* cell instance $16979 m0 *1 5.64,103.74
X$16979 81 590 82 644 645 cell_1rw
* cell instance $16980 r0 *1 5.64,101.01
X$16980 81 589 82 644 645 cell_1rw
* cell instance $16981 r0 *1 5.64,103.74
X$16981 81 591 82 644 645 cell_1rw
* cell instance $16982 m0 *1 5.64,106.47
X$16982 81 593 82 644 645 cell_1rw
* cell instance $16983 r0 *1 5.64,106.47
X$16983 81 592 82 644 645 cell_1rw
* cell instance $16984 m0 *1 5.64,109.2
X$16984 81 594 82 644 645 cell_1rw
* cell instance $16985 r0 *1 5.64,109.2
X$16985 81 595 82 644 645 cell_1rw
* cell instance $16986 m0 *1 5.64,111.93
X$16986 81 597 82 644 645 cell_1rw
* cell instance $16987 m0 *1 5.64,114.66
X$16987 81 598 82 644 645 cell_1rw
* cell instance $16988 r0 *1 5.64,111.93
X$16988 81 596 82 644 645 cell_1rw
* cell instance $16989 r0 *1 5.64,114.66
X$16989 81 599 82 644 645 cell_1rw
* cell instance $16990 m0 *1 5.64,117.39
X$16990 81 600 82 644 645 cell_1rw
* cell instance $16991 m0 *1 5.64,120.12
X$16991 81 602 82 644 645 cell_1rw
* cell instance $16992 r0 *1 5.64,117.39
X$16992 81 601 82 644 645 cell_1rw
* cell instance $16993 r0 *1 5.64,120.12
X$16993 81 603 82 644 645 cell_1rw
* cell instance $16994 m0 *1 5.64,122.85
X$16994 81 604 82 644 645 cell_1rw
* cell instance $16995 r0 *1 5.64,122.85
X$16995 81 605 82 644 645 cell_1rw
* cell instance $16996 m0 *1 5.64,125.58
X$16996 81 606 82 644 645 cell_1rw
* cell instance $16997 r0 *1 5.64,125.58
X$16997 81 607 82 644 645 cell_1rw
* cell instance $16998 m0 *1 5.64,128.31
X$16998 81 609 82 644 645 cell_1rw
* cell instance $16999 r0 *1 5.64,128.31
X$16999 81 608 82 644 645 cell_1rw
* cell instance $17000 m0 *1 5.64,131.04
X$17000 81 610 82 644 645 cell_1rw
* cell instance $17001 r0 *1 5.64,131.04
X$17001 81 611 82 644 645 cell_1rw
* cell instance $17002 m0 *1 5.64,133.77
X$17002 81 612 82 644 645 cell_1rw
* cell instance $17003 r0 *1 5.64,133.77
X$17003 81 613 82 644 645 cell_1rw
* cell instance $17004 m0 *1 5.64,136.5
X$17004 81 615 82 644 645 cell_1rw
* cell instance $17005 r0 *1 5.64,136.5
X$17005 81 614 82 644 645 cell_1rw
* cell instance $17006 m0 *1 5.64,139.23
X$17006 81 617 82 644 645 cell_1rw
* cell instance $17007 r0 *1 5.64,139.23
X$17007 81 616 82 644 645 cell_1rw
* cell instance $17008 m0 *1 5.64,141.96
X$17008 81 618 82 644 645 cell_1rw
* cell instance $17009 r0 *1 5.64,141.96
X$17009 81 619 82 644 645 cell_1rw
* cell instance $17010 m0 *1 5.64,144.69
X$17010 81 620 82 644 645 cell_1rw
* cell instance $17011 r0 *1 5.64,144.69
X$17011 81 621 82 644 645 cell_1rw
* cell instance $17012 m0 *1 5.64,147.42
X$17012 81 622 82 644 645 cell_1rw
* cell instance $17013 r0 *1 5.64,147.42
X$17013 81 623 82 644 645 cell_1rw
* cell instance $17014 m0 *1 5.64,150.15
X$17014 81 624 82 644 645 cell_1rw
* cell instance $17015 r0 *1 5.64,150.15
X$17015 81 625 82 644 645 cell_1rw
* cell instance $17016 m0 *1 5.64,152.88
X$17016 81 626 82 644 645 cell_1rw
* cell instance $17017 r0 *1 5.64,152.88
X$17017 81 627 82 644 645 cell_1rw
* cell instance $17018 m0 *1 5.64,155.61
X$17018 81 628 82 644 645 cell_1rw
* cell instance $17019 r0 *1 5.64,155.61
X$17019 81 629 82 644 645 cell_1rw
* cell instance $17020 m0 *1 5.64,158.34
X$17020 81 630 82 644 645 cell_1rw
* cell instance $17021 r0 *1 5.64,158.34
X$17021 81 631 82 644 645 cell_1rw
* cell instance $17022 m0 *1 5.64,161.07
X$17022 81 632 82 644 645 cell_1rw
* cell instance $17023 r0 *1 5.64,161.07
X$17023 81 633 82 644 645 cell_1rw
* cell instance $17024 m0 *1 5.64,163.8
X$17024 81 634 82 644 645 cell_1rw
* cell instance $17025 r0 *1 5.64,163.8
X$17025 81 635 82 644 645 cell_1rw
* cell instance $17026 m0 *1 5.64,166.53
X$17026 81 637 82 644 645 cell_1rw
* cell instance $17027 r0 *1 5.64,166.53
X$17027 81 636 82 644 645 cell_1rw
* cell instance $17028 m0 *1 5.64,169.26
X$17028 81 639 82 644 645 cell_1rw
* cell instance $17029 r0 *1 5.64,169.26
X$17029 81 638 82 644 645 cell_1rw
* cell instance $17030 m0 *1 5.64,171.99
X$17030 81 640 82 644 645 cell_1rw
* cell instance $17031 r0 *1 5.64,171.99
X$17031 81 641 82 644 645 cell_1rw
* cell instance $17032 m0 *1 5.64,174.72
X$17032 81 642 82 644 645 cell_1rw
* cell instance $17033 r0 *1 5.64,174.72
X$17033 81 643 82 644 645 cell_1rw
* cell instance $17034 m0 *1 6.345,90.09
X$17034 83 581 84 644 645 cell_1rw
* cell instance $17035 r0 *1 6.345,87.36
X$17035 83 322 84 644 645 cell_1rw
* cell instance $17036 m0 *1 6.345,92.82
X$17036 83 583 84 644 645 cell_1rw
* cell instance $17037 r0 *1 6.345,90.09
X$17037 83 580 84 644 645 cell_1rw
* cell instance $17038 m0 *1 6.345,95.55
X$17038 83 584 84 644 645 cell_1rw
* cell instance $17039 r0 *1 6.345,92.82
X$17039 83 582 84 644 645 cell_1rw
* cell instance $17040 r0 *1 6.345,95.55
X$17040 83 585 84 644 645 cell_1rw
* cell instance $17041 m0 *1 6.345,98.28
X$17041 83 586 84 644 645 cell_1rw
* cell instance $17042 r0 *1 6.345,98.28
X$17042 83 587 84 644 645 cell_1rw
* cell instance $17043 m0 *1 6.345,101.01
X$17043 83 588 84 644 645 cell_1rw
* cell instance $17044 r0 *1 6.345,101.01
X$17044 83 589 84 644 645 cell_1rw
* cell instance $17045 m0 *1 6.345,103.74
X$17045 83 590 84 644 645 cell_1rw
* cell instance $17046 m0 *1 6.345,106.47
X$17046 83 593 84 644 645 cell_1rw
* cell instance $17047 r0 *1 6.345,103.74
X$17047 83 591 84 644 645 cell_1rw
* cell instance $17048 r0 *1 6.345,106.47
X$17048 83 592 84 644 645 cell_1rw
* cell instance $17049 m0 *1 6.345,109.2
X$17049 83 594 84 644 645 cell_1rw
* cell instance $17050 r0 *1 6.345,109.2
X$17050 83 595 84 644 645 cell_1rw
* cell instance $17051 m0 *1 6.345,111.93
X$17051 83 597 84 644 645 cell_1rw
* cell instance $17052 r0 *1 6.345,111.93
X$17052 83 596 84 644 645 cell_1rw
* cell instance $17053 m0 *1 6.345,114.66
X$17053 83 598 84 644 645 cell_1rw
* cell instance $17054 r0 *1 6.345,114.66
X$17054 83 599 84 644 645 cell_1rw
* cell instance $17055 m0 *1 6.345,117.39
X$17055 83 600 84 644 645 cell_1rw
* cell instance $17056 r0 *1 6.345,117.39
X$17056 83 601 84 644 645 cell_1rw
* cell instance $17057 m0 *1 6.345,120.12
X$17057 83 602 84 644 645 cell_1rw
* cell instance $17058 r0 *1 6.345,120.12
X$17058 83 603 84 644 645 cell_1rw
* cell instance $17059 m0 *1 6.345,122.85
X$17059 83 604 84 644 645 cell_1rw
* cell instance $17060 r0 *1 6.345,122.85
X$17060 83 605 84 644 645 cell_1rw
* cell instance $17061 m0 *1 6.345,125.58
X$17061 83 606 84 644 645 cell_1rw
* cell instance $17062 r0 *1 6.345,125.58
X$17062 83 607 84 644 645 cell_1rw
* cell instance $17063 m0 *1 6.345,128.31
X$17063 83 609 84 644 645 cell_1rw
* cell instance $17064 r0 *1 6.345,128.31
X$17064 83 608 84 644 645 cell_1rw
* cell instance $17065 m0 *1 6.345,131.04
X$17065 83 610 84 644 645 cell_1rw
* cell instance $17066 r0 *1 6.345,131.04
X$17066 83 611 84 644 645 cell_1rw
* cell instance $17067 m0 *1 6.345,133.77
X$17067 83 612 84 644 645 cell_1rw
* cell instance $17068 r0 *1 6.345,133.77
X$17068 83 613 84 644 645 cell_1rw
* cell instance $17069 m0 *1 6.345,136.5
X$17069 83 615 84 644 645 cell_1rw
* cell instance $17070 m0 *1 6.345,139.23
X$17070 83 617 84 644 645 cell_1rw
* cell instance $17071 r0 *1 6.345,136.5
X$17071 83 614 84 644 645 cell_1rw
* cell instance $17072 r0 *1 6.345,139.23
X$17072 83 616 84 644 645 cell_1rw
* cell instance $17073 m0 *1 6.345,141.96
X$17073 83 618 84 644 645 cell_1rw
* cell instance $17074 m0 *1 6.345,144.69
X$17074 83 620 84 644 645 cell_1rw
* cell instance $17075 r0 *1 6.345,141.96
X$17075 83 619 84 644 645 cell_1rw
* cell instance $17076 m0 *1 6.345,147.42
X$17076 83 622 84 644 645 cell_1rw
* cell instance $17077 r0 *1 6.345,144.69
X$17077 83 621 84 644 645 cell_1rw
* cell instance $17078 r0 *1 6.345,147.42
X$17078 83 623 84 644 645 cell_1rw
* cell instance $17079 m0 *1 6.345,150.15
X$17079 83 624 84 644 645 cell_1rw
* cell instance $17080 r0 *1 6.345,150.15
X$17080 83 625 84 644 645 cell_1rw
* cell instance $17081 m0 *1 6.345,152.88
X$17081 83 626 84 644 645 cell_1rw
* cell instance $17082 r0 *1 6.345,152.88
X$17082 83 627 84 644 645 cell_1rw
* cell instance $17083 m0 *1 6.345,155.61
X$17083 83 628 84 644 645 cell_1rw
* cell instance $17084 m0 *1 6.345,158.34
X$17084 83 630 84 644 645 cell_1rw
* cell instance $17085 r0 *1 6.345,155.61
X$17085 83 629 84 644 645 cell_1rw
* cell instance $17086 r0 *1 6.345,158.34
X$17086 83 631 84 644 645 cell_1rw
* cell instance $17087 m0 *1 6.345,161.07
X$17087 83 632 84 644 645 cell_1rw
* cell instance $17088 r0 *1 6.345,161.07
X$17088 83 633 84 644 645 cell_1rw
* cell instance $17089 m0 *1 6.345,163.8
X$17089 83 634 84 644 645 cell_1rw
* cell instance $17090 r0 *1 6.345,163.8
X$17090 83 635 84 644 645 cell_1rw
* cell instance $17091 m0 *1 6.345,166.53
X$17091 83 637 84 644 645 cell_1rw
* cell instance $17092 r0 *1 6.345,166.53
X$17092 83 636 84 644 645 cell_1rw
* cell instance $17093 m0 *1 6.345,169.26
X$17093 83 639 84 644 645 cell_1rw
* cell instance $17094 r0 *1 6.345,169.26
X$17094 83 638 84 644 645 cell_1rw
* cell instance $17095 m0 *1 6.345,171.99
X$17095 83 640 84 644 645 cell_1rw
* cell instance $17096 r0 *1 6.345,171.99
X$17096 83 641 84 644 645 cell_1rw
* cell instance $17097 m0 *1 6.345,174.72
X$17097 83 642 84 644 645 cell_1rw
* cell instance $17098 r0 *1 6.345,174.72
X$17098 83 643 84 644 645 cell_1rw
* cell instance $17099 r0 *1 7.05,87.36
X$17099 85 322 86 644 645 cell_1rw
* cell instance $17100 m0 *1 7.05,90.09
X$17100 85 581 86 644 645 cell_1rw
* cell instance $17101 r0 *1 7.05,90.09
X$17101 85 580 86 644 645 cell_1rw
* cell instance $17102 m0 *1 7.05,92.82
X$17102 85 583 86 644 645 cell_1rw
* cell instance $17103 r0 *1 7.05,92.82
X$17103 85 582 86 644 645 cell_1rw
* cell instance $17104 m0 *1 7.05,95.55
X$17104 85 584 86 644 645 cell_1rw
* cell instance $17105 r0 *1 7.05,95.55
X$17105 85 585 86 644 645 cell_1rw
* cell instance $17106 m0 *1 7.05,98.28
X$17106 85 586 86 644 645 cell_1rw
* cell instance $17107 m0 *1 7.05,101.01
X$17107 85 588 86 644 645 cell_1rw
* cell instance $17108 r0 *1 7.05,98.28
X$17108 85 587 86 644 645 cell_1rw
* cell instance $17109 r0 *1 7.05,101.01
X$17109 85 589 86 644 645 cell_1rw
* cell instance $17110 m0 *1 7.05,103.74
X$17110 85 590 86 644 645 cell_1rw
* cell instance $17111 r0 *1 7.05,103.74
X$17111 85 591 86 644 645 cell_1rw
* cell instance $17112 m0 *1 7.05,106.47
X$17112 85 593 86 644 645 cell_1rw
* cell instance $17113 r0 *1 7.05,106.47
X$17113 85 592 86 644 645 cell_1rw
* cell instance $17114 m0 *1 7.05,109.2
X$17114 85 594 86 644 645 cell_1rw
* cell instance $17115 m0 *1 7.05,111.93
X$17115 85 597 86 644 645 cell_1rw
* cell instance $17116 r0 *1 7.05,109.2
X$17116 85 595 86 644 645 cell_1rw
* cell instance $17117 r0 *1 7.05,111.93
X$17117 85 596 86 644 645 cell_1rw
* cell instance $17118 m0 *1 7.05,114.66
X$17118 85 598 86 644 645 cell_1rw
* cell instance $17119 r0 *1 7.05,114.66
X$17119 85 599 86 644 645 cell_1rw
* cell instance $17120 m0 *1 7.05,117.39
X$17120 85 600 86 644 645 cell_1rw
* cell instance $17121 m0 *1 7.05,120.12
X$17121 85 602 86 644 645 cell_1rw
* cell instance $17122 r0 *1 7.05,117.39
X$17122 85 601 86 644 645 cell_1rw
* cell instance $17123 r0 *1 7.05,120.12
X$17123 85 603 86 644 645 cell_1rw
* cell instance $17124 m0 *1 7.05,122.85
X$17124 85 604 86 644 645 cell_1rw
* cell instance $17125 r0 *1 7.05,122.85
X$17125 85 605 86 644 645 cell_1rw
* cell instance $17126 m0 *1 7.05,125.58
X$17126 85 606 86 644 645 cell_1rw
* cell instance $17127 r0 *1 7.05,125.58
X$17127 85 607 86 644 645 cell_1rw
* cell instance $17128 m0 *1 7.05,128.31
X$17128 85 609 86 644 645 cell_1rw
* cell instance $17129 r0 *1 7.05,128.31
X$17129 85 608 86 644 645 cell_1rw
* cell instance $17130 m0 *1 7.05,131.04
X$17130 85 610 86 644 645 cell_1rw
* cell instance $17131 r0 *1 7.05,131.04
X$17131 85 611 86 644 645 cell_1rw
* cell instance $17132 m0 *1 7.05,133.77
X$17132 85 612 86 644 645 cell_1rw
* cell instance $17133 r0 *1 7.05,133.77
X$17133 85 613 86 644 645 cell_1rw
* cell instance $17134 m0 *1 7.05,136.5
X$17134 85 615 86 644 645 cell_1rw
* cell instance $17135 m0 *1 7.05,139.23
X$17135 85 617 86 644 645 cell_1rw
* cell instance $17136 r0 *1 7.05,136.5
X$17136 85 614 86 644 645 cell_1rw
* cell instance $17137 r0 *1 7.05,139.23
X$17137 85 616 86 644 645 cell_1rw
* cell instance $17138 m0 *1 7.05,141.96
X$17138 85 618 86 644 645 cell_1rw
* cell instance $17139 r0 *1 7.05,141.96
X$17139 85 619 86 644 645 cell_1rw
* cell instance $17140 m0 *1 7.05,144.69
X$17140 85 620 86 644 645 cell_1rw
* cell instance $17141 r0 *1 7.05,144.69
X$17141 85 621 86 644 645 cell_1rw
* cell instance $17142 m0 *1 7.05,147.42
X$17142 85 622 86 644 645 cell_1rw
* cell instance $17143 r0 *1 7.05,147.42
X$17143 85 623 86 644 645 cell_1rw
* cell instance $17144 m0 *1 7.05,150.15
X$17144 85 624 86 644 645 cell_1rw
* cell instance $17145 r0 *1 7.05,150.15
X$17145 85 625 86 644 645 cell_1rw
* cell instance $17146 m0 *1 7.05,152.88
X$17146 85 626 86 644 645 cell_1rw
* cell instance $17147 r0 *1 7.05,152.88
X$17147 85 627 86 644 645 cell_1rw
* cell instance $17148 m0 *1 7.05,155.61
X$17148 85 628 86 644 645 cell_1rw
* cell instance $17149 m0 *1 7.05,158.34
X$17149 85 630 86 644 645 cell_1rw
* cell instance $17150 r0 *1 7.05,155.61
X$17150 85 629 86 644 645 cell_1rw
* cell instance $17151 m0 *1 7.05,161.07
X$17151 85 632 86 644 645 cell_1rw
* cell instance $17152 r0 *1 7.05,158.34
X$17152 85 631 86 644 645 cell_1rw
* cell instance $17153 r0 *1 7.05,161.07
X$17153 85 633 86 644 645 cell_1rw
* cell instance $17154 m0 *1 7.05,163.8
X$17154 85 634 86 644 645 cell_1rw
* cell instance $17155 r0 *1 7.05,163.8
X$17155 85 635 86 644 645 cell_1rw
* cell instance $17156 m0 *1 7.05,166.53
X$17156 85 637 86 644 645 cell_1rw
* cell instance $17157 m0 *1 7.05,169.26
X$17157 85 639 86 644 645 cell_1rw
* cell instance $17158 r0 *1 7.05,166.53
X$17158 85 636 86 644 645 cell_1rw
* cell instance $17159 r0 *1 7.05,169.26
X$17159 85 638 86 644 645 cell_1rw
* cell instance $17160 m0 *1 7.05,171.99
X$17160 85 640 86 644 645 cell_1rw
* cell instance $17161 r0 *1 7.05,171.99
X$17161 85 641 86 644 645 cell_1rw
* cell instance $17162 m0 *1 7.05,174.72
X$17162 85 642 86 644 645 cell_1rw
* cell instance $17163 r0 *1 7.05,174.72
X$17163 85 643 86 644 645 cell_1rw
* cell instance $17164 r0 *1 7.755,87.36
X$17164 87 322 88 644 645 cell_1rw
* cell instance $17165 m0 *1 7.755,90.09
X$17165 87 581 88 644 645 cell_1rw
* cell instance $17166 r0 *1 7.755,90.09
X$17166 87 580 88 644 645 cell_1rw
* cell instance $17167 m0 *1 7.755,92.82
X$17167 87 583 88 644 645 cell_1rw
* cell instance $17168 m0 *1 7.755,95.55
X$17168 87 584 88 644 645 cell_1rw
* cell instance $17169 r0 *1 7.755,92.82
X$17169 87 582 88 644 645 cell_1rw
* cell instance $17170 r0 *1 7.755,95.55
X$17170 87 585 88 644 645 cell_1rw
* cell instance $17171 m0 *1 7.755,98.28
X$17171 87 586 88 644 645 cell_1rw
* cell instance $17172 r0 *1 7.755,98.28
X$17172 87 587 88 644 645 cell_1rw
* cell instance $17173 m0 *1 7.755,101.01
X$17173 87 588 88 644 645 cell_1rw
* cell instance $17174 r0 *1 7.755,101.01
X$17174 87 589 88 644 645 cell_1rw
* cell instance $17175 m0 *1 7.755,103.74
X$17175 87 590 88 644 645 cell_1rw
* cell instance $17176 r0 *1 7.755,103.74
X$17176 87 591 88 644 645 cell_1rw
* cell instance $17177 m0 *1 7.755,106.47
X$17177 87 593 88 644 645 cell_1rw
* cell instance $17178 r0 *1 7.755,106.47
X$17178 87 592 88 644 645 cell_1rw
* cell instance $17179 m0 *1 7.755,109.2
X$17179 87 594 88 644 645 cell_1rw
* cell instance $17180 r0 *1 7.755,109.2
X$17180 87 595 88 644 645 cell_1rw
* cell instance $17181 m0 *1 7.755,111.93
X$17181 87 597 88 644 645 cell_1rw
* cell instance $17182 r0 *1 7.755,111.93
X$17182 87 596 88 644 645 cell_1rw
* cell instance $17183 m0 *1 7.755,114.66
X$17183 87 598 88 644 645 cell_1rw
* cell instance $17184 r0 *1 7.755,114.66
X$17184 87 599 88 644 645 cell_1rw
* cell instance $17185 m0 *1 7.755,117.39
X$17185 87 600 88 644 645 cell_1rw
* cell instance $17186 r0 *1 7.755,117.39
X$17186 87 601 88 644 645 cell_1rw
* cell instance $17187 m0 *1 7.755,120.12
X$17187 87 602 88 644 645 cell_1rw
* cell instance $17188 r0 *1 7.755,120.12
X$17188 87 603 88 644 645 cell_1rw
* cell instance $17189 m0 *1 7.755,122.85
X$17189 87 604 88 644 645 cell_1rw
* cell instance $17190 r0 *1 7.755,122.85
X$17190 87 605 88 644 645 cell_1rw
* cell instance $17191 m0 *1 7.755,125.58
X$17191 87 606 88 644 645 cell_1rw
* cell instance $17192 r0 *1 7.755,125.58
X$17192 87 607 88 644 645 cell_1rw
* cell instance $17193 m0 *1 7.755,128.31
X$17193 87 609 88 644 645 cell_1rw
* cell instance $17194 r0 *1 7.755,128.31
X$17194 87 608 88 644 645 cell_1rw
* cell instance $17195 m0 *1 7.755,131.04
X$17195 87 610 88 644 645 cell_1rw
* cell instance $17196 m0 *1 7.755,133.77
X$17196 87 612 88 644 645 cell_1rw
* cell instance $17197 r0 *1 7.755,131.04
X$17197 87 611 88 644 645 cell_1rw
* cell instance $17198 r0 *1 7.755,133.77
X$17198 87 613 88 644 645 cell_1rw
* cell instance $17199 m0 *1 7.755,136.5
X$17199 87 615 88 644 645 cell_1rw
* cell instance $17200 r0 *1 7.755,136.5
X$17200 87 614 88 644 645 cell_1rw
* cell instance $17201 m0 *1 7.755,139.23
X$17201 87 617 88 644 645 cell_1rw
* cell instance $17202 r0 *1 7.755,139.23
X$17202 87 616 88 644 645 cell_1rw
* cell instance $17203 m0 *1 7.755,141.96
X$17203 87 618 88 644 645 cell_1rw
* cell instance $17204 r0 *1 7.755,141.96
X$17204 87 619 88 644 645 cell_1rw
* cell instance $17205 m0 *1 7.755,144.69
X$17205 87 620 88 644 645 cell_1rw
* cell instance $17206 r0 *1 7.755,144.69
X$17206 87 621 88 644 645 cell_1rw
* cell instance $17207 m0 *1 7.755,147.42
X$17207 87 622 88 644 645 cell_1rw
* cell instance $17208 r0 *1 7.755,147.42
X$17208 87 623 88 644 645 cell_1rw
* cell instance $17209 m0 *1 7.755,150.15
X$17209 87 624 88 644 645 cell_1rw
* cell instance $17210 m0 *1 7.755,152.88
X$17210 87 626 88 644 645 cell_1rw
* cell instance $17211 r0 *1 7.755,150.15
X$17211 87 625 88 644 645 cell_1rw
* cell instance $17212 r0 *1 7.755,152.88
X$17212 87 627 88 644 645 cell_1rw
* cell instance $17213 m0 *1 7.755,155.61
X$17213 87 628 88 644 645 cell_1rw
* cell instance $17214 r0 *1 7.755,155.61
X$17214 87 629 88 644 645 cell_1rw
* cell instance $17215 m0 *1 7.755,158.34
X$17215 87 630 88 644 645 cell_1rw
* cell instance $17216 r0 *1 7.755,158.34
X$17216 87 631 88 644 645 cell_1rw
* cell instance $17217 m0 *1 7.755,161.07
X$17217 87 632 88 644 645 cell_1rw
* cell instance $17218 r0 *1 7.755,161.07
X$17218 87 633 88 644 645 cell_1rw
* cell instance $17219 m0 *1 7.755,163.8
X$17219 87 634 88 644 645 cell_1rw
* cell instance $17220 r0 *1 7.755,163.8
X$17220 87 635 88 644 645 cell_1rw
* cell instance $17221 m0 *1 7.755,166.53
X$17221 87 637 88 644 645 cell_1rw
* cell instance $17222 r0 *1 7.755,166.53
X$17222 87 636 88 644 645 cell_1rw
* cell instance $17223 m0 *1 7.755,169.26
X$17223 87 639 88 644 645 cell_1rw
* cell instance $17224 r0 *1 7.755,169.26
X$17224 87 638 88 644 645 cell_1rw
* cell instance $17225 m0 *1 7.755,171.99
X$17225 87 640 88 644 645 cell_1rw
* cell instance $17226 r0 *1 7.755,171.99
X$17226 87 641 88 644 645 cell_1rw
* cell instance $17227 m0 *1 7.755,174.72
X$17227 87 642 88 644 645 cell_1rw
* cell instance $17228 r0 *1 7.755,174.72
X$17228 87 643 88 644 645 cell_1rw
* cell instance $17229 r0 *1 8.46,87.36
X$17229 89 322 90 644 645 cell_1rw
* cell instance $17230 m0 *1 8.46,90.09
X$17230 89 581 90 644 645 cell_1rw
* cell instance $17231 r0 *1 8.46,90.09
X$17231 89 580 90 644 645 cell_1rw
* cell instance $17232 m0 *1 8.46,92.82
X$17232 89 583 90 644 645 cell_1rw
* cell instance $17233 r0 *1 8.46,92.82
X$17233 89 582 90 644 645 cell_1rw
* cell instance $17234 m0 *1 8.46,95.55
X$17234 89 584 90 644 645 cell_1rw
* cell instance $17235 r0 *1 8.46,95.55
X$17235 89 585 90 644 645 cell_1rw
* cell instance $17236 m0 *1 8.46,98.28
X$17236 89 586 90 644 645 cell_1rw
* cell instance $17237 r0 *1 8.46,98.28
X$17237 89 587 90 644 645 cell_1rw
* cell instance $17238 m0 *1 8.46,101.01
X$17238 89 588 90 644 645 cell_1rw
* cell instance $17239 r0 *1 8.46,101.01
X$17239 89 589 90 644 645 cell_1rw
* cell instance $17240 m0 *1 8.46,103.74
X$17240 89 590 90 644 645 cell_1rw
* cell instance $17241 m0 *1 8.46,106.47
X$17241 89 593 90 644 645 cell_1rw
* cell instance $17242 r0 *1 8.46,103.74
X$17242 89 591 90 644 645 cell_1rw
* cell instance $17243 r0 *1 8.46,106.47
X$17243 89 592 90 644 645 cell_1rw
* cell instance $17244 m0 *1 8.46,109.2
X$17244 89 594 90 644 645 cell_1rw
* cell instance $17245 r0 *1 8.46,109.2
X$17245 89 595 90 644 645 cell_1rw
* cell instance $17246 m0 *1 8.46,111.93
X$17246 89 597 90 644 645 cell_1rw
* cell instance $17247 m0 *1 8.46,114.66
X$17247 89 598 90 644 645 cell_1rw
* cell instance $17248 r0 *1 8.46,111.93
X$17248 89 596 90 644 645 cell_1rw
* cell instance $17249 r0 *1 8.46,114.66
X$17249 89 599 90 644 645 cell_1rw
* cell instance $17250 m0 *1 8.46,117.39
X$17250 89 600 90 644 645 cell_1rw
* cell instance $17251 r0 *1 8.46,117.39
X$17251 89 601 90 644 645 cell_1rw
* cell instance $17252 m0 *1 8.46,120.12
X$17252 89 602 90 644 645 cell_1rw
* cell instance $17253 r0 *1 8.46,120.12
X$17253 89 603 90 644 645 cell_1rw
* cell instance $17254 m0 *1 8.46,122.85
X$17254 89 604 90 644 645 cell_1rw
* cell instance $17255 m0 *1 8.46,125.58
X$17255 89 606 90 644 645 cell_1rw
* cell instance $17256 r0 *1 8.46,122.85
X$17256 89 605 90 644 645 cell_1rw
* cell instance $17257 r0 *1 8.46,125.58
X$17257 89 607 90 644 645 cell_1rw
* cell instance $17258 m0 *1 8.46,128.31
X$17258 89 609 90 644 645 cell_1rw
* cell instance $17259 r0 *1 8.46,128.31
X$17259 89 608 90 644 645 cell_1rw
* cell instance $17260 m0 *1 8.46,131.04
X$17260 89 610 90 644 645 cell_1rw
* cell instance $17261 r0 *1 8.46,131.04
X$17261 89 611 90 644 645 cell_1rw
* cell instance $17262 m0 *1 8.46,133.77
X$17262 89 612 90 644 645 cell_1rw
* cell instance $17263 m0 *1 8.46,136.5
X$17263 89 615 90 644 645 cell_1rw
* cell instance $17264 r0 *1 8.46,133.77
X$17264 89 613 90 644 645 cell_1rw
* cell instance $17265 r0 *1 8.46,136.5
X$17265 89 614 90 644 645 cell_1rw
* cell instance $17266 m0 *1 8.46,139.23
X$17266 89 617 90 644 645 cell_1rw
* cell instance $17267 r0 *1 8.46,139.23
X$17267 89 616 90 644 645 cell_1rw
* cell instance $17268 m0 *1 8.46,141.96
X$17268 89 618 90 644 645 cell_1rw
* cell instance $17269 r0 *1 8.46,141.96
X$17269 89 619 90 644 645 cell_1rw
* cell instance $17270 m0 *1 8.46,144.69
X$17270 89 620 90 644 645 cell_1rw
* cell instance $17271 r0 *1 8.46,144.69
X$17271 89 621 90 644 645 cell_1rw
* cell instance $17272 m0 *1 8.46,147.42
X$17272 89 622 90 644 645 cell_1rw
* cell instance $17273 r0 *1 8.46,147.42
X$17273 89 623 90 644 645 cell_1rw
* cell instance $17274 m0 *1 8.46,150.15
X$17274 89 624 90 644 645 cell_1rw
* cell instance $17275 r0 *1 8.46,150.15
X$17275 89 625 90 644 645 cell_1rw
* cell instance $17276 m0 *1 8.46,152.88
X$17276 89 626 90 644 645 cell_1rw
* cell instance $17277 r0 *1 8.46,152.88
X$17277 89 627 90 644 645 cell_1rw
* cell instance $17278 m0 *1 8.46,155.61
X$17278 89 628 90 644 645 cell_1rw
* cell instance $17279 r0 *1 8.46,155.61
X$17279 89 629 90 644 645 cell_1rw
* cell instance $17280 m0 *1 8.46,158.34
X$17280 89 630 90 644 645 cell_1rw
* cell instance $17281 r0 *1 8.46,158.34
X$17281 89 631 90 644 645 cell_1rw
* cell instance $17282 m0 *1 8.46,161.07
X$17282 89 632 90 644 645 cell_1rw
* cell instance $17283 r0 *1 8.46,161.07
X$17283 89 633 90 644 645 cell_1rw
* cell instance $17284 m0 *1 8.46,163.8
X$17284 89 634 90 644 645 cell_1rw
* cell instance $17285 r0 *1 8.46,163.8
X$17285 89 635 90 644 645 cell_1rw
* cell instance $17286 m0 *1 8.46,166.53
X$17286 89 637 90 644 645 cell_1rw
* cell instance $17287 r0 *1 8.46,166.53
X$17287 89 636 90 644 645 cell_1rw
* cell instance $17288 m0 *1 8.46,169.26
X$17288 89 639 90 644 645 cell_1rw
* cell instance $17289 r0 *1 8.46,169.26
X$17289 89 638 90 644 645 cell_1rw
* cell instance $17290 m0 *1 8.46,171.99
X$17290 89 640 90 644 645 cell_1rw
* cell instance $17291 r0 *1 8.46,171.99
X$17291 89 641 90 644 645 cell_1rw
* cell instance $17292 m0 *1 8.46,174.72
X$17292 89 642 90 644 645 cell_1rw
* cell instance $17293 r0 *1 8.46,174.72
X$17293 89 643 90 644 645 cell_1rw
* cell instance $17294 r0 *1 9.165,87.36
X$17294 91 322 92 644 645 cell_1rw
* cell instance $17295 m0 *1 9.165,90.09
X$17295 91 581 92 644 645 cell_1rw
* cell instance $17296 r0 *1 9.165,90.09
X$17296 91 580 92 644 645 cell_1rw
* cell instance $17297 m0 *1 9.165,92.82
X$17297 91 583 92 644 645 cell_1rw
* cell instance $17298 r0 *1 9.165,92.82
X$17298 91 582 92 644 645 cell_1rw
* cell instance $17299 m0 *1 9.165,95.55
X$17299 91 584 92 644 645 cell_1rw
* cell instance $17300 r0 *1 9.165,95.55
X$17300 91 585 92 644 645 cell_1rw
* cell instance $17301 m0 *1 9.165,98.28
X$17301 91 586 92 644 645 cell_1rw
* cell instance $17302 r0 *1 9.165,98.28
X$17302 91 587 92 644 645 cell_1rw
* cell instance $17303 m0 *1 9.165,101.01
X$17303 91 588 92 644 645 cell_1rw
* cell instance $17304 r0 *1 9.165,101.01
X$17304 91 589 92 644 645 cell_1rw
* cell instance $17305 m0 *1 9.165,103.74
X$17305 91 590 92 644 645 cell_1rw
* cell instance $17306 r0 *1 9.165,103.74
X$17306 91 591 92 644 645 cell_1rw
* cell instance $17307 m0 *1 9.165,106.47
X$17307 91 593 92 644 645 cell_1rw
* cell instance $17308 r0 *1 9.165,106.47
X$17308 91 592 92 644 645 cell_1rw
* cell instance $17309 m0 *1 9.165,109.2
X$17309 91 594 92 644 645 cell_1rw
* cell instance $17310 r0 *1 9.165,109.2
X$17310 91 595 92 644 645 cell_1rw
* cell instance $17311 m0 *1 9.165,111.93
X$17311 91 597 92 644 645 cell_1rw
* cell instance $17312 r0 *1 9.165,111.93
X$17312 91 596 92 644 645 cell_1rw
* cell instance $17313 m0 *1 9.165,114.66
X$17313 91 598 92 644 645 cell_1rw
* cell instance $17314 r0 *1 9.165,114.66
X$17314 91 599 92 644 645 cell_1rw
* cell instance $17315 m0 *1 9.165,117.39
X$17315 91 600 92 644 645 cell_1rw
* cell instance $17316 r0 *1 9.165,117.39
X$17316 91 601 92 644 645 cell_1rw
* cell instance $17317 m0 *1 9.165,120.12
X$17317 91 602 92 644 645 cell_1rw
* cell instance $17318 r0 *1 9.165,120.12
X$17318 91 603 92 644 645 cell_1rw
* cell instance $17319 m0 *1 9.165,122.85
X$17319 91 604 92 644 645 cell_1rw
* cell instance $17320 r0 *1 9.165,122.85
X$17320 91 605 92 644 645 cell_1rw
* cell instance $17321 m0 *1 9.165,125.58
X$17321 91 606 92 644 645 cell_1rw
* cell instance $17322 r0 *1 9.165,125.58
X$17322 91 607 92 644 645 cell_1rw
* cell instance $17323 m0 *1 9.165,128.31
X$17323 91 609 92 644 645 cell_1rw
* cell instance $17324 r0 *1 9.165,128.31
X$17324 91 608 92 644 645 cell_1rw
* cell instance $17325 m0 *1 9.165,131.04
X$17325 91 610 92 644 645 cell_1rw
* cell instance $17326 r0 *1 9.165,131.04
X$17326 91 611 92 644 645 cell_1rw
* cell instance $17327 m0 *1 9.165,133.77
X$17327 91 612 92 644 645 cell_1rw
* cell instance $17328 r0 *1 9.165,133.77
X$17328 91 613 92 644 645 cell_1rw
* cell instance $17329 m0 *1 9.165,136.5
X$17329 91 615 92 644 645 cell_1rw
* cell instance $17330 m0 *1 9.165,139.23
X$17330 91 617 92 644 645 cell_1rw
* cell instance $17331 r0 *1 9.165,136.5
X$17331 91 614 92 644 645 cell_1rw
* cell instance $17332 r0 *1 9.165,139.23
X$17332 91 616 92 644 645 cell_1rw
* cell instance $17333 m0 *1 9.165,141.96
X$17333 91 618 92 644 645 cell_1rw
* cell instance $17334 m0 *1 9.165,144.69
X$17334 91 620 92 644 645 cell_1rw
* cell instance $17335 r0 *1 9.165,141.96
X$17335 91 619 92 644 645 cell_1rw
* cell instance $17336 r0 *1 9.165,144.69
X$17336 91 621 92 644 645 cell_1rw
* cell instance $17337 m0 *1 9.165,147.42
X$17337 91 622 92 644 645 cell_1rw
* cell instance $17338 r0 *1 9.165,147.42
X$17338 91 623 92 644 645 cell_1rw
* cell instance $17339 m0 *1 9.165,150.15
X$17339 91 624 92 644 645 cell_1rw
* cell instance $17340 r0 *1 9.165,150.15
X$17340 91 625 92 644 645 cell_1rw
* cell instance $17341 m0 *1 9.165,152.88
X$17341 91 626 92 644 645 cell_1rw
* cell instance $17342 r0 *1 9.165,152.88
X$17342 91 627 92 644 645 cell_1rw
* cell instance $17343 m0 *1 9.165,155.61
X$17343 91 628 92 644 645 cell_1rw
* cell instance $17344 r0 *1 9.165,155.61
X$17344 91 629 92 644 645 cell_1rw
* cell instance $17345 m0 *1 9.165,158.34
X$17345 91 630 92 644 645 cell_1rw
* cell instance $17346 r0 *1 9.165,158.34
X$17346 91 631 92 644 645 cell_1rw
* cell instance $17347 m0 *1 9.165,161.07
X$17347 91 632 92 644 645 cell_1rw
* cell instance $17348 r0 *1 9.165,161.07
X$17348 91 633 92 644 645 cell_1rw
* cell instance $17349 m0 *1 9.165,163.8
X$17349 91 634 92 644 645 cell_1rw
* cell instance $17350 r0 *1 9.165,163.8
X$17350 91 635 92 644 645 cell_1rw
* cell instance $17351 m0 *1 9.165,166.53
X$17351 91 637 92 644 645 cell_1rw
* cell instance $17352 r0 *1 9.165,166.53
X$17352 91 636 92 644 645 cell_1rw
* cell instance $17353 m0 *1 9.165,169.26
X$17353 91 639 92 644 645 cell_1rw
* cell instance $17354 r0 *1 9.165,169.26
X$17354 91 638 92 644 645 cell_1rw
* cell instance $17355 m0 *1 9.165,171.99
X$17355 91 640 92 644 645 cell_1rw
* cell instance $17356 m0 *1 9.165,174.72
X$17356 91 642 92 644 645 cell_1rw
* cell instance $17357 r0 *1 9.165,171.99
X$17357 91 641 92 644 645 cell_1rw
* cell instance $17358 r0 *1 9.165,174.72
X$17358 91 643 92 644 645 cell_1rw
* cell instance $17359 m0 *1 9.87,90.09
X$17359 93 581 94 644 645 cell_1rw
* cell instance $17360 r0 *1 9.87,87.36
X$17360 93 322 94 644 645 cell_1rw
* cell instance $17361 r0 *1 9.87,90.09
X$17361 93 580 94 644 645 cell_1rw
* cell instance $17362 m0 *1 9.87,92.82
X$17362 93 583 94 644 645 cell_1rw
* cell instance $17363 r0 *1 9.87,92.82
X$17363 93 582 94 644 645 cell_1rw
* cell instance $17364 m0 *1 9.87,95.55
X$17364 93 584 94 644 645 cell_1rw
* cell instance $17365 m0 *1 9.87,98.28
X$17365 93 586 94 644 645 cell_1rw
* cell instance $17366 r0 *1 9.87,95.55
X$17366 93 585 94 644 645 cell_1rw
* cell instance $17367 r0 *1 9.87,98.28
X$17367 93 587 94 644 645 cell_1rw
* cell instance $17368 m0 *1 9.87,101.01
X$17368 93 588 94 644 645 cell_1rw
* cell instance $17369 r0 *1 9.87,101.01
X$17369 93 589 94 644 645 cell_1rw
* cell instance $17370 m0 *1 9.87,103.74
X$17370 93 590 94 644 645 cell_1rw
* cell instance $17371 r0 *1 9.87,103.74
X$17371 93 591 94 644 645 cell_1rw
* cell instance $17372 m0 *1 9.87,106.47
X$17372 93 593 94 644 645 cell_1rw
* cell instance $17373 r0 *1 9.87,106.47
X$17373 93 592 94 644 645 cell_1rw
* cell instance $17374 m0 *1 9.87,109.2
X$17374 93 594 94 644 645 cell_1rw
* cell instance $17375 r0 *1 9.87,109.2
X$17375 93 595 94 644 645 cell_1rw
* cell instance $17376 m0 *1 9.87,111.93
X$17376 93 597 94 644 645 cell_1rw
* cell instance $17377 r0 *1 9.87,111.93
X$17377 93 596 94 644 645 cell_1rw
* cell instance $17378 m0 *1 9.87,114.66
X$17378 93 598 94 644 645 cell_1rw
* cell instance $17379 r0 *1 9.87,114.66
X$17379 93 599 94 644 645 cell_1rw
* cell instance $17380 m0 *1 9.87,117.39
X$17380 93 600 94 644 645 cell_1rw
* cell instance $17381 m0 *1 9.87,120.12
X$17381 93 602 94 644 645 cell_1rw
* cell instance $17382 r0 *1 9.87,117.39
X$17382 93 601 94 644 645 cell_1rw
* cell instance $17383 m0 *1 9.87,122.85
X$17383 93 604 94 644 645 cell_1rw
* cell instance $17384 r0 *1 9.87,120.12
X$17384 93 603 94 644 645 cell_1rw
* cell instance $17385 r0 *1 9.87,122.85
X$17385 93 605 94 644 645 cell_1rw
* cell instance $17386 m0 *1 9.87,125.58
X$17386 93 606 94 644 645 cell_1rw
* cell instance $17387 r0 *1 9.87,125.58
X$17387 93 607 94 644 645 cell_1rw
* cell instance $17388 m0 *1 9.87,128.31
X$17388 93 609 94 644 645 cell_1rw
* cell instance $17389 m0 *1 9.87,131.04
X$17389 93 610 94 644 645 cell_1rw
* cell instance $17390 r0 *1 9.87,128.31
X$17390 93 608 94 644 645 cell_1rw
* cell instance $17391 r0 *1 9.87,131.04
X$17391 93 611 94 644 645 cell_1rw
* cell instance $17392 m0 *1 9.87,133.77
X$17392 93 612 94 644 645 cell_1rw
* cell instance $17393 r0 *1 9.87,133.77
X$17393 93 613 94 644 645 cell_1rw
* cell instance $17394 m0 *1 9.87,136.5
X$17394 93 615 94 644 645 cell_1rw
* cell instance $17395 r0 *1 9.87,136.5
X$17395 93 614 94 644 645 cell_1rw
* cell instance $17396 m0 *1 9.87,139.23
X$17396 93 617 94 644 645 cell_1rw
* cell instance $17397 r0 *1 9.87,139.23
X$17397 93 616 94 644 645 cell_1rw
* cell instance $17398 m0 *1 9.87,141.96
X$17398 93 618 94 644 645 cell_1rw
* cell instance $17399 r0 *1 9.87,141.96
X$17399 93 619 94 644 645 cell_1rw
* cell instance $17400 m0 *1 9.87,144.69
X$17400 93 620 94 644 645 cell_1rw
* cell instance $17401 r0 *1 9.87,144.69
X$17401 93 621 94 644 645 cell_1rw
* cell instance $17402 m0 *1 9.87,147.42
X$17402 93 622 94 644 645 cell_1rw
* cell instance $17403 m0 *1 9.87,150.15
X$17403 93 624 94 644 645 cell_1rw
* cell instance $17404 r0 *1 9.87,147.42
X$17404 93 623 94 644 645 cell_1rw
* cell instance $17405 r0 *1 9.87,150.15
X$17405 93 625 94 644 645 cell_1rw
* cell instance $17406 m0 *1 9.87,152.88
X$17406 93 626 94 644 645 cell_1rw
* cell instance $17407 r0 *1 9.87,152.88
X$17407 93 627 94 644 645 cell_1rw
* cell instance $17408 m0 *1 9.87,155.61
X$17408 93 628 94 644 645 cell_1rw
* cell instance $17409 r0 *1 9.87,155.61
X$17409 93 629 94 644 645 cell_1rw
* cell instance $17410 m0 *1 9.87,158.34
X$17410 93 630 94 644 645 cell_1rw
* cell instance $17411 r0 *1 9.87,158.34
X$17411 93 631 94 644 645 cell_1rw
* cell instance $17412 m0 *1 9.87,161.07
X$17412 93 632 94 644 645 cell_1rw
* cell instance $17413 r0 *1 9.87,161.07
X$17413 93 633 94 644 645 cell_1rw
* cell instance $17414 m0 *1 9.87,163.8
X$17414 93 634 94 644 645 cell_1rw
* cell instance $17415 m0 *1 9.87,166.53
X$17415 93 637 94 644 645 cell_1rw
* cell instance $17416 r0 *1 9.87,163.8
X$17416 93 635 94 644 645 cell_1rw
* cell instance $17417 r0 *1 9.87,166.53
X$17417 93 636 94 644 645 cell_1rw
* cell instance $17418 m0 *1 9.87,169.26
X$17418 93 639 94 644 645 cell_1rw
* cell instance $17419 r0 *1 9.87,169.26
X$17419 93 638 94 644 645 cell_1rw
* cell instance $17420 m0 *1 9.87,171.99
X$17420 93 640 94 644 645 cell_1rw
* cell instance $17421 r0 *1 9.87,171.99
X$17421 93 641 94 644 645 cell_1rw
* cell instance $17422 m0 *1 9.87,174.72
X$17422 93 642 94 644 645 cell_1rw
* cell instance $17423 r0 *1 9.87,174.72
X$17423 93 643 94 644 645 cell_1rw
* cell instance $17424 r0 *1 10.575,87.36
X$17424 95 322 96 644 645 cell_1rw
* cell instance $17425 m0 *1 10.575,90.09
X$17425 95 581 96 644 645 cell_1rw
* cell instance $17426 r0 *1 10.575,90.09
X$17426 95 580 96 644 645 cell_1rw
* cell instance $17427 m0 *1 10.575,92.82
X$17427 95 583 96 644 645 cell_1rw
* cell instance $17428 r0 *1 10.575,92.82
X$17428 95 582 96 644 645 cell_1rw
* cell instance $17429 m0 *1 10.575,95.55
X$17429 95 584 96 644 645 cell_1rw
* cell instance $17430 r0 *1 10.575,95.55
X$17430 95 585 96 644 645 cell_1rw
* cell instance $17431 m0 *1 10.575,98.28
X$17431 95 586 96 644 645 cell_1rw
* cell instance $17432 r0 *1 10.575,98.28
X$17432 95 587 96 644 645 cell_1rw
* cell instance $17433 m0 *1 10.575,101.01
X$17433 95 588 96 644 645 cell_1rw
* cell instance $17434 r0 *1 10.575,101.01
X$17434 95 589 96 644 645 cell_1rw
* cell instance $17435 m0 *1 10.575,103.74
X$17435 95 590 96 644 645 cell_1rw
* cell instance $17436 r0 *1 10.575,103.74
X$17436 95 591 96 644 645 cell_1rw
* cell instance $17437 m0 *1 10.575,106.47
X$17437 95 593 96 644 645 cell_1rw
* cell instance $17438 r0 *1 10.575,106.47
X$17438 95 592 96 644 645 cell_1rw
* cell instance $17439 m0 *1 10.575,109.2
X$17439 95 594 96 644 645 cell_1rw
* cell instance $17440 m0 *1 10.575,111.93
X$17440 95 597 96 644 645 cell_1rw
* cell instance $17441 r0 *1 10.575,109.2
X$17441 95 595 96 644 645 cell_1rw
* cell instance $17442 r0 *1 10.575,111.93
X$17442 95 596 96 644 645 cell_1rw
* cell instance $17443 m0 *1 10.575,114.66
X$17443 95 598 96 644 645 cell_1rw
* cell instance $17444 r0 *1 10.575,114.66
X$17444 95 599 96 644 645 cell_1rw
* cell instance $17445 m0 *1 10.575,117.39
X$17445 95 600 96 644 645 cell_1rw
* cell instance $17446 r0 *1 10.575,117.39
X$17446 95 601 96 644 645 cell_1rw
* cell instance $17447 m0 *1 10.575,120.12
X$17447 95 602 96 644 645 cell_1rw
* cell instance $17448 r0 *1 10.575,120.12
X$17448 95 603 96 644 645 cell_1rw
* cell instance $17449 m0 *1 10.575,122.85
X$17449 95 604 96 644 645 cell_1rw
* cell instance $17450 m0 *1 10.575,125.58
X$17450 95 606 96 644 645 cell_1rw
* cell instance $17451 r0 *1 10.575,122.85
X$17451 95 605 96 644 645 cell_1rw
* cell instance $17452 r0 *1 10.575,125.58
X$17452 95 607 96 644 645 cell_1rw
* cell instance $17453 m0 *1 10.575,128.31
X$17453 95 609 96 644 645 cell_1rw
* cell instance $17454 r0 *1 10.575,128.31
X$17454 95 608 96 644 645 cell_1rw
* cell instance $17455 m0 *1 10.575,131.04
X$17455 95 610 96 644 645 cell_1rw
* cell instance $17456 r0 *1 10.575,131.04
X$17456 95 611 96 644 645 cell_1rw
* cell instance $17457 m0 *1 10.575,133.77
X$17457 95 612 96 644 645 cell_1rw
* cell instance $17458 r0 *1 10.575,133.77
X$17458 95 613 96 644 645 cell_1rw
* cell instance $17459 m0 *1 10.575,136.5
X$17459 95 615 96 644 645 cell_1rw
* cell instance $17460 m0 *1 10.575,139.23
X$17460 95 617 96 644 645 cell_1rw
* cell instance $17461 r0 *1 10.575,136.5
X$17461 95 614 96 644 645 cell_1rw
* cell instance $17462 r0 *1 10.575,139.23
X$17462 95 616 96 644 645 cell_1rw
* cell instance $17463 m0 *1 10.575,141.96
X$17463 95 618 96 644 645 cell_1rw
* cell instance $17464 r0 *1 10.575,141.96
X$17464 95 619 96 644 645 cell_1rw
* cell instance $17465 m0 *1 10.575,144.69
X$17465 95 620 96 644 645 cell_1rw
* cell instance $17466 r0 *1 10.575,144.69
X$17466 95 621 96 644 645 cell_1rw
* cell instance $17467 m0 *1 10.575,147.42
X$17467 95 622 96 644 645 cell_1rw
* cell instance $17468 r0 *1 10.575,147.42
X$17468 95 623 96 644 645 cell_1rw
* cell instance $17469 m0 *1 10.575,150.15
X$17469 95 624 96 644 645 cell_1rw
* cell instance $17470 r0 *1 10.575,150.15
X$17470 95 625 96 644 645 cell_1rw
* cell instance $17471 m0 *1 10.575,152.88
X$17471 95 626 96 644 645 cell_1rw
* cell instance $17472 r0 *1 10.575,152.88
X$17472 95 627 96 644 645 cell_1rw
* cell instance $17473 m0 *1 10.575,155.61
X$17473 95 628 96 644 645 cell_1rw
* cell instance $17474 r0 *1 10.575,155.61
X$17474 95 629 96 644 645 cell_1rw
* cell instance $17475 m0 *1 10.575,158.34
X$17475 95 630 96 644 645 cell_1rw
* cell instance $17476 r0 *1 10.575,158.34
X$17476 95 631 96 644 645 cell_1rw
* cell instance $17477 m0 *1 10.575,161.07
X$17477 95 632 96 644 645 cell_1rw
* cell instance $17478 r0 *1 10.575,161.07
X$17478 95 633 96 644 645 cell_1rw
* cell instance $17479 m0 *1 10.575,163.8
X$17479 95 634 96 644 645 cell_1rw
* cell instance $17480 r0 *1 10.575,163.8
X$17480 95 635 96 644 645 cell_1rw
* cell instance $17481 m0 *1 10.575,166.53
X$17481 95 637 96 644 645 cell_1rw
* cell instance $17482 m0 *1 10.575,169.26
X$17482 95 639 96 644 645 cell_1rw
* cell instance $17483 r0 *1 10.575,166.53
X$17483 95 636 96 644 645 cell_1rw
* cell instance $17484 m0 *1 10.575,171.99
X$17484 95 640 96 644 645 cell_1rw
* cell instance $17485 r0 *1 10.575,169.26
X$17485 95 638 96 644 645 cell_1rw
* cell instance $17486 m0 *1 10.575,174.72
X$17486 95 642 96 644 645 cell_1rw
* cell instance $17487 r0 *1 10.575,171.99
X$17487 95 641 96 644 645 cell_1rw
* cell instance $17488 r0 *1 10.575,174.72
X$17488 95 643 96 644 645 cell_1rw
* cell instance $17489 r0 *1 11.28,87.36
X$17489 97 322 98 644 645 cell_1rw
* cell instance $17490 m0 *1 11.28,90.09
X$17490 97 581 98 644 645 cell_1rw
* cell instance $17491 r0 *1 11.28,90.09
X$17491 97 580 98 644 645 cell_1rw
* cell instance $17492 m0 *1 11.28,92.82
X$17492 97 583 98 644 645 cell_1rw
* cell instance $17493 m0 *1 11.28,95.55
X$17493 97 584 98 644 645 cell_1rw
* cell instance $17494 r0 *1 11.28,92.82
X$17494 97 582 98 644 645 cell_1rw
* cell instance $17495 m0 *1 11.28,98.28
X$17495 97 586 98 644 645 cell_1rw
* cell instance $17496 r0 *1 11.28,95.55
X$17496 97 585 98 644 645 cell_1rw
* cell instance $17497 r0 *1 11.28,98.28
X$17497 97 587 98 644 645 cell_1rw
* cell instance $17498 m0 *1 11.28,101.01
X$17498 97 588 98 644 645 cell_1rw
* cell instance $17499 m0 *1 11.28,103.74
X$17499 97 590 98 644 645 cell_1rw
* cell instance $17500 r0 *1 11.28,101.01
X$17500 97 589 98 644 645 cell_1rw
* cell instance $17501 m0 *1 11.28,106.47
X$17501 97 593 98 644 645 cell_1rw
* cell instance $17502 r0 *1 11.28,103.74
X$17502 97 591 98 644 645 cell_1rw
* cell instance $17503 r0 *1 11.28,106.47
X$17503 97 592 98 644 645 cell_1rw
* cell instance $17504 m0 *1 11.28,109.2
X$17504 97 594 98 644 645 cell_1rw
* cell instance $17505 r0 *1 11.28,109.2
X$17505 97 595 98 644 645 cell_1rw
* cell instance $17506 m0 *1 11.28,111.93
X$17506 97 597 98 644 645 cell_1rw
* cell instance $17507 r0 *1 11.28,111.93
X$17507 97 596 98 644 645 cell_1rw
* cell instance $17508 m0 *1 11.28,114.66
X$17508 97 598 98 644 645 cell_1rw
* cell instance $17509 r0 *1 11.28,114.66
X$17509 97 599 98 644 645 cell_1rw
* cell instance $17510 m0 *1 11.28,117.39
X$17510 97 600 98 644 645 cell_1rw
* cell instance $17511 m0 *1 11.28,120.12
X$17511 97 602 98 644 645 cell_1rw
* cell instance $17512 r0 *1 11.28,117.39
X$17512 97 601 98 644 645 cell_1rw
* cell instance $17513 r0 *1 11.28,120.12
X$17513 97 603 98 644 645 cell_1rw
* cell instance $17514 m0 *1 11.28,122.85
X$17514 97 604 98 644 645 cell_1rw
* cell instance $17515 r0 *1 11.28,122.85
X$17515 97 605 98 644 645 cell_1rw
* cell instance $17516 m0 *1 11.28,125.58
X$17516 97 606 98 644 645 cell_1rw
* cell instance $17517 r0 *1 11.28,125.58
X$17517 97 607 98 644 645 cell_1rw
* cell instance $17518 m0 *1 11.28,128.31
X$17518 97 609 98 644 645 cell_1rw
* cell instance $17519 m0 *1 11.28,131.04
X$17519 97 610 98 644 645 cell_1rw
* cell instance $17520 r0 *1 11.28,128.31
X$17520 97 608 98 644 645 cell_1rw
* cell instance $17521 m0 *1 11.28,133.77
X$17521 97 612 98 644 645 cell_1rw
* cell instance $17522 r0 *1 11.28,131.04
X$17522 97 611 98 644 645 cell_1rw
* cell instance $17523 r0 *1 11.28,133.77
X$17523 97 613 98 644 645 cell_1rw
* cell instance $17524 m0 *1 11.28,136.5
X$17524 97 615 98 644 645 cell_1rw
* cell instance $17525 r0 *1 11.28,136.5
X$17525 97 614 98 644 645 cell_1rw
* cell instance $17526 m0 *1 11.28,139.23
X$17526 97 617 98 644 645 cell_1rw
* cell instance $17527 r0 *1 11.28,139.23
X$17527 97 616 98 644 645 cell_1rw
* cell instance $17528 m0 *1 11.28,141.96
X$17528 97 618 98 644 645 cell_1rw
* cell instance $17529 r0 *1 11.28,141.96
X$17529 97 619 98 644 645 cell_1rw
* cell instance $17530 m0 *1 11.28,144.69
X$17530 97 620 98 644 645 cell_1rw
* cell instance $17531 r0 *1 11.28,144.69
X$17531 97 621 98 644 645 cell_1rw
* cell instance $17532 m0 *1 11.28,147.42
X$17532 97 622 98 644 645 cell_1rw
* cell instance $17533 r0 *1 11.28,147.42
X$17533 97 623 98 644 645 cell_1rw
* cell instance $17534 m0 *1 11.28,150.15
X$17534 97 624 98 644 645 cell_1rw
* cell instance $17535 r0 *1 11.28,150.15
X$17535 97 625 98 644 645 cell_1rw
* cell instance $17536 m0 *1 11.28,152.88
X$17536 97 626 98 644 645 cell_1rw
* cell instance $17537 r0 *1 11.28,152.88
X$17537 97 627 98 644 645 cell_1rw
* cell instance $17538 m0 *1 11.28,155.61
X$17538 97 628 98 644 645 cell_1rw
* cell instance $17539 r0 *1 11.28,155.61
X$17539 97 629 98 644 645 cell_1rw
* cell instance $17540 m0 *1 11.28,158.34
X$17540 97 630 98 644 645 cell_1rw
* cell instance $17541 m0 *1 11.28,161.07
X$17541 97 632 98 644 645 cell_1rw
* cell instance $17542 r0 *1 11.28,158.34
X$17542 97 631 98 644 645 cell_1rw
* cell instance $17543 r0 *1 11.28,161.07
X$17543 97 633 98 644 645 cell_1rw
* cell instance $17544 m0 *1 11.28,163.8
X$17544 97 634 98 644 645 cell_1rw
* cell instance $17545 r0 *1 11.28,163.8
X$17545 97 635 98 644 645 cell_1rw
* cell instance $17546 m0 *1 11.28,166.53
X$17546 97 637 98 644 645 cell_1rw
* cell instance $17547 m0 *1 11.28,169.26
X$17547 97 639 98 644 645 cell_1rw
* cell instance $17548 r0 *1 11.28,166.53
X$17548 97 636 98 644 645 cell_1rw
* cell instance $17549 r0 *1 11.28,169.26
X$17549 97 638 98 644 645 cell_1rw
* cell instance $17550 m0 *1 11.28,171.99
X$17550 97 640 98 644 645 cell_1rw
* cell instance $17551 m0 *1 11.28,174.72
X$17551 97 642 98 644 645 cell_1rw
* cell instance $17552 r0 *1 11.28,171.99
X$17552 97 641 98 644 645 cell_1rw
* cell instance $17553 r0 *1 11.28,174.72
X$17553 97 643 98 644 645 cell_1rw
* cell instance $17554 r0 *1 11.985,87.36
X$17554 99 322 100 644 645 cell_1rw
* cell instance $17555 m0 *1 11.985,90.09
X$17555 99 581 100 644 645 cell_1rw
* cell instance $17556 r0 *1 11.985,90.09
X$17556 99 580 100 644 645 cell_1rw
* cell instance $17557 m0 *1 11.985,92.82
X$17557 99 583 100 644 645 cell_1rw
* cell instance $17558 r0 *1 11.985,92.82
X$17558 99 582 100 644 645 cell_1rw
* cell instance $17559 m0 *1 11.985,95.55
X$17559 99 584 100 644 645 cell_1rw
* cell instance $17560 m0 *1 11.985,98.28
X$17560 99 586 100 644 645 cell_1rw
* cell instance $17561 r0 *1 11.985,95.55
X$17561 99 585 100 644 645 cell_1rw
* cell instance $17562 r0 *1 11.985,98.28
X$17562 99 587 100 644 645 cell_1rw
* cell instance $17563 m0 *1 11.985,101.01
X$17563 99 588 100 644 645 cell_1rw
* cell instance $17564 r0 *1 11.985,101.01
X$17564 99 589 100 644 645 cell_1rw
* cell instance $17565 m0 *1 11.985,103.74
X$17565 99 590 100 644 645 cell_1rw
* cell instance $17566 r0 *1 11.985,103.74
X$17566 99 591 100 644 645 cell_1rw
* cell instance $17567 m0 *1 11.985,106.47
X$17567 99 593 100 644 645 cell_1rw
* cell instance $17568 r0 *1 11.985,106.47
X$17568 99 592 100 644 645 cell_1rw
* cell instance $17569 m0 *1 11.985,109.2
X$17569 99 594 100 644 645 cell_1rw
* cell instance $17570 r0 *1 11.985,109.2
X$17570 99 595 100 644 645 cell_1rw
* cell instance $17571 m0 *1 11.985,111.93
X$17571 99 597 100 644 645 cell_1rw
* cell instance $17572 m0 *1 11.985,114.66
X$17572 99 598 100 644 645 cell_1rw
* cell instance $17573 r0 *1 11.985,111.93
X$17573 99 596 100 644 645 cell_1rw
* cell instance $17574 r0 *1 11.985,114.66
X$17574 99 599 100 644 645 cell_1rw
* cell instance $17575 m0 *1 11.985,117.39
X$17575 99 600 100 644 645 cell_1rw
* cell instance $17576 r0 *1 11.985,117.39
X$17576 99 601 100 644 645 cell_1rw
* cell instance $17577 m0 *1 11.985,120.12
X$17577 99 602 100 644 645 cell_1rw
* cell instance $17578 r0 *1 11.985,120.12
X$17578 99 603 100 644 645 cell_1rw
* cell instance $17579 m0 *1 11.985,122.85
X$17579 99 604 100 644 645 cell_1rw
* cell instance $17580 r0 *1 11.985,122.85
X$17580 99 605 100 644 645 cell_1rw
* cell instance $17581 m0 *1 11.985,125.58
X$17581 99 606 100 644 645 cell_1rw
* cell instance $17582 r0 *1 11.985,125.58
X$17582 99 607 100 644 645 cell_1rw
* cell instance $17583 m0 *1 11.985,128.31
X$17583 99 609 100 644 645 cell_1rw
* cell instance $17584 m0 *1 11.985,131.04
X$17584 99 610 100 644 645 cell_1rw
* cell instance $17585 r0 *1 11.985,128.31
X$17585 99 608 100 644 645 cell_1rw
* cell instance $17586 r0 *1 11.985,131.04
X$17586 99 611 100 644 645 cell_1rw
* cell instance $17587 m0 *1 11.985,133.77
X$17587 99 612 100 644 645 cell_1rw
* cell instance $17588 r0 *1 11.985,133.77
X$17588 99 613 100 644 645 cell_1rw
* cell instance $17589 m0 *1 11.985,136.5
X$17589 99 615 100 644 645 cell_1rw
* cell instance $17590 r0 *1 11.985,136.5
X$17590 99 614 100 644 645 cell_1rw
* cell instance $17591 m0 *1 11.985,139.23
X$17591 99 617 100 644 645 cell_1rw
* cell instance $17592 r0 *1 11.985,139.23
X$17592 99 616 100 644 645 cell_1rw
* cell instance $17593 m0 *1 11.985,141.96
X$17593 99 618 100 644 645 cell_1rw
* cell instance $17594 r0 *1 11.985,141.96
X$17594 99 619 100 644 645 cell_1rw
* cell instance $17595 m0 *1 11.985,144.69
X$17595 99 620 100 644 645 cell_1rw
* cell instance $17596 m0 *1 11.985,147.42
X$17596 99 622 100 644 645 cell_1rw
* cell instance $17597 r0 *1 11.985,144.69
X$17597 99 621 100 644 645 cell_1rw
* cell instance $17598 r0 *1 11.985,147.42
X$17598 99 623 100 644 645 cell_1rw
* cell instance $17599 m0 *1 11.985,150.15
X$17599 99 624 100 644 645 cell_1rw
* cell instance $17600 r0 *1 11.985,150.15
X$17600 99 625 100 644 645 cell_1rw
* cell instance $17601 m0 *1 11.985,152.88
X$17601 99 626 100 644 645 cell_1rw
* cell instance $17602 r0 *1 11.985,152.88
X$17602 99 627 100 644 645 cell_1rw
* cell instance $17603 m0 *1 11.985,155.61
X$17603 99 628 100 644 645 cell_1rw
* cell instance $17604 r0 *1 11.985,155.61
X$17604 99 629 100 644 645 cell_1rw
* cell instance $17605 m0 *1 11.985,158.34
X$17605 99 630 100 644 645 cell_1rw
* cell instance $17606 r0 *1 11.985,158.34
X$17606 99 631 100 644 645 cell_1rw
* cell instance $17607 m0 *1 11.985,161.07
X$17607 99 632 100 644 645 cell_1rw
* cell instance $17608 m0 *1 11.985,163.8
X$17608 99 634 100 644 645 cell_1rw
* cell instance $17609 r0 *1 11.985,161.07
X$17609 99 633 100 644 645 cell_1rw
* cell instance $17610 r0 *1 11.985,163.8
X$17610 99 635 100 644 645 cell_1rw
* cell instance $17611 m0 *1 11.985,166.53
X$17611 99 637 100 644 645 cell_1rw
* cell instance $17612 r0 *1 11.985,166.53
X$17612 99 636 100 644 645 cell_1rw
* cell instance $17613 m0 *1 11.985,169.26
X$17613 99 639 100 644 645 cell_1rw
* cell instance $17614 m0 *1 11.985,171.99
X$17614 99 640 100 644 645 cell_1rw
* cell instance $17615 r0 *1 11.985,169.26
X$17615 99 638 100 644 645 cell_1rw
* cell instance $17616 r0 *1 11.985,171.99
X$17616 99 641 100 644 645 cell_1rw
* cell instance $17617 m0 *1 11.985,174.72
X$17617 99 642 100 644 645 cell_1rw
* cell instance $17618 r0 *1 11.985,174.72
X$17618 99 643 100 644 645 cell_1rw
* cell instance $17619 m0 *1 12.69,90.09
X$17619 101 581 102 644 645 cell_1rw
* cell instance $17620 r0 *1 12.69,87.36
X$17620 101 322 102 644 645 cell_1rw
* cell instance $17621 r0 *1 12.69,90.09
X$17621 101 580 102 644 645 cell_1rw
* cell instance $17622 m0 *1 12.69,92.82
X$17622 101 583 102 644 645 cell_1rw
* cell instance $17623 r0 *1 12.69,92.82
X$17623 101 582 102 644 645 cell_1rw
* cell instance $17624 m0 *1 12.69,95.55
X$17624 101 584 102 644 645 cell_1rw
* cell instance $17625 r0 *1 12.69,95.55
X$17625 101 585 102 644 645 cell_1rw
* cell instance $17626 m0 *1 12.69,98.28
X$17626 101 586 102 644 645 cell_1rw
* cell instance $17627 r0 *1 12.69,98.28
X$17627 101 587 102 644 645 cell_1rw
* cell instance $17628 m0 *1 12.69,101.01
X$17628 101 588 102 644 645 cell_1rw
* cell instance $17629 r0 *1 12.69,101.01
X$17629 101 589 102 644 645 cell_1rw
* cell instance $17630 m0 *1 12.69,103.74
X$17630 101 590 102 644 645 cell_1rw
* cell instance $17631 r0 *1 12.69,103.74
X$17631 101 591 102 644 645 cell_1rw
* cell instance $17632 m0 *1 12.69,106.47
X$17632 101 593 102 644 645 cell_1rw
* cell instance $17633 r0 *1 12.69,106.47
X$17633 101 592 102 644 645 cell_1rw
* cell instance $17634 m0 *1 12.69,109.2
X$17634 101 594 102 644 645 cell_1rw
* cell instance $17635 r0 *1 12.69,109.2
X$17635 101 595 102 644 645 cell_1rw
* cell instance $17636 m0 *1 12.69,111.93
X$17636 101 597 102 644 645 cell_1rw
* cell instance $17637 m0 *1 12.69,114.66
X$17637 101 598 102 644 645 cell_1rw
* cell instance $17638 r0 *1 12.69,111.93
X$17638 101 596 102 644 645 cell_1rw
* cell instance $17639 r0 *1 12.69,114.66
X$17639 101 599 102 644 645 cell_1rw
* cell instance $17640 m0 *1 12.69,117.39
X$17640 101 600 102 644 645 cell_1rw
* cell instance $17641 r0 *1 12.69,117.39
X$17641 101 601 102 644 645 cell_1rw
* cell instance $17642 m0 *1 12.69,120.12
X$17642 101 602 102 644 645 cell_1rw
* cell instance $17643 r0 *1 12.69,120.12
X$17643 101 603 102 644 645 cell_1rw
* cell instance $17644 m0 *1 12.69,122.85
X$17644 101 604 102 644 645 cell_1rw
* cell instance $17645 r0 *1 12.69,122.85
X$17645 101 605 102 644 645 cell_1rw
* cell instance $17646 m0 *1 12.69,125.58
X$17646 101 606 102 644 645 cell_1rw
* cell instance $17647 m0 *1 12.69,128.31
X$17647 101 609 102 644 645 cell_1rw
* cell instance $17648 r0 *1 12.69,125.58
X$17648 101 607 102 644 645 cell_1rw
* cell instance $17649 r0 *1 12.69,128.31
X$17649 101 608 102 644 645 cell_1rw
* cell instance $17650 m0 *1 12.69,131.04
X$17650 101 610 102 644 645 cell_1rw
* cell instance $17651 r0 *1 12.69,131.04
X$17651 101 611 102 644 645 cell_1rw
* cell instance $17652 m0 *1 12.69,133.77
X$17652 101 612 102 644 645 cell_1rw
* cell instance $17653 r0 *1 12.69,133.77
X$17653 101 613 102 644 645 cell_1rw
* cell instance $17654 m0 *1 12.69,136.5
X$17654 101 615 102 644 645 cell_1rw
* cell instance $17655 r0 *1 12.69,136.5
X$17655 101 614 102 644 645 cell_1rw
* cell instance $17656 m0 *1 12.69,139.23
X$17656 101 617 102 644 645 cell_1rw
* cell instance $17657 r0 *1 12.69,139.23
X$17657 101 616 102 644 645 cell_1rw
* cell instance $17658 m0 *1 12.69,141.96
X$17658 101 618 102 644 645 cell_1rw
* cell instance $17659 r0 *1 12.69,141.96
X$17659 101 619 102 644 645 cell_1rw
* cell instance $17660 m0 *1 12.69,144.69
X$17660 101 620 102 644 645 cell_1rw
* cell instance $17661 m0 *1 12.69,147.42
X$17661 101 622 102 644 645 cell_1rw
* cell instance $17662 r0 *1 12.69,144.69
X$17662 101 621 102 644 645 cell_1rw
* cell instance $17663 r0 *1 12.69,147.42
X$17663 101 623 102 644 645 cell_1rw
* cell instance $17664 m0 *1 12.69,150.15
X$17664 101 624 102 644 645 cell_1rw
* cell instance $17665 r0 *1 12.69,150.15
X$17665 101 625 102 644 645 cell_1rw
* cell instance $17666 m0 *1 12.69,152.88
X$17666 101 626 102 644 645 cell_1rw
* cell instance $17667 r0 *1 12.69,152.88
X$17667 101 627 102 644 645 cell_1rw
* cell instance $17668 m0 *1 12.69,155.61
X$17668 101 628 102 644 645 cell_1rw
* cell instance $17669 m0 *1 12.69,158.34
X$17669 101 630 102 644 645 cell_1rw
* cell instance $17670 r0 *1 12.69,155.61
X$17670 101 629 102 644 645 cell_1rw
* cell instance $17671 r0 *1 12.69,158.34
X$17671 101 631 102 644 645 cell_1rw
* cell instance $17672 m0 *1 12.69,161.07
X$17672 101 632 102 644 645 cell_1rw
* cell instance $17673 r0 *1 12.69,161.07
X$17673 101 633 102 644 645 cell_1rw
* cell instance $17674 m0 *1 12.69,163.8
X$17674 101 634 102 644 645 cell_1rw
* cell instance $17675 r0 *1 12.69,163.8
X$17675 101 635 102 644 645 cell_1rw
* cell instance $17676 m0 *1 12.69,166.53
X$17676 101 637 102 644 645 cell_1rw
* cell instance $17677 r0 *1 12.69,166.53
X$17677 101 636 102 644 645 cell_1rw
* cell instance $17678 m0 *1 12.69,169.26
X$17678 101 639 102 644 645 cell_1rw
* cell instance $17679 m0 *1 12.69,171.99
X$17679 101 640 102 644 645 cell_1rw
* cell instance $17680 r0 *1 12.69,169.26
X$17680 101 638 102 644 645 cell_1rw
* cell instance $17681 r0 *1 12.69,171.99
X$17681 101 641 102 644 645 cell_1rw
* cell instance $17682 m0 *1 12.69,174.72
X$17682 101 642 102 644 645 cell_1rw
* cell instance $17683 r0 *1 12.69,174.72
X$17683 101 643 102 644 645 cell_1rw
* cell instance $17684 m0 *1 13.395,90.09
X$17684 103 581 104 644 645 cell_1rw
* cell instance $17685 r0 *1 13.395,87.36
X$17685 103 322 104 644 645 cell_1rw
* cell instance $17686 r0 *1 13.395,90.09
X$17686 103 580 104 644 645 cell_1rw
* cell instance $17687 m0 *1 13.395,92.82
X$17687 103 583 104 644 645 cell_1rw
* cell instance $17688 r0 *1 13.395,92.82
X$17688 103 582 104 644 645 cell_1rw
* cell instance $17689 m0 *1 13.395,95.55
X$17689 103 584 104 644 645 cell_1rw
* cell instance $17690 r0 *1 13.395,95.55
X$17690 103 585 104 644 645 cell_1rw
* cell instance $17691 m0 *1 13.395,98.28
X$17691 103 586 104 644 645 cell_1rw
* cell instance $17692 r0 *1 13.395,98.28
X$17692 103 587 104 644 645 cell_1rw
* cell instance $17693 m0 *1 13.395,101.01
X$17693 103 588 104 644 645 cell_1rw
* cell instance $17694 r0 *1 13.395,101.01
X$17694 103 589 104 644 645 cell_1rw
* cell instance $17695 m0 *1 13.395,103.74
X$17695 103 590 104 644 645 cell_1rw
* cell instance $17696 r0 *1 13.395,103.74
X$17696 103 591 104 644 645 cell_1rw
* cell instance $17697 m0 *1 13.395,106.47
X$17697 103 593 104 644 645 cell_1rw
* cell instance $17698 r0 *1 13.395,106.47
X$17698 103 592 104 644 645 cell_1rw
* cell instance $17699 m0 *1 13.395,109.2
X$17699 103 594 104 644 645 cell_1rw
* cell instance $17700 r0 *1 13.395,109.2
X$17700 103 595 104 644 645 cell_1rw
* cell instance $17701 m0 *1 13.395,111.93
X$17701 103 597 104 644 645 cell_1rw
* cell instance $17702 r0 *1 13.395,111.93
X$17702 103 596 104 644 645 cell_1rw
* cell instance $17703 m0 *1 13.395,114.66
X$17703 103 598 104 644 645 cell_1rw
* cell instance $17704 r0 *1 13.395,114.66
X$17704 103 599 104 644 645 cell_1rw
* cell instance $17705 m0 *1 13.395,117.39
X$17705 103 600 104 644 645 cell_1rw
* cell instance $17706 r0 *1 13.395,117.39
X$17706 103 601 104 644 645 cell_1rw
* cell instance $17707 m0 *1 13.395,120.12
X$17707 103 602 104 644 645 cell_1rw
* cell instance $17708 r0 *1 13.395,120.12
X$17708 103 603 104 644 645 cell_1rw
* cell instance $17709 m0 *1 13.395,122.85
X$17709 103 604 104 644 645 cell_1rw
* cell instance $17710 r0 *1 13.395,122.85
X$17710 103 605 104 644 645 cell_1rw
* cell instance $17711 m0 *1 13.395,125.58
X$17711 103 606 104 644 645 cell_1rw
* cell instance $17712 r0 *1 13.395,125.58
X$17712 103 607 104 644 645 cell_1rw
* cell instance $17713 m0 *1 13.395,128.31
X$17713 103 609 104 644 645 cell_1rw
* cell instance $17714 r0 *1 13.395,128.31
X$17714 103 608 104 644 645 cell_1rw
* cell instance $17715 m0 *1 13.395,131.04
X$17715 103 610 104 644 645 cell_1rw
* cell instance $17716 r0 *1 13.395,131.04
X$17716 103 611 104 644 645 cell_1rw
* cell instance $17717 m0 *1 13.395,133.77
X$17717 103 612 104 644 645 cell_1rw
* cell instance $17718 m0 *1 13.395,136.5
X$17718 103 615 104 644 645 cell_1rw
* cell instance $17719 r0 *1 13.395,133.77
X$17719 103 613 104 644 645 cell_1rw
* cell instance $17720 m0 *1 13.395,139.23
X$17720 103 617 104 644 645 cell_1rw
* cell instance $17721 r0 *1 13.395,136.5
X$17721 103 614 104 644 645 cell_1rw
* cell instance $17722 r0 *1 13.395,139.23
X$17722 103 616 104 644 645 cell_1rw
* cell instance $17723 m0 *1 13.395,141.96
X$17723 103 618 104 644 645 cell_1rw
* cell instance $17724 r0 *1 13.395,141.96
X$17724 103 619 104 644 645 cell_1rw
* cell instance $17725 m0 *1 13.395,144.69
X$17725 103 620 104 644 645 cell_1rw
* cell instance $17726 r0 *1 13.395,144.69
X$17726 103 621 104 644 645 cell_1rw
* cell instance $17727 m0 *1 13.395,147.42
X$17727 103 622 104 644 645 cell_1rw
* cell instance $17728 r0 *1 13.395,147.42
X$17728 103 623 104 644 645 cell_1rw
* cell instance $17729 m0 *1 13.395,150.15
X$17729 103 624 104 644 645 cell_1rw
* cell instance $17730 r0 *1 13.395,150.15
X$17730 103 625 104 644 645 cell_1rw
* cell instance $17731 m0 *1 13.395,152.88
X$17731 103 626 104 644 645 cell_1rw
* cell instance $17732 r0 *1 13.395,152.88
X$17732 103 627 104 644 645 cell_1rw
* cell instance $17733 m0 *1 13.395,155.61
X$17733 103 628 104 644 645 cell_1rw
* cell instance $17734 r0 *1 13.395,155.61
X$17734 103 629 104 644 645 cell_1rw
* cell instance $17735 m0 *1 13.395,158.34
X$17735 103 630 104 644 645 cell_1rw
* cell instance $17736 r0 *1 13.395,158.34
X$17736 103 631 104 644 645 cell_1rw
* cell instance $17737 m0 *1 13.395,161.07
X$17737 103 632 104 644 645 cell_1rw
* cell instance $17738 r0 *1 13.395,161.07
X$17738 103 633 104 644 645 cell_1rw
* cell instance $17739 m0 *1 13.395,163.8
X$17739 103 634 104 644 645 cell_1rw
* cell instance $17740 r0 *1 13.395,163.8
X$17740 103 635 104 644 645 cell_1rw
* cell instance $17741 m0 *1 13.395,166.53
X$17741 103 637 104 644 645 cell_1rw
* cell instance $17742 r0 *1 13.395,166.53
X$17742 103 636 104 644 645 cell_1rw
* cell instance $17743 m0 *1 13.395,169.26
X$17743 103 639 104 644 645 cell_1rw
* cell instance $17744 r0 *1 13.395,169.26
X$17744 103 638 104 644 645 cell_1rw
* cell instance $17745 m0 *1 13.395,171.99
X$17745 103 640 104 644 645 cell_1rw
* cell instance $17746 m0 *1 13.395,174.72
X$17746 103 642 104 644 645 cell_1rw
* cell instance $17747 r0 *1 13.395,171.99
X$17747 103 641 104 644 645 cell_1rw
* cell instance $17748 r0 *1 13.395,174.72
X$17748 103 643 104 644 645 cell_1rw
* cell instance $17749 m0 *1 14.1,90.09
X$17749 105 581 106 644 645 cell_1rw
* cell instance $17750 r0 *1 14.1,87.36
X$17750 105 322 106 644 645 cell_1rw
* cell instance $17751 r0 *1 14.1,90.09
X$17751 105 580 106 644 645 cell_1rw
* cell instance $17752 m0 *1 14.1,92.82
X$17752 105 583 106 644 645 cell_1rw
* cell instance $17753 m0 *1 14.1,95.55
X$17753 105 584 106 644 645 cell_1rw
* cell instance $17754 r0 *1 14.1,92.82
X$17754 105 582 106 644 645 cell_1rw
* cell instance $17755 r0 *1 14.1,95.55
X$17755 105 585 106 644 645 cell_1rw
* cell instance $17756 m0 *1 14.1,98.28
X$17756 105 586 106 644 645 cell_1rw
* cell instance $17757 r0 *1 14.1,98.28
X$17757 105 587 106 644 645 cell_1rw
* cell instance $17758 m0 *1 14.1,101.01
X$17758 105 588 106 644 645 cell_1rw
* cell instance $17759 r0 *1 14.1,101.01
X$17759 105 589 106 644 645 cell_1rw
* cell instance $17760 m0 *1 14.1,103.74
X$17760 105 590 106 644 645 cell_1rw
* cell instance $17761 r0 *1 14.1,103.74
X$17761 105 591 106 644 645 cell_1rw
* cell instance $17762 m0 *1 14.1,106.47
X$17762 105 593 106 644 645 cell_1rw
* cell instance $17763 r0 *1 14.1,106.47
X$17763 105 592 106 644 645 cell_1rw
* cell instance $17764 m0 *1 14.1,109.2
X$17764 105 594 106 644 645 cell_1rw
* cell instance $17765 r0 *1 14.1,109.2
X$17765 105 595 106 644 645 cell_1rw
* cell instance $17766 m0 *1 14.1,111.93
X$17766 105 597 106 644 645 cell_1rw
* cell instance $17767 r0 *1 14.1,111.93
X$17767 105 596 106 644 645 cell_1rw
* cell instance $17768 m0 *1 14.1,114.66
X$17768 105 598 106 644 645 cell_1rw
* cell instance $17769 m0 *1 14.1,117.39
X$17769 105 600 106 644 645 cell_1rw
* cell instance $17770 r0 *1 14.1,114.66
X$17770 105 599 106 644 645 cell_1rw
* cell instance $17771 r0 *1 14.1,117.39
X$17771 105 601 106 644 645 cell_1rw
* cell instance $17772 m0 *1 14.1,120.12
X$17772 105 602 106 644 645 cell_1rw
* cell instance $17773 r0 *1 14.1,120.12
X$17773 105 603 106 644 645 cell_1rw
* cell instance $17774 m0 *1 14.1,122.85
X$17774 105 604 106 644 645 cell_1rw
* cell instance $17775 r0 *1 14.1,122.85
X$17775 105 605 106 644 645 cell_1rw
* cell instance $17776 m0 *1 14.1,125.58
X$17776 105 606 106 644 645 cell_1rw
* cell instance $17777 r0 *1 14.1,125.58
X$17777 105 607 106 644 645 cell_1rw
* cell instance $17778 m0 *1 14.1,128.31
X$17778 105 609 106 644 645 cell_1rw
* cell instance $17779 r0 *1 14.1,128.31
X$17779 105 608 106 644 645 cell_1rw
* cell instance $17780 m0 *1 14.1,131.04
X$17780 105 610 106 644 645 cell_1rw
* cell instance $17781 r0 *1 14.1,131.04
X$17781 105 611 106 644 645 cell_1rw
* cell instance $17782 m0 *1 14.1,133.77
X$17782 105 612 106 644 645 cell_1rw
* cell instance $17783 r0 *1 14.1,133.77
X$17783 105 613 106 644 645 cell_1rw
* cell instance $17784 m0 *1 14.1,136.5
X$17784 105 615 106 644 645 cell_1rw
* cell instance $17785 r0 *1 14.1,136.5
X$17785 105 614 106 644 645 cell_1rw
* cell instance $17786 m0 *1 14.1,139.23
X$17786 105 617 106 644 645 cell_1rw
* cell instance $17787 r0 *1 14.1,139.23
X$17787 105 616 106 644 645 cell_1rw
* cell instance $17788 m0 *1 14.1,141.96
X$17788 105 618 106 644 645 cell_1rw
* cell instance $17789 r0 *1 14.1,141.96
X$17789 105 619 106 644 645 cell_1rw
* cell instance $17790 m0 *1 14.1,144.69
X$17790 105 620 106 644 645 cell_1rw
* cell instance $17791 r0 *1 14.1,144.69
X$17791 105 621 106 644 645 cell_1rw
* cell instance $17792 m0 *1 14.1,147.42
X$17792 105 622 106 644 645 cell_1rw
* cell instance $17793 r0 *1 14.1,147.42
X$17793 105 623 106 644 645 cell_1rw
* cell instance $17794 m0 *1 14.1,150.15
X$17794 105 624 106 644 645 cell_1rw
* cell instance $17795 r0 *1 14.1,150.15
X$17795 105 625 106 644 645 cell_1rw
* cell instance $17796 m0 *1 14.1,152.88
X$17796 105 626 106 644 645 cell_1rw
* cell instance $17797 r0 *1 14.1,152.88
X$17797 105 627 106 644 645 cell_1rw
* cell instance $17798 m0 *1 14.1,155.61
X$17798 105 628 106 644 645 cell_1rw
* cell instance $17799 r0 *1 14.1,155.61
X$17799 105 629 106 644 645 cell_1rw
* cell instance $17800 m0 *1 14.1,158.34
X$17800 105 630 106 644 645 cell_1rw
* cell instance $17801 r0 *1 14.1,158.34
X$17801 105 631 106 644 645 cell_1rw
* cell instance $17802 m0 *1 14.1,161.07
X$17802 105 632 106 644 645 cell_1rw
* cell instance $17803 r0 *1 14.1,161.07
X$17803 105 633 106 644 645 cell_1rw
* cell instance $17804 m0 *1 14.1,163.8
X$17804 105 634 106 644 645 cell_1rw
* cell instance $17805 r0 *1 14.1,163.8
X$17805 105 635 106 644 645 cell_1rw
* cell instance $17806 m0 *1 14.1,166.53
X$17806 105 637 106 644 645 cell_1rw
* cell instance $17807 r0 *1 14.1,166.53
X$17807 105 636 106 644 645 cell_1rw
* cell instance $17808 m0 *1 14.1,169.26
X$17808 105 639 106 644 645 cell_1rw
* cell instance $17809 m0 *1 14.1,171.99
X$17809 105 640 106 644 645 cell_1rw
* cell instance $17810 r0 *1 14.1,169.26
X$17810 105 638 106 644 645 cell_1rw
* cell instance $17811 r0 *1 14.1,171.99
X$17811 105 641 106 644 645 cell_1rw
* cell instance $17812 m0 *1 14.1,174.72
X$17812 105 642 106 644 645 cell_1rw
* cell instance $17813 r0 *1 14.1,174.72
X$17813 105 643 106 644 645 cell_1rw
* cell instance $17814 m0 *1 14.805,90.09
X$17814 107 581 108 644 645 cell_1rw
* cell instance $17815 r0 *1 14.805,87.36
X$17815 107 322 108 644 645 cell_1rw
* cell instance $17816 r0 *1 14.805,90.09
X$17816 107 580 108 644 645 cell_1rw
* cell instance $17817 m0 *1 14.805,92.82
X$17817 107 583 108 644 645 cell_1rw
* cell instance $17818 r0 *1 14.805,92.82
X$17818 107 582 108 644 645 cell_1rw
* cell instance $17819 m0 *1 14.805,95.55
X$17819 107 584 108 644 645 cell_1rw
* cell instance $17820 r0 *1 14.805,95.55
X$17820 107 585 108 644 645 cell_1rw
* cell instance $17821 m0 *1 14.805,98.28
X$17821 107 586 108 644 645 cell_1rw
* cell instance $17822 r0 *1 14.805,98.28
X$17822 107 587 108 644 645 cell_1rw
* cell instance $17823 m0 *1 14.805,101.01
X$17823 107 588 108 644 645 cell_1rw
* cell instance $17824 m0 *1 14.805,103.74
X$17824 107 590 108 644 645 cell_1rw
* cell instance $17825 r0 *1 14.805,101.01
X$17825 107 589 108 644 645 cell_1rw
* cell instance $17826 r0 *1 14.805,103.74
X$17826 107 591 108 644 645 cell_1rw
* cell instance $17827 m0 *1 14.805,106.47
X$17827 107 593 108 644 645 cell_1rw
* cell instance $17828 r0 *1 14.805,106.47
X$17828 107 592 108 644 645 cell_1rw
* cell instance $17829 m0 *1 14.805,109.2
X$17829 107 594 108 644 645 cell_1rw
* cell instance $17830 r0 *1 14.805,109.2
X$17830 107 595 108 644 645 cell_1rw
* cell instance $17831 m0 *1 14.805,111.93
X$17831 107 597 108 644 645 cell_1rw
* cell instance $17832 r0 *1 14.805,111.93
X$17832 107 596 108 644 645 cell_1rw
* cell instance $17833 m0 *1 14.805,114.66
X$17833 107 598 108 644 645 cell_1rw
* cell instance $17834 r0 *1 14.805,114.66
X$17834 107 599 108 644 645 cell_1rw
* cell instance $17835 m0 *1 14.805,117.39
X$17835 107 600 108 644 645 cell_1rw
* cell instance $17836 r0 *1 14.805,117.39
X$17836 107 601 108 644 645 cell_1rw
* cell instance $17837 m0 *1 14.805,120.12
X$17837 107 602 108 644 645 cell_1rw
* cell instance $17838 r0 *1 14.805,120.12
X$17838 107 603 108 644 645 cell_1rw
* cell instance $17839 m0 *1 14.805,122.85
X$17839 107 604 108 644 645 cell_1rw
* cell instance $17840 r0 *1 14.805,122.85
X$17840 107 605 108 644 645 cell_1rw
* cell instance $17841 m0 *1 14.805,125.58
X$17841 107 606 108 644 645 cell_1rw
* cell instance $17842 m0 *1 14.805,128.31
X$17842 107 609 108 644 645 cell_1rw
* cell instance $17843 r0 *1 14.805,125.58
X$17843 107 607 108 644 645 cell_1rw
* cell instance $17844 r0 *1 14.805,128.31
X$17844 107 608 108 644 645 cell_1rw
* cell instance $17845 m0 *1 14.805,131.04
X$17845 107 610 108 644 645 cell_1rw
* cell instance $17846 r0 *1 14.805,131.04
X$17846 107 611 108 644 645 cell_1rw
* cell instance $17847 m0 *1 14.805,133.77
X$17847 107 612 108 644 645 cell_1rw
* cell instance $17848 r0 *1 14.805,133.77
X$17848 107 613 108 644 645 cell_1rw
* cell instance $17849 m0 *1 14.805,136.5
X$17849 107 615 108 644 645 cell_1rw
* cell instance $17850 r0 *1 14.805,136.5
X$17850 107 614 108 644 645 cell_1rw
* cell instance $17851 m0 *1 14.805,139.23
X$17851 107 617 108 644 645 cell_1rw
* cell instance $17852 r0 *1 14.805,139.23
X$17852 107 616 108 644 645 cell_1rw
* cell instance $17853 m0 *1 14.805,141.96
X$17853 107 618 108 644 645 cell_1rw
* cell instance $17854 r0 *1 14.805,141.96
X$17854 107 619 108 644 645 cell_1rw
* cell instance $17855 m0 *1 14.805,144.69
X$17855 107 620 108 644 645 cell_1rw
* cell instance $17856 r0 *1 14.805,144.69
X$17856 107 621 108 644 645 cell_1rw
* cell instance $17857 m0 *1 14.805,147.42
X$17857 107 622 108 644 645 cell_1rw
* cell instance $17858 r0 *1 14.805,147.42
X$17858 107 623 108 644 645 cell_1rw
* cell instance $17859 m0 *1 14.805,150.15
X$17859 107 624 108 644 645 cell_1rw
* cell instance $17860 r0 *1 14.805,150.15
X$17860 107 625 108 644 645 cell_1rw
* cell instance $17861 m0 *1 14.805,152.88
X$17861 107 626 108 644 645 cell_1rw
* cell instance $17862 r0 *1 14.805,152.88
X$17862 107 627 108 644 645 cell_1rw
* cell instance $17863 m0 *1 14.805,155.61
X$17863 107 628 108 644 645 cell_1rw
* cell instance $17864 r0 *1 14.805,155.61
X$17864 107 629 108 644 645 cell_1rw
* cell instance $17865 m0 *1 14.805,158.34
X$17865 107 630 108 644 645 cell_1rw
* cell instance $17866 r0 *1 14.805,158.34
X$17866 107 631 108 644 645 cell_1rw
* cell instance $17867 m0 *1 14.805,161.07
X$17867 107 632 108 644 645 cell_1rw
* cell instance $17868 r0 *1 14.805,161.07
X$17868 107 633 108 644 645 cell_1rw
* cell instance $17869 m0 *1 14.805,163.8
X$17869 107 634 108 644 645 cell_1rw
* cell instance $17870 r0 *1 14.805,163.8
X$17870 107 635 108 644 645 cell_1rw
* cell instance $17871 m0 *1 14.805,166.53
X$17871 107 637 108 644 645 cell_1rw
* cell instance $17872 r0 *1 14.805,166.53
X$17872 107 636 108 644 645 cell_1rw
* cell instance $17873 m0 *1 14.805,169.26
X$17873 107 639 108 644 645 cell_1rw
* cell instance $17874 r0 *1 14.805,169.26
X$17874 107 638 108 644 645 cell_1rw
* cell instance $17875 m0 *1 14.805,171.99
X$17875 107 640 108 644 645 cell_1rw
* cell instance $17876 r0 *1 14.805,171.99
X$17876 107 641 108 644 645 cell_1rw
* cell instance $17877 m0 *1 14.805,174.72
X$17877 107 642 108 644 645 cell_1rw
* cell instance $17878 r0 *1 14.805,174.72
X$17878 107 643 108 644 645 cell_1rw
* cell instance $17879 r0 *1 15.51,87.36
X$17879 109 322 110 644 645 cell_1rw
* cell instance $17880 m0 *1 15.51,90.09
X$17880 109 581 110 644 645 cell_1rw
* cell instance $17881 r0 *1 15.51,90.09
X$17881 109 580 110 644 645 cell_1rw
* cell instance $17882 m0 *1 15.51,92.82
X$17882 109 583 110 644 645 cell_1rw
* cell instance $17883 r0 *1 15.51,92.82
X$17883 109 582 110 644 645 cell_1rw
* cell instance $17884 m0 *1 15.51,95.55
X$17884 109 584 110 644 645 cell_1rw
* cell instance $17885 r0 *1 15.51,95.55
X$17885 109 585 110 644 645 cell_1rw
* cell instance $17886 m0 *1 15.51,98.28
X$17886 109 586 110 644 645 cell_1rw
* cell instance $17887 r0 *1 15.51,98.28
X$17887 109 587 110 644 645 cell_1rw
* cell instance $17888 m0 *1 15.51,101.01
X$17888 109 588 110 644 645 cell_1rw
* cell instance $17889 r0 *1 15.51,101.01
X$17889 109 589 110 644 645 cell_1rw
* cell instance $17890 m0 *1 15.51,103.74
X$17890 109 590 110 644 645 cell_1rw
* cell instance $17891 r0 *1 15.51,103.74
X$17891 109 591 110 644 645 cell_1rw
* cell instance $17892 m0 *1 15.51,106.47
X$17892 109 593 110 644 645 cell_1rw
* cell instance $17893 m0 *1 15.51,109.2
X$17893 109 594 110 644 645 cell_1rw
* cell instance $17894 r0 *1 15.51,106.47
X$17894 109 592 110 644 645 cell_1rw
* cell instance $17895 r0 *1 15.51,109.2
X$17895 109 595 110 644 645 cell_1rw
* cell instance $17896 m0 *1 15.51,111.93
X$17896 109 597 110 644 645 cell_1rw
* cell instance $17897 r0 *1 15.51,111.93
X$17897 109 596 110 644 645 cell_1rw
* cell instance $17898 m0 *1 15.51,114.66
X$17898 109 598 110 644 645 cell_1rw
* cell instance $17899 r0 *1 15.51,114.66
X$17899 109 599 110 644 645 cell_1rw
* cell instance $17900 m0 *1 15.51,117.39
X$17900 109 600 110 644 645 cell_1rw
* cell instance $17901 r0 *1 15.51,117.39
X$17901 109 601 110 644 645 cell_1rw
* cell instance $17902 m0 *1 15.51,120.12
X$17902 109 602 110 644 645 cell_1rw
* cell instance $17903 r0 *1 15.51,120.12
X$17903 109 603 110 644 645 cell_1rw
* cell instance $17904 m0 *1 15.51,122.85
X$17904 109 604 110 644 645 cell_1rw
* cell instance $17905 r0 *1 15.51,122.85
X$17905 109 605 110 644 645 cell_1rw
* cell instance $17906 m0 *1 15.51,125.58
X$17906 109 606 110 644 645 cell_1rw
* cell instance $17907 r0 *1 15.51,125.58
X$17907 109 607 110 644 645 cell_1rw
* cell instance $17908 m0 *1 15.51,128.31
X$17908 109 609 110 644 645 cell_1rw
* cell instance $17909 r0 *1 15.51,128.31
X$17909 109 608 110 644 645 cell_1rw
* cell instance $17910 m0 *1 15.51,131.04
X$17910 109 610 110 644 645 cell_1rw
* cell instance $17911 r0 *1 15.51,131.04
X$17911 109 611 110 644 645 cell_1rw
* cell instance $17912 m0 *1 15.51,133.77
X$17912 109 612 110 644 645 cell_1rw
* cell instance $17913 r0 *1 15.51,133.77
X$17913 109 613 110 644 645 cell_1rw
* cell instance $17914 m0 *1 15.51,136.5
X$17914 109 615 110 644 645 cell_1rw
* cell instance $17915 r0 *1 15.51,136.5
X$17915 109 614 110 644 645 cell_1rw
* cell instance $17916 m0 *1 15.51,139.23
X$17916 109 617 110 644 645 cell_1rw
* cell instance $17917 m0 *1 15.51,141.96
X$17917 109 618 110 644 645 cell_1rw
* cell instance $17918 r0 *1 15.51,139.23
X$17918 109 616 110 644 645 cell_1rw
* cell instance $17919 r0 *1 15.51,141.96
X$17919 109 619 110 644 645 cell_1rw
* cell instance $17920 m0 *1 15.51,144.69
X$17920 109 620 110 644 645 cell_1rw
* cell instance $17921 r0 *1 15.51,144.69
X$17921 109 621 110 644 645 cell_1rw
* cell instance $17922 m0 *1 15.51,147.42
X$17922 109 622 110 644 645 cell_1rw
* cell instance $17923 r0 *1 15.51,147.42
X$17923 109 623 110 644 645 cell_1rw
* cell instance $17924 m0 *1 15.51,150.15
X$17924 109 624 110 644 645 cell_1rw
* cell instance $17925 r0 *1 15.51,150.15
X$17925 109 625 110 644 645 cell_1rw
* cell instance $17926 m0 *1 15.51,152.88
X$17926 109 626 110 644 645 cell_1rw
* cell instance $17927 r0 *1 15.51,152.88
X$17927 109 627 110 644 645 cell_1rw
* cell instance $17928 m0 *1 15.51,155.61
X$17928 109 628 110 644 645 cell_1rw
* cell instance $17929 r0 *1 15.51,155.61
X$17929 109 629 110 644 645 cell_1rw
* cell instance $17930 m0 *1 15.51,158.34
X$17930 109 630 110 644 645 cell_1rw
* cell instance $17931 r0 *1 15.51,158.34
X$17931 109 631 110 644 645 cell_1rw
* cell instance $17932 m0 *1 15.51,161.07
X$17932 109 632 110 644 645 cell_1rw
* cell instance $17933 m0 *1 15.51,163.8
X$17933 109 634 110 644 645 cell_1rw
* cell instance $17934 r0 *1 15.51,161.07
X$17934 109 633 110 644 645 cell_1rw
* cell instance $17935 m0 *1 15.51,166.53
X$17935 109 637 110 644 645 cell_1rw
* cell instance $17936 r0 *1 15.51,163.8
X$17936 109 635 110 644 645 cell_1rw
* cell instance $17937 r0 *1 15.51,166.53
X$17937 109 636 110 644 645 cell_1rw
* cell instance $17938 m0 *1 15.51,169.26
X$17938 109 639 110 644 645 cell_1rw
* cell instance $17939 m0 *1 15.51,171.99
X$17939 109 640 110 644 645 cell_1rw
* cell instance $17940 r0 *1 15.51,169.26
X$17940 109 638 110 644 645 cell_1rw
* cell instance $17941 r0 *1 15.51,171.99
X$17941 109 641 110 644 645 cell_1rw
* cell instance $17942 m0 *1 15.51,174.72
X$17942 109 642 110 644 645 cell_1rw
* cell instance $17943 r0 *1 15.51,174.72
X$17943 109 643 110 644 645 cell_1rw
* cell instance $17944 r0 *1 16.215,87.36
X$17944 111 322 112 644 645 cell_1rw
* cell instance $17945 m0 *1 16.215,90.09
X$17945 111 581 112 644 645 cell_1rw
* cell instance $17946 r0 *1 16.215,90.09
X$17946 111 580 112 644 645 cell_1rw
* cell instance $17947 m0 *1 16.215,92.82
X$17947 111 583 112 644 645 cell_1rw
* cell instance $17948 r0 *1 16.215,92.82
X$17948 111 582 112 644 645 cell_1rw
* cell instance $17949 m0 *1 16.215,95.55
X$17949 111 584 112 644 645 cell_1rw
* cell instance $17950 r0 *1 16.215,95.55
X$17950 111 585 112 644 645 cell_1rw
* cell instance $17951 m0 *1 16.215,98.28
X$17951 111 586 112 644 645 cell_1rw
* cell instance $17952 r0 *1 16.215,98.28
X$17952 111 587 112 644 645 cell_1rw
* cell instance $17953 m0 *1 16.215,101.01
X$17953 111 588 112 644 645 cell_1rw
* cell instance $17954 r0 *1 16.215,101.01
X$17954 111 589 112 644 645 cell_1rw
* cell instance $17955 m0 *1 16.215,103.74
X$17955 111 590 112 644 645 cell_1rw
* cell instance $17956 m0 *1 16.215,106.47
X$17956 111 593 112 644 645 cell_1rw
* cell instance $17957 r0 *1 16.215,103.74
X$17957 111 591 112 644 645 cell_1rw
* cell instance $17958 r0 *1 16.215,106.47
X$17958 111 592 112 644 645 cell_1rw
* cell instance $17959 m0 *1 16.215,109.2
X$17959 111 594 112 644 645 cell_1rw
* cell instance $17960 r0 *1 16.215,109.2
X$17960 111 595 112 644 645 cell_1rw
* cell instance $17961 m0 *1 16.215,111.93
X$17961 111 597 112 644 645 cell_1rw
* cell instance $17962 r0 *1 16.215,111.93
X$17962 111 596 112 644 645 cell_1rw
* cell instance $17963 m0 *1 16.215,114.66
X$17963 111 598 112 644 645 cell_1rw
* cell instance $17964 r0 *1 16.215,114.66
X$17964 111 599 112 644 645 cell_1rw
* cell instance $17965 m0 *1 16.215,117.39
X$17965 111 600 112 644 645 cell_1rw
* cell instance $17966 m0 *1 16.215,120.12
X$17966 111 602 112 644 645 cell_1rw
* cell instance $17967 r0 *1 16.215,117.39
X$17967 111 601 112 644 645 cell_1rw
* cell instance $17968 r0 *1 16.215,120.12
X$17968 111 603 112 644 645 cell_1rw
* cell instance $17969 m0 *1 16.215,122.85
X$17969 111 604 112 644 645 cell_1rw
* cell instance $17970 r0 *1 16.215,122.85
X$17970 111 605 112 644 645 cell_1rw
* cell instance $17971 m0 *1 16.215,125.58
X$17971 111 606 112 644 645 cell_1rw
* cell instance $17972 r0 *1 16.215,125.58
X$17972 111 607 112 644 645 cell_1rw
* cell instance $17973 m0 *1 16.215,128.31
X$17973 111 609 112 644 645 cell_1rw
* cell instance $17974 r0 *1 16.215,128.31
X$17974 111 608 112 644 645 cell_1rw
* cell instance $17975 m0 *1 16.215,131.04
X$17975 111 610 112 644 645 cell_1rw
* cell instance $17976 m0 *1 16.215,133.77
X$17976 111 612 112 644 645 cell_1rw
* cell instance $17977 r0 *1 16.215,131.04
X$17977 111 611 112 644 645 cell_1rw
* cell instance $17978 r0 *1 16.215,133.77
X$17978 111 613 112 644 645 cell_1rw
* cell instance $17979 m0 *1 16.215,136.5
X$17979 111 615 112 644 645 cell_1rw
* cell instance $17980 r0 *1 16.215,136.5
X$17980 111 614 112 644 645 cell_1rw
* cell instance $17981 m0 *1 16.215,139.23
X$17981 111 617 112 644 645 cell_1rw
* cell instance $17982 r0 *1 16.215,139.23
X$17982 111 616 112 644 645 cell_1rw
* cell instance $17983 m0 *1 16.215,141.96
X$17983 111 618 112 644 645 cell_1rw
* cell instance $17984 m0 *1 16.215,144.69
X$17984 111 620 112 644 645 cell_1rw
* cell instance $17985 r0 *1 16.215,141.96
X$17985 111 619 112 644 645 cell_1rw
* cell instance $17986 r0 *1 16.215,144.69
X$17986 111 621 112 644 645 cell_1rw
* cell instance $17987 m0 *1 16.215,147.42
X$17987 111 622 112 644 645 cell_1rw
* cell instance $17988 r0 *1 16.215,147.42
X$17988 111 623 112 644 645 cell_1rw
* cell instance $17989 m0 *1 16.215,150.15
X$17989 111 624 112 644 645 cell_1rw
* cell instance $17990 r0 *1 16.215,150.15
X$17990 111 625 112 644 645 cell_1rw
* cell instance $17991 m0 *1 16.215,152.88
X$17991 111 626 112 644 645 cell_1rw
* cell instance $17992 r0 *1 16.215,152.88
X$17992 111 627 112 644 645 cell_1rw
* cell instance $17993 m0 *1 16.215,155.61
X$17993 111 628 112 644 645 cell_1rw
* cell instance $17994 m0 *1 16.215,158.34
X$17994 111 630 112 644 645 cell_1rw
* cell instance $17995 r0 *1 16.215,155.61
X$17995 111 629 112 644 645 cell_1rw
* cell instance $17996 m0 *1 16.215,161.07
X$17996 111 632 112 644 645 cell_1rw
* cell instance $17997 r0 *1 16.215,158.34
X$17997 111 631 112 644 645 cell_1rw
* cell instance $17998 r0 *1 16.215,161.07
X$17998 111 633 112 644 645 cell_1rw
* cell instance $17999 m0 *1 16.215,163.8
X$17999 111 634 112 644 645 cell_1rw
* cell instance $18000 m0 *1 16.215,166.53
X$18000 111 637 112 644 645 cell_1rw
* cell instance $18001 r0 *1 16.215,163.8
X$18001 111 635 112 644 645 cell_1rw
* cell instance $18002 r0 *1 16.215,166.53
X$18002 111 636 112 644 645 cell_1rw
* cell instance $18003 m0 *1 16.215,169.26
X$18003 111 639 112 644 645 cell_1rw
* cell instance $18004 r0 *1 16.215,169.26
X$18004 111 638 112 644 645 cell_1rw
* cell instance $18005 m0 *1 16.215,171.99
X$18005 111 640 112 644 645 cell_1rw
* cell instance $18006 r0 *1 16.215,171.99
X$18006 111 641 112 644 645 cell_1rw
* cell instance $18007 m0 *1 16.215,174.72
X$18007 111 642 112 644 645 cell_1rw
* cell instance $18008 r0 *1 16.215,174.72
X$18008 111 643 112 644 645 cell_1rw
* cell instance $18009 r0 *1 16.92,87.36
X$18009 113 322 114 644 645 cell_1rw
* cell instance $18010 m0 *1 16.92,90.09
X$18010 113 581 114 644 645 cell_1rw
* cell instance $18011 r0 *1 16.92,90.09
X$18011 113 580 114 644 645 cell_1rw
* cell instance $18012 m0 *1 16.92,92.82
X$18012 113 583 114 644 645 cell_1rw
* cell instance $18013 m0 *1 16.92,95.55
X$18013 113 584 114 644 645 cell_1rw
* cell instance $18014 r0 *1 16.92,92.82
X$18014 113 582 114 644 645 cell_1rw
* cell instance $18015 r0 *1 16.92,95.55
X$18015 113 585 114 644 645 cell_1rw
* cell instance $18016 m0 *1 16.92,98.28
X$18016 113 586 114 644 645 cell_1rw
* cell instance $18017 r0 *1 16.92,98.28
X$18017 113 587 114 644 645 cell_1rw
* cell instance $18018 m0 *1 16.92,101.01
X$18018 113 588 114 644 645 cell_1rw
* cell instance $18019 r0 *1 16.92,101.01
X$18019 113 589 114 644 645 cell_1rw
* cell instance $18020 m0 *1 16.92,103.74
X$18020 113 590 114 644 645 cell_1rw
* cell instance $18021 r0 *1 16.92,103.74
X$18021 113 591 114 644 645 cell_1rw
* cell instance $18022 m0 *1 16.92,106.47
X$18022 113 593 114 644 645 cell_1rw
* cell instance $18023 r0 *1 16.92,106.47
X$18023 113 592 114 644 645 cell_1rw
* cell instance $18024 m0 *1 16.92,109.2
X$18024 113 594 114 644 645 cell_1rw
* cell instance $18025 r0 *1 16.92,109.2
X$18025 113 595 114 644 645 cell_1rw
* cell instance $18026 m0 *1 16.92,111.93
X$18026 113 597 114 644 645 cell_1rw
* cell instance $18027 m0 *1 16.92,114.66
X$18027 113 598 114 644 645 cell_1rw
* cell instance $18028 r0 *1 16.92,111.93
X$18028 113 596 114 644 645 cell_1rw
* cell instance $18029 r0 *1 16.92,114.66
X$18029 113 599 114 644 645 cell_1rw
* cell instance $18030 m0 *1 16.92,117.39
X$18030 113 600 114 644 645 cell_1rw
* cell instance $18031 r0 *1 16.92,117.39
X$18031 113 601 114 644 645 cell_1rw
* cell instance $18032 m0 *1 16.92,120.12
X$18032 113 602 114 644 645 cell_1rw
* cell instance $18033 r0 *1 16.92,120.12
X$18033 113 603 114 644 645 cell_1rw
* cell instance $18034 m0 *1 16.92,122.85
X$18034 113 604 114 644 645 cell_1rw
* cell instance $18035 r0 *1 16.92,122.85
X$18035 113 605 114 644 645 cell_1rw
* cell instance $18036 m0 *1 16.92,125.58
X$18036 113 606 114 644 645 cell_1rw
* cell instance $18037 r0 *1 16.92,125.58
X$18037 113 607 114 644 645 cell_1rw
* cell instance $18038 m0 *1 16.92,128.31
X$18038 113 609 114 644 645 cell_1rw
* cell instance $18039 r0 *1 16.92,128.31
X$18039 113 608 114 644 645 cell_1rw
* cell instance $18040 m0 *1 16.92,131.04
X$18040 113 610 114 644 645 cell_1rw
* cell instance $18041 r0 *1 16.92,131.04
X$18041 113 611 114 644 645 cell_1rw
* cell instance $18042 m0 *1 16.92,133.77
X$18042 113 612 114 644 645 cell_1rw
* cell instance $18043 r0 *1 16.92,133.77
X$18043 113 613 114 644 645 cell_1rw
* cell instance $18044 m0 *1 16.92,136.5
X$18044 113 615 114 644 645 cell_1rw
* cell instance $18045 r0 *1 16.92,136.5
X$18045 113 614 114 644 645 cell_1rw
* cell instance $18046 m0 *1 16.92,139.23
X$18046 113 617 114 644 645 cell_1rw
* cell instance $18047 r0 *1 16.92,139.23
X$18047 113 616 114 644 645 cell_1rw
* cell instance $18048 m0 *1 16.92,141.96
X$18048 113 618 114 644 645 cell_1rw
* cell instance $18049 r0 *1 16.92,141.96
X$18049 113 619 114 644 645 cell_1rw
* cell instance $18050 m0 *1 16.92,144.69
X$18050 113 620 114 644 645 cell_1rw
* cell instance $18051 r0 *1 16.92,144.69
X$18051 113 621 114 644 645 cell_1rw
* cell instance $18052 m0 *1 16.92,147.42
X$18052 113 622 114 644 645 cell_1rw
* cell instance $18053 r0 *1 16.92,147.42
X$18053 113 623 114 644 645 cell_1rw
* cell instance $18054 m0 *1 16.92,150.15
X$18054 113 624 114 644 645 cell_1rw
* cell instance $18055 r0 *1 16.92,150.15
X$18055 113 625 114 644 645 cell_1rw
* cell instance $18056 m0 *1 16.92,152.88
X$18056 113 626 114 644 645 cell_1rw
* cell instance $18057 r0 *1 16.92,152.88
X$18057 113 627 114 644 645 cell_1rw
* cell instance $18058 m0 *1 16.92,155.61
X$18058 113 628 114 644 645 cell_1rw
* cell instance $18059 r0 *1 16.92,155.61
X$18059 113 629 114 644 645 cell_1rw
* cell instance $18060 m0 *1 16.92,158.34
X$18060 113 630 114 644 645 cell_1rw
* cell instance $18061 r0 *1 16.92,158.34
X$18061 113 631 114 644 645 cell_1rw
* cell instance $18062 m0 *1 16.92,161.07
X$18062 113 632 114 644 645 cell_1rw
* cell instance $18063 r0 *1 16.92,161.07
X$18063 113 633 114 644 645 cell_1rw
* cell instance $18064 m0 *1 16.92,163.8
X$18064 113 634 114 644 645 cell_1rw
* cell instance $18065 r0 *1 16.92,163.8
X$18065 113 635 114 644 645 cell_1rw
* cell instance $18066 m0 *1 16.92,166.53
X$18066 113 637 114 644 645 cell_1rw
* cell instance $18067 r0 *1 16.92,166.53
X$18067 113 636 114 644 645 cell_1rw
* cell instance $18068 m0 *1 16.92,169.26
X$18068 113 639 114 644 645 cell_1rw
* cell instance $18069 r0 *1 16.92,169.26
X$18069 113 638 114 644 645 cell_1rw
* cell instance $18070 m0 *1 16.92,171.99
X$18070 113 640 114 644 645 cell_1rw
* cell instance $18071 r0 *1 16.92,171.99
X$18071 113 641 114 644 645 cell_1rw
* cell instance $18072 m0 *1 16.92,174.72
X$18072 113 642 114 644 645 cell_1rw
* cell instance $18073 r0 *1 16.92,174.72
X$18073 113 643 114 644 645 cell_1rw
* cell instance $18074 m0 *1 17.625,90.09
X$18074 115 581 116 644 645 cell_1rw
* cell instance $18075 r0 *1 17.625,87.36
X$18075 115 322 116 644 645 cell_1rw
* cell instance $18076 m0 *1 17.625,92.82
X$18076 115 583 116 644 645 cell_1rw
* cell instance $18077 r0 *1 17.625,90.09
X$18077 115 580 116 644 645 cell_1rw
* cell instance $18078 r0 *1 17.625,92.82
X$18078 115 582 116 644 645 cell_1rw
* cell instance $18079 m0 *1 17.625,95.55
X$18079 115 584 116 644 645 cell_1rw
* cell instance $18080 r0 *1 17.625,95.55
X$18080 115 585 116 644 645 cell_1rw
* cell instance $18081 m0 *1 17.625,98.28
X$18081 115 586 116 644 645 cell_1rw
* cell instance $18082 r0 *1 17.625,98.28
X$18082 115 587 116 644 645 cell_1rw
* cell instance $18083 m0 *1 17.625,101.01
X$18083 115 588 116 644 645 cell_1rw
* cell instance $18084 r0 *1 17.625,101.01
X$18084 115 589 116 644 645 cell_1rw
* cell instance $18085 m0 *1 17.625,103.74
X$18085 115 590 116 644 645 cell_1rw
* cell instance $18086 r0 *1 17.625,103.74
X$18086 115 591 116 644 645 cell_1rw
* cell instance $18087 m0 *1 17.625,106.47
X$18087 115 593 116 644 645 cell_1rw
* cell instance $18088 r0 *1 17.625,106.47
X$18088 115 592 116 644 645 cell_1rw
* cell instance $18089 m0 *1 17.625,109.2
X$18089 115 594 116 644 645 cell_1rw
* cell instance $18090 r0 *1 17.625,109.2
X$18090 115 595 116 644 645 cell_1rw
* cell instance $18091 m0 *1 17.625,111.93
X$18091 115 597 116 644 645 cell_1rw
* cell instance $18092 r0 *1 17.625,111.93
X$18092 115 596 116 644 645 cell_1rw
* cell instance $18093 m0 *1 17.625,114.66
X$18093 115 598 116 644 645 cell_1rw
* cell instance $18094 m0 *1 17.625,117.39
X$18094 115 600 116 644 645 cell_1rw
* cell instance $18095 r0 *1 17.625,114.66
X$18095 115 599 116 644 645 cell_1rw
* cell instance $18096 m0 *1 17.625,120.12
X$18096 115 602 116 644 645 cell_1rw
* cell instance $18097 r0 *1 17.625,117.39
X$18097 115 601 116 644 645 cell_1rw
* cell instance $18098 r0 *1 17.625,120.12
X$18098 115 603 116 644 645 cell_1rw
* cell instance $18099 m0 *1 17.625,122.85
X$18099 115 604 116 644 645 cell_1rw
* cell instance $18100 r0 *1 17.625,122.85
X$18100 115 605 116 644 645 cell_1rw
* cell instance $18101 m0 *1 17.625,125.58
X$18101 115 606 116 644 645 cell_1rw
* cell instance $18102 r0 *1 17.625,125.58
X$18102 115 607 116 644 645 cell_1rw
* cell instance $18103 m0 *1 17.625,128.31
X$18103 115 609 116 644 645 cell_1rw
* cell instance $18104 m0 *1 17.625,131.04
X$18104 115 610 116 644 645 cell_1rw
* cell instance $18105 r0 *1 17.625,128.31
X$18105 115 608 116 644 645 cell_1rw
* cell instance $18106 r0 *1 17.625,131.04
X$18106 115 611 116 644 645 cell_1rw
* cell instance $18107 m0 *1 17.625,133.77
X$18107 115 612 116 644 645 cell_1rw
* cell instance $18108 r0 *1 17.625,133.77
X$18108 115 613 116 644 645 cell_1rw
* cell instance $18109 m0 *1 17.625,136.5
X$18109 115 615 116 644 645 cell_1rw
* cell instance $18110 r0 *1 17.625,136.5
X$18110 115 614 116 644 645 cell_1rw
* cell instance $18111 m0 *1 17.625,139.23
X$18111 115 617 116 644 645 cell_1rw
* cell instance $18112 r0 *1 17.625,139.23
X$18112 115 616 116 644 645 cell_1rw
* cell instance $18113 m0 *1 17.625,141.96
X$18113 115 618 116 644 645 cell_1rw
* cell instance $18114 r0 *1 17.625,141.96
X$18114 115 619 116 644 645 cell_1rw
* cell instance $18115 m0 *1 17.625,144.69
X$18115 115 620 116 644 645 cell_1rw
* cell instance $18116 r0 *1 17.625,144.69
X$18116 115 621 116 644 645 cell_1rw
* cell instance $18117 m0 *1 17.625,147.42
X$18117 115 622 116 644 645 cell_1rw
* cell instance $18118 r0 *1 17.625,147.42
X$18118 115 623 116 644 645 cell_1rw
* cell instance $18119 m0 *1 17.625,150.15
X$18119 115 624 116 644 645 cell_1rw
* cell instance $18120 r0 *1 17.625,150.15
X$18120 115 625 116 644 645 cell_1rw
* cell instance $18121 m0 *1 17.625,152.88
X$18121 115 626 116 644 645 cell_1rw
* cell instance $18122 r0 *1 17.625,152.88
X$18122 115 627 116 644 645 cell_1rw
* cell instance $18123 m0 *1 17.625,155.61
X$18123 115 628 116 644 645 cell_1rw
* cell instance $18124 r0 *1 17.625,155.61
X$18124 115 629 116 644 645 cell_1rw
* cell instance $18125 m0 *1 17.625,158.34
X$18125 115 630 116 644 645 cell_1rw
* cell instance $18126 r0 *1 17.625,158.34
X$18126 115 631 116 644 645 cell_1rw
* cell instance $18127 m0 *1 17.625,161.07
X$18127 115 632 116 644 645 cell_1rw
* cell instance $18128 r0 *1 17.625,161.07
X$18128 115 633 116 644 645 cell_1rw
* cell instance $18129 m0 *1 17.625,163.8
X$18129 115 634 116 644 645 cell_1rw
* cell instance $18130 r0 *1 17.625,163.8
X$18130 115 635 116 644 645 cell_1rw
* cell instance $18131 m0 *1 17.625,166.53
X$18131 115 637 116 644 645 cell_1rw
* cell instance $18132 r0 *1 17.625,166.53
X$18132 115 636 116 644 645 cell_1rw
* cell instance $18133 m0 *1 17.625,169.26
X$18133 115 639 116 644 645 cell_1rw
* cell instance $18134 m0 *1 17.625,171.99
X$18134 115 640 116 644 645 cell_1rw
* cell instance $18135 r0 *1 17.625,169.26
X$18135 115 638 116 644 645 cell_1rw
* cell instance $18136 r0 *1 17.625,171.99
X$18136 115 641 116 644 645 cell_1rw
* cell instance $18137 m0 *1 17.625,174.72
X$18137 115 642 116 644 645 cell_1rw
* cell instance $18138 r0 *1 17.625,174.72
X$18138 115 643 116 644 645 cell_1rw
* cell instance $18139 r0 *1 18.33,87.36
X$18139 117 322 118 644 645 cell_1rw
* cell instance $18140 m0 *1 18.33,90.09
X$18140 117 581 118 644 645 cell_1rw
* cell instance $18141 m0 *1 18.33,92.82
X$18141 117 583 118 644 645 cell_1rw
* cell instance $18142 r0 *1 18.33,90.09
X$18142 117 580 118 644 645 cell_1rw
* cell instance $18143 r0 *1 18.33,92.82
X$18143 117 582 118 644 645 cell_1rw
* cell instance $18144 m0 *1 18.33,95.55
X$18144 117 584 118 644 645 cell_1rw
* cell instance $18145 m0 *1 18.33,98.28
X$18145 117 586 118 644 645 cell_1rw
* cell instance $18146 r0 *1 18.33,95.55
X$18146 117 585 118 644 645 cell_1rw
* cell instance $18147 r0 *1 18.33,98.28
X$18147 117 587 118 644 645 cell_1rw
* cell instance $18148 m0 *1 18.33,101.01
X$18148 117 588 118 644 645 cell_1rw
* cell instance $18149 r0 *1 18.33,101.01
X$18149 117 589 118 644 645 cell_1rw
* cell instance $18150 m0 *1 18.33,103.74
X$18150 117 590 118 644 645 cell_1rw
* cell instance $18151 r0 *1 18.33,103.74
X$18151 117 591 118 644 645 cell_1rw
* cell instance $18152 m0 *1 18.33,106.47
X$18152 117 593 118 644 645 cell_1rw
* cell instance $18153 m0 *1 18.33,109.2
X$18153 117 594 118 644 645 cell_1rw
* cell instance $18154 r0 *1 18.33,106.47
X$18154 117 592 118 644 645 cell_1rw
* cell instance $18155 r0 *1 18.33,109.2
X$18155 117 595 118 644 645 cell_1rw
* cell instance $18156 m0 *1 18.33,111.93
X$18156 117 597 118 644 645 cell_1rw
* cell instance $18157 r0 *1 18.33,111.93
X$18157 117 596 118 644 645 cell_1rw
* cell instance $18158 m0 *1 18.33,114.66
X$18158 117 598 118 644 645 cell_1rw
* cell instance $18159 r0 *1 18.33,114.66
X$18159 117 599 118 644 645 cell_1rw
* cell instance $18160 m0 *1 18.33,117.39
X$18160 117 600 118 644 645 cell_1rw
* cell instance $18161 r0 *1 18.33,117.39
X$18161 117 601 118 644 645 cell_1rw
* cell instance $18162 m0 *1 18.33,120.12
X$18162 117 602 118 644 645 cell_1rw
* cell instance $18163 r0 *1 18.33,120.12
X$18163 117 603 118 644 645 cell_1rw
* cell instance $18164 m0 *1 18.33,122.85
X$18164 117 604 118 644 645 cell_1rw
* cell instance $18165 r0 *1 18.33,122.85
X$18165 117 605 118 644 645 cell_1rw
* cell instance $18166 m0 *1 18.33,125.58
X$18166 117 606 118 644 645 cell_1rw
* cell instance $18167 r0 *1 18.33,125.58
X$18167 117 607 118 644 645 cell_1rw
* cell instance $18168 m0 *1 18.33,128.31
X$18168 117 609 118 644 645 cell_1rw
* cell instance $18169 r0 *1 18.33,128.31
X$18169 117 608 118 644 645 cell_1rw
* cell instance $18170 m0 *1 18.33,131.04
X$18170 117 610 118 644 645 cell_1rw
* cell instance $18171 r0 *1 18.33,131.04
X$18171 117 611 118 644 645 cell_1rw
* cell instance $18172 m0 *1 18.33,133.77
X$18172 117 612 118 644 645 cell_1rw
* cell instance $18173 r0 *1 18.33,133.77
X$18173 117 613 118 644 645 cell_1rw
* cell instance $18174 m0 *1 18.33,136.5
X$18174 117 615 118 644 645 cell_1rw
* cell instance $18175 m0 *1 18.33,139.23
X$18175 117 617 118 644 645 cell_1rw
* cell instance $18176 r0 *1 18.33,136.5
X$18176 117 614 118 644 645 cell_1rw
* cell instance $18177 r0 *1 18.33,139.23
X$18177 117 616 118 644 645 cell_1rw
* cell instance $18178 m0 *1 18.33,141.96
X$18178 117 618 118 644 645 cell_1rw
* cell instance $18179 r0 *1 18.33,141.96
X$18179 117 619 118 644 645 cell_1rw
* cell instance $18180 m0 *1 18.33,144.69
X$18180 117 620 118 644 645 cell_1rw
* cell instance $18181 r0 *1 18.33,144.69
X$18181 117 621 118 644 645 cell_1rw
* cell instance $18182 m0 *1 18.33,147.42
X$18182 117 622 118 644 645 cell_1rw
* cell instance $18183 r0 *1 18.33,147.42
X$18183 117 623 118 644 645 cell_1rw
* cell instance $18184 m0 *1 18.33,150.15
X$18184 117 624 118 644 645 cell_1rw
* cell instance $18185 r0 *1 18.33,150.15
X$18185 117 625 118 644 645 cell_1rw
* cell instance $18186 m0 *1 18.33,152.88
X$18186 117 626 118 644 645 cell_1rw
* cell instance $18187 r0 *1 18.33,152.88
X$18187 117 627 118 644 645 cell_1rw
* cell instance $18188 m0 *1 18.33,155.61
X$18188 117 628 118 644 645 cell_1rw
* cell instance $18189 r0 *1 18.33,155.61
X$18189 117 629 118 644 645 cell_1rw
* cell instance $18190 m0 *1 18.33,158.34
X$18190 117 630 118 644 645 cell_1rw
* cell instance $18191 r0 *1 18.33,158.34
X$18191 117 631 118 644 645 cell_1rw
* cell instance $18192 m0 *1 18.33,161.07
X$18192 117 632 118 644 645 cell_1rw
* cell instance $18193 r0 *1 18.33,161.07
X$18193 117 633 118 644 645 cell_1rw
* cell instance $18194 m0 *1 18.33,163.8
X$18194 117 634 118 644 645 cell_1rw
* cell instance $18195 r0 *1 18.33,163.8
X$18195 117 635 118 644 645 cell_1rw
* cell instance $18196 m0 *1 18.33,166.53
X$18196 117 637 118 644 645 cell_1rw
* cell instance $18197 r0 *1 18.33,166.53
X$18197 117 636 118 644 645 cell_1rw
* cell instance $18198 m0 *1 18.33,169.26
X$18198 117 639 118 644 645 cell_1rw
* cell instance $18199 r0 *1 18.33,169.26
X$18199 117 638 118 644 645 cell_1rw
* cell instance $18200 m0 *1 18.33,171.99
X$18200 117 640 118 644 645 cell_1rw
* cell instance $18201 r0 *1 18.33,171.99
X$18201 117 641 118 644 645 cell_1rw
* cell instance $18202 m0 *1 18.33,174.72
X$18202 117 642 118 644 645 cell_1rw
* cell instance $18203 r0 *1 18.33,174.72
X$18203 117 643 118 644 645 cell_1rw
* cell instance $18204 r0 *1 19.035,87.36
X$18204 119 322 120 644 645 cell_1rw
* cell instance $18205 m0 *1 19.035,90.09
X$18205 119 581 120 644 645 cell_1rw
* cell instance $18206 r0 *1 19.035,90.09
X$18206 119 580 120 644 645 cell_1rw
* cell instance $18207 m0 *1 19.035,92.82
X$18207 119 583 120 644 645 cell_1rw
* cell instance $18208 r0 *1 19.035,92.82
X$18208 119 582 120 644 645 cell_1rw
* cell instance $18209 m0 *1 19.035,95.55
X$18209 119 584 120 644 645 cell_1rw
* cell instance $18210 r0 *1 19.035,95.55
X$18210 119 585 120 644 645 cell_1rw
* cell instance $18211 m0 *1 19.035,98.28
X$18211 119 586 120 644 645 cell_1rw
* cell instance $18212 r0 *1 19.035,98.28
X$18212 119 587 120 644 645 cell_1rw
* cell instance $18213 m0 *1 19.035,101.01
X$18213 119 588 120 644 645 cell_1rw
* cell instance $18214 r0 *1 19.035,101.01
X$18214 119 589 120 644 645 cell_1rw
* cell instance $18215 m0 *1 19.035,103.74
X$18215 119 590 120 644 645 cell_1rw
* cell instance $18216 r0 *1 19.035,103.74
X$18216 119 591 120 644 645 cell_1rw
* cell instance $18217 m0 *1 19.035,106.47
X$18217 119 593 120 644 645 cell_1rw
* cell instance $18218 m0 *1 19.035,109.2
X$18218 119 594 120 644 645 cell_1rw
* cell instance $18219 r0 *1 19.035,106.47
X$18219 119 592 120 644 645 cell_1rw
* cell instance $18220 r0 *1 19.035,109.2
X$18220 119 595 120 644 645 cell_1rw
* cell instance $18221 m0 *1 19.035,111.93
X$18221 119 597 120 644 645 cell_1rw
* cell instance $18222 r0 *1 19.035,111.93
X$18222 119 596 120 644 645 cell_1rw
* cell instance $18223 m0 *1 19.035,114.66
X$18223 119 598 120 644 645 cell_1rw
* cell instance $18224 r0 *1 19.035,114.66
X$18224 119 599 120 644 645 cell_1rw
* cell instance $18225 m0 *1 19.035,117.39
X$18225 119 600 120 644 645 cell_1rw
* cell instance $18226 r0 *1 19.035,117.39
X$18226 119 601 120 644 645 cell_1rw
* cell instance $18227 m0 *1 19.035,120.12
X$18227 119 602 120 644 645 cell_1rw
* cell instance $18228 r0 *1 19.035,120.12
X$18228 119 603 120 644 645 cell_1rw
* cell instance $18229 m0 *1 19.035,122.85
X$18229 119 604 120 644 645 cell_1rw
* cell instance $18230 r0 *1 19.035,122.85
X$18230 119 605 120 644 645 cell_1rw
* cell instance $18231 m0 *1 19.035,125.58
X$18231 119 606 120 644 645 cell_1rw
* cell instance $18232 r0 *1 19.035,125.58
X$18232 119 607 120 644 645 cell_1rw
* cell instance $18233 m0 *1 19.035,128.31
X$18233 119 609 120 644 645 cell_1rw
* cell instance $18234 m0 *1 19.035,131.04
X$18234 119 610 120 644 645 cell_1rw
* cell instance $18235 r0 *1 19.035,128.31
X$18235 119 608 120 644 645 cell_1rw
* cell instance $18236 r0 *1 19.035,131.04
X$18236 119 611 120 644 645 cell_1rw
* cell instance $18237 m0 *1 19.035,133.77
X$18237 119 612 120 644 645 cell_1rw
* cell instance $18238 r0 *1 19.035,133.77
X$18238 119 613 120 644 645 cell_1rw
* cell instance $18239 m0 *1 19.035,136.5
X$18239 119 615 120 644 645 cell_1rw
* cell instance $18240 r0 *1 19.035,136.5
X$18240 119 614 120 644 645 cell_1rw
* cell instance $18241 m0 *1 19.035,139.23
X$18241 119 617 120 644 645 cell_1rw
* cell instance $18242 r0 *1 19.035,139.23
X$18242 119 616 120 644 645 cell_1rw
* cell instance $18243 m0 *1 19.035,141.96
X$18243 119 618 120 644 645 cell_1rw
* cell instance $18244 r0 *1 19.035,141.96
X$18244 119 619 120 644 645 cell_1rw
* cell instance $18245 m0 *1 19.035,144.69
X$18245 119 620 120 644 645 cell_1rw
* cell instance $18246 m0 *1 19.035,147.42
X$18246 119 622 120 644 645 cell_1rw
* cell instance $18247 r0 *1 19.035,144.69
X$18247 119 621 120 644 645 cell_1rw
* cell instance $18248 r0 *1 19.035,147.42
X$18248 119 623 120 644 645 cell_1rw
* cell instance $18249 m0 *1 19.035,150.15
X$18249 119 624 120 644 645 cell_1rw
* cell instance $18250 r0 *1 19.035,150.15
X$18250 119 625 120 644 645 cell_1rw
* cell instance $18251 m0 *1 19.035,152.88
X$18251 119 626 120 644 645 cell_1rw
* cell instance $18252 r0 *1 19.035,152.88
X$18252 119 627 120 644 645 cell_1rw
* cell instance $18253 m0 *1 19.035,155.61
X$18253 119 628 120 644 645 cell_1rw
* cell instance $18254 r0 *1 19.035,155.61
X$18254 119 629 120 644 645 cell_1rw
* cell instance $18255 m0 *1 19.035,158.34
X$18255 119 630 120 644 645 cell_1rw
* cell instance $18256 r0 *1 19.035,158.34
X$18256 119 631 120 644 645 cell_1rw
* cell instance $18257 m0 *1 19.035,161.07
X$18257 119 632 120 644 645 cell_1rw
* cell instance $18258 r0 *1 19.035,161.07
X$18258 119 633 120 644 645 cell_1rw
* cell instance $18259 m0 *1 19.035,163.8
X$18259 119 634 120 644 645 cell_1rw
* cell instance $18260 r0 *1 19.035,163.8
X$18260 119 635 120 644 645 cell_1rw
* cell instance $18261 m0 *1 19.035,166.53
X$18261 119 637 120 644 645 cell_1rw
* cell instance $18262 r0 *1 19.035,166.53
X$18262 119 636 120 644 645 cell_1rw
* cell instance $18263 m0 *1 19.035,169.26
X$18263 119 639 120 644 645 cell_1rw
* cell instance $18264 r0 *1 19.035,169.26
X$18264 119 638 120 644 645 cell_1rw
* cell instance $18265 m0 *1 19.035,171.99
X$18265 119 640 120 644 645 cell_1rw
* cell instance $18266 r0 *1 19.035,171.99
X$18266 119 641 120 644 645 cell_1rw
* cell instance $18267 m0 *1 19.035,174.72
X$18267 119 642 120 644 645 cell_1rw
* cell instance $18268 r0 *1 19.035,174.72
X$18268 119 643 120 644 645 cell_1rw
* cell instance $18269 r0 *1 19.74,87.36
X$18269 121 322 122 644 645 cell_1rw
* cell instance $18270 m0 *1 19.74,90.09
X$18270 121 581 122 644 645 cell_1rw
* cell instance $18271 r0 *1 19.74,90.09
X$18271 121 580 122 644 645 cell_1rw
* cell instance $18272 m0 *1 19.74,92.82
X$18272 121 583 122 644 645 cell_1rw
* cell instance $18273 r0 *1 19.74,92.82
X$18273 121 582 122 644 645 cell_1rw
* cell instance $18274 m0 *1 19.74,95.55
X$18274 121 584 122 644 645 cell_1rw
* cell instance $18275 r0 *1 19.74,95.55
X$18275 121 585 122 644 645 cell_1rw
* cell instance $18276 m0 *1 19.74,98.28
X$18276 121 586 122 644 645 cell_1rw
* cell instance $18277 r0 *1 19.74,98.28
X$18277 121 587 122 644 645 cell_1rw
* cell instance $18278 m0 *1 19.74,101.01
X$18278 121 588 122 644 645 cell_1rw
* cell instance $18279 r0 *1 19.74,101.01
X$18279 121 589 122 644 645 cell_1rw
* cell instance $18280 m0 *1 19.74,103.74
X$18280 121 590 122 644 645 cell_1rw
* cell instance $18281 r0 *1 19.74,103.74
X$18281 121 591 122 644 645 cell_1rw
* cell instance $18282 m0 *1 19.74,106.47
X$18282 121 593 122 644 645 cell_1rw
* cell instance $18283 r0 *1 19.74,106.47
X$18283 121 592 122 644 645 cell_1rw
* cell instance $18284 m0 *1 19.74,109.2
X$18284 121 594 122 644 645 cell_1rw
* cell instance $18285 r0 *1 19.74,109.2
X$18285 121 595 122 644 645 cell_1rw
* cell instance $18286 m0 *1 19.74,111.93
X$18286 121 597 122 644 645 cell_1rw
* cell instance $18287 r0 *1 19.74,111.93
X$18287 121 596 122 644 645 cell_1rw
* cell instance $18288 m0 *1 19.74,114.66
X$18288 121 598 122 644 645 cell_1rw
* cell instance $18289 r0 *1 19.74,114.66
X$18289 121 599 122 644 645 cell_1rw
* cell instance $18290 m0 *1 19.74,117.39
X$18290 121 600 122 644 645 cell_1rw
* cell instance $18291 r0 *1 19.74,117.39
X$18291 121 601 122 644 645 cell_1rw
* cell instance $18292 m0 *1 19.74,120.12
X$18292 121 602 122 644 645 cell_1rw
* cell instance $18293 r0 *1 19.74,120.12
X$18293 121 603 122 644 645 cell_1rw
* cell instance $18294 m0 *1 19.74,122.85
X$18294 121 604 122 644 645 cell_1rw
* cell instance $18295 r0 *1 19.74,122.85
X$18295 121 605 122 644 645 cell_1rw
* cell instance $18296 m0 *1 19.74,125.58
X$18296 121 606 122 644 645 cell_1rw
* cell instance $18297 r0 *1 19.74,125.58
X$18297 121 607 122 644 645 cell_1rw
* cell instance $18298 m0 *1 19.74,128.31
X$18298 121 609 122 644 645 cell_1rw
* cell instance $18299 m0 *1 19.74,131.04
X$18299 121 610 122 644 645 cell_1rw
* cell instance $18300 r0 *1 19.74,128.31
X$18300 121 608 122 644 645 cell_1rw
* cell instance $18301 r0 *1 19.74,131.04
X$18301 121 611 122 644 645 cell_1rw
* cell instance $18302 m0 *1 19.74,133.77
X$18302 121 612 122 644 645 cell_1rw
* cell instance $18303 m0 *1 19.74,136.5
X$18303 121 615 122 644 645 cell_1rw
* cell instance $18304 r0 *1 19.74,133.77
X$18304 121 613 122 644 645 cell_1rw
* cell instance $18305 r0 *1 19.74,136.5
X$18305 121 614 122 644 645 cell_1rw
* cell instance $18306 m0 *1 19.74,139.23
X$18306 121 617 122 644 645 cell_1rw
* cell instance $18307 r0 *1 19.74,139.23
X$18307 121 616 122 644 645 cell_1rw
* cell instance $18308 m0 *1 19.74,141.96
X$18308 121 618 122 644 645 cell_1rw
* cell instance $18309 r0 *1 19.74,141.96
X$18309 121 619 122 644 645 cell_1rw
* cell instance $18310 m0 *1 19.74,144.69
X$18310 121 620 122 644 645 cell_1rw
* cell instance $18311 r0 *1 19.74,144.69
X$18311 121 621 122 644 645 cell_1rw
* cell instance $18312 m0 *1 19.74,147.42
X$18312 121 622 122 644 645 cell_1rw
* cell instance $18313 m0 *1 19.74,150.15
X$18313 121 624 122 644 645 cell_1rw
* cell instance $18314 r0 *1 19.74,147.42
X$18314 121 623 122 644 645 cell_1rw
* cell instance $18315 r0 *1 19.74,150.15
X$18315 121 625 122 644 645 cell_1rw
* cell instance $18316 m0 *1 19.74,152.88
X$18316 121 626 122 644 645 cell_1rw
* cell instance $18317 r0 *1 19.74,152.88
X$18317 121 627 122 644 645 cell_1rw
* cell instance $18318 m0 *1 19.74,155.61
X$18318 121 628 122 644 645 cell_1rw
* cell instance $18319 r0 *1 19.74,155.61
X$18319 121 629 122 644 645 cell_1rw
* cell instance $18320 m0 *1 19.74,158.34
X$18320 121 630 122 644 645 cell_1rw
* cell instance $18321 r0 *1 19.74,158.34
X$18321 121 631 122 644 645 cell_1rw
* cell instance $18322 m0 *1 19.74,161.07
X$18322 121 632 122 644 645 cell_1rw
* cell instance $18323 m0 *1 19.74,163.8
X$18323 121 634 122 644 645 cell_1rw
* cell instance $18324 r0 *1 19.74,161.07
X$18324 121 633 122 644 645 cell_1rw
* cell instance $18325 r0 *1 19.74,163.8
X$18325 121 635 122 644 645 cell_1rw
* cell instance $18326 m0 *1 19.74,166.53
X$18326 121 637 122 644 645 cell_1rw
* cell instance $18327 r0 *1 19.74,166.53
X$18327 121 636 122 644 645 cell_1rw
* cell instance $18328 m0 *1 19.74,169.26
X$18328 121 639 122 644 645 cell_1rw
* cell instance $18329 r0 *1 19.74,169.26
X$18329 121 638 122 644 645 cell_1rw
* cell instance $18330 m0 *1 19.74,171.99
X$18330 121 640 122 644 645 cell_1rw
* cell instance $18331 r0 *1 19.74,171.99
X$18331 121 641 122 644 645 cell_1rw
* cell instance $18332 m0 *1 19.74,174.72
X$18332 121 642 122 644 645 cell_1rw
* cell instance $18333 r0 *1 19.74,174.72
X$18333 121 643 122 644 645 cell_1rw
* cell instance $18334 r0 *1 20.445,87.36
X$18334 123 322 124 644 645 cell_1rw
* cell instance $18335 m0 *1 20.445,90.09
X$18335 123 581 124 644 645 cell_1rw
* cell instance $18336 r0 *1 20.445,90.09
X$18336 123 580 124 644 645 cell_1rw
* cell instance $18337 m0 *1 20.445,92.82
X$18337 123 583 124 644 645 cell_1rw
* cell instance $18338 r0 *1 20.445,92.82
X$18338 123 582 124 644 645 cell_1rw
* cell instance $18339 m0 *1 20.445,95.55
X$18339 123 584 124 644 645 cell_1rw
* cell instance $18340 r0 *1 20.445,95.55
X$18340 123 585 124 644 645 cell_1rw
* cell instance $18341 m0 *1 20.445,98.28
X$18341 123 586 124 644 645 cell_1rw
* cell instance $18342 r0 *1 20.445,98.28
X$18342 123 587 124 644 645 cell_1rw
* cell instance $18343 m0 *1 20.445,101.01
X$18343 123 588 124 644 645 cell_1rw
* cell instance $18344 r0 *1 20.445,101.01
X$18344 123 589 124 644 645 cell_1rw
* cell instance $18345 m0 *1 20.445,103.74
X$18345 123 590 124 644 645 cell_1rw
* cell instance $18346 r0 *1 20.445,103.74
X$18346 123 591 124 644 645 cell_1rw
* cell instance $18347 m0 *1 20.445,106.47
X$18347 123 593 124 644 645 cell_1rw
* cell instance $18348 r0 *1 20.445,106.47
X$18348 123 592 124 644 645 cell_1rw
* cell instance $18349 m0 *1 20.445,109.2
X$18349 123 594 124 644 645 cell_1rw
* cell instance $18350 r0 *1 20.445,109.2
X$18350 123 595 124 644 645 cell_1rw
* cell instance $18351 m0 *1 20.445,111.93
X$18351 123 597 124 644 645 cell_1rw
* cell instance $18352 r0 *1 20.445,111.93
X$18352 123 596 124 644 645 cell_1rw
* cell instance $18353 m0 *1 20.445,114.66
X$18353 123 598 124 644 645 cell_1rw
* cell instance $18354 m0 *1 20.445,117.39
X$18354 123 600 124 644 645 cell_1rw
* cell instance $18355 r0 *1 20.445,114.66
X$18355 123 599 124 644 645 cell_1rw
* cell instance $18356 r0 *1 20.445,117.39
X$18356 123 601 124 644 645 cell_1rw
* cell instance $18357 m0 *1 20.445,120.12
X$18357 123 602 124 644 645 cell_1rw
* cell instance $18358 r0 *1 20.445,120.12
X$18358 123 603 124 644 645 cell_1rw
* cell instance $18359 m0 *1 20.445,122.85
X$18359 123 604 124 644 645 cell_1rw
* cell instance $18360 r0 *1 20.445,122.85
X$18360 123 605 124 644 645 cell_1rw
* cell instance $18361 m0 *1 20.445,125.58
X$18361 123 606 124 644 645 cell_1rw
* cell instance $18362 r0 *1 20.445,125.58
X$18362 123 607 124 644 645 cell_1rw
* cell instance $18363 m0 *1 20.445,128.31
X$18363 123 609 124 644 645 cell_1rw
* cell instance $18364 m0 *1 20.445,131.04
X$18364 123 610 124 644 645 cell_1rw
* cell instance $18365 r0 *1 20.445,128.31
X$18365 123 608 124 644 645 cell_1rw
* cell instance $18366 r0 *1 20.445,131.04
X$18366 123 611 124 644 645 cell_1rw
* cell instance $18367 m0 *1 20.445,133.77
X$18367 123 612 124 644 645 cell_1rw
* cell instance $18368 r0 *1 20.445,133.77
X$18368 123 613 124 644 645 cell_1rw
* cell instance $18369 m0 *1 20.445,136.5
X$18369 123 615 124 644 645 cell_1rw
* cell instance $18370 m0 *1 20.445,139.23
X$18370 123 617 124 644 645 cell_1rw
* cell instance $18371 r0 *1 20.445,136.5
X$18371 123 614 124 644 645 cell_1rw
* cell instance $18372 r0 *1 20.445,139.23
X$18372 123 616 124 644 645 cell_1rw
* cell instance $18373 m0 *1 20.445,141.96
X$18373 123 618 124 644 645 cell_1rw
* cell instance $18374 r0 *1 20.445,141.96
X$18374 123 619 124 644 645 cell_1rw
* cell instance $18375 m0 *1 20.445,144.69
X$18375 123 620 124 644 645 cell_1rw
* cell instance $18376 r0 *1 20.445,144.69
X$18376 123 621 124 644 645 cell_1rw
* cell instance $18377 m0 *1 20.445,147.42
X$18377 123 622 124 644 645 cell_1rw
* cell instance $18378 r0 *1 20.445,147.42
X$18378 123 623 124 644 645 cell_1rw
* cell instance $18379 m0 *1 20.445,150.15
X$18379 123 624 124 644 645 cell_1rw
* cell instance $18380 r0 *1 20.445,150.15
X$18380 123 625 124 644 645 cell_1rw
* cell instance $18381 m0 *1 20.445,152.88
X$18381 123 626 124 644 645 cell_1rw
* cell instance $18382 r0 *1 20.445,152.88
X$18382 123 627 124 644 645 cell_1rw
* cell instance $18383 m0 *1 20.445,155.61
X$18383 123 628 124 644 645 cell_1rw
* cell instance $18384 r0 *1 20.445,155.61
X$18384 123 629 124 644 645 cell_1rw
* cell instance $18385 m0 *1 20.445,158.34
X$18385 123 630 124 644 645 cell_1rw
* cell instance $18386 r0 *1 20.445,158.34
X$18386 123 631 124 644 645 cell_1rw
* cell instance $18387 m0 *1 20.445,161.07
X$18387 123 632 124 644 645 cell_1rw
* cell instance $18388 r0 *1 20.445,161.07
X$18388 123 633 124 644 645 cell_1rw
* cell instance $18389 m0 *1 20.445,163.8
X$18389 123 634 124 644 645 cell_1rw
* cell instance $18390 r0 *1 20.445,163.8
X$18390 123 635 124 644 645 cell_1rw
* cell instance $18391 m0 *1 20.445,166.53
X$18391 123 637 124 644 645 cell_1rw
* cell instance $18392 r0 *1 20.445,166.53
X$18392 123 636 124 644 645 cell_1rw
* cell instance $18393 m0 *1 20.445,169.26
X$18393 123 639 124 644 645 cell_1rw
* cell instance $18394 r0 *1 20.445,169.26
X$18394 123 638 124 644 645 cell_1rw
* cell instance $18395 m0 *1 20.445,171.99
X$18395 123 640 124 644 645 cell_1rw
* cell instance $18396 r0 *1 20.445,171.99
X$18396 123 641 124 644 645 cell_1rw
* cell instance $18397 m0 *1 20.445,174.72
X$18397 123 642 124 644 645 cell_1rw
* cell instance $18398 r0 *1 20.445,174.72
X$18398 123 643 124 644 645 cell_1rw
* cell instance $18399 r0 *1 21.15,87.36
X$18399 125 322 126 644 645 cell_1rw
* cell instance $18400 m0 *1 21.15,90.09
X$18400 125 581 126 644 645 cell_1rw
* cell instance $18401 r0 *1 21.15,90.09
X$18401 125 580 126 644 645 cell_1rw
* cell instance $18402 m0 *1 21.15,92.82
X$18402 125 583 126 644 645 cell_1rw
* cell instance $18403 r0 *1 21.15,92.82
X$18403 125 582 126 644 645 cell_1rw
* cell instance $18404 m0 *1 21.15,95.55
X$18404 125 584 126 644 645 cell_1rw
* cell instance $18405 r0 *1 21.15,95.55
X$18405 125 585 126 644 645 cell_1rw
* cell instance $18406 m0 *1 21.15,98.28
X$18406 125 586 126 644 645 cell_1rw
* cell instance $18407 r0 *1 21.15,98.28
X$18407 125 587 126 644 645 cell_1rw
* cell instance $18408 m0 *1 21.15,101.01
X$18408 125 588 126 644 645 cell_1rw
* cell instance $18409 r0 *1 21.15,101.01
X$18409 125 589 126 644 645 cell_1rw
* cell instance $18410 m0 *1 21.15,103.74
X$18410 125 590 126 644 645 cell_1rw
* cell instance $18411 r0 *1 21.15,103.74
X$18411 125 591 126 644 645 cell_1rw
* cell instance $18412 m0 *1 21.15,106.47
X$18412 125 593 126 644 645 cell_1rw
* cell instance $18413 m0 *1 21.15,109.2
X$18413 125 594 126 644 645 cell_1rw
* cell instance $18414 r0 *1 21.15,106.47
X$18414 125 592 126 644 645 cell_1rw
* cell instance $18415 r0 *1 21.15,109.2
X$18415 125 595 126 644 645 cell_1rw
* cell instance $18416 m0 *1 21.15,111.93
X$18416 125 597 126 644 645 cell_1rw
* cell instance $18417 r0 *1 21.15,111.93
X$18417 125 596 126 644 645 cell_1rw
* cell instance $18418 m0 *1 21.15,114.66
X$18418 125 598 126 644 645 cell_1rw
* cell instance $18419 r0 *1 21.15,114.66
X$18419 125 599 126 644 645 cell_1rw
* cell instance $18420 m0 *1 21.15,117.39
X$18420 125 600 126 644 645 cell_1rw
* cell instance $18421 r0 *1 21.15,117.39
X$18421 125 601 126 644 645 cell_1rw
* cell instance $18422 m0 *1 21.15,120.12
X$18422 125 602 126 644 645 cell_1rw
* cell instance $18423 r0 *1 21.15,120.12
X$18423 125 603 126 644 645 cell_1rw
* cell instance $18424 m0 *1 21.15,122.85
X$18424 125 604 126 644 645 cell_1rw
* cell instance $18425 r0 *1 21.15,122.85
X$18425 125 605 126 644 645 cell_1rw
* cell instance $18426 m0 *1 21.15,125.58
X$18426 125 606 126 644 645 cell_1rw
* cell instance $18427 r0 *1 21.15,125.58
X$18427 125 607 126 644 645 cell_1rw
* cell instance $18428 m0 *1 21.15,128.31
X$18428 125 609 126 644 645 cell_1rw
* cell instance $18429 r0 *1 21.15,128.31
X$18429 125 608 126 644 645 cell_1rw
* cell instance $18430 m0 *1 21.15,131.04
X$18430 125 610 126 644 645 cell_1rw
* cell instance $18431 r0 *1 21.15,131.04
X$18431 125 611 126 644 645 cell_1rw
* cell instance $18432 m0 *1 21.15,133.77
X$18432 125 612 126 644 645 cell_1rw
* cell instance $18433 r0 *1 21.15,133.77
X$18433 125 613 126 644 645 cell_1rw
* cell instance $18434 m0 *1 21.15,136.5
X$18434 125 615 126 644 645 cell_1rw
* cell instance $18435 r0 *1 21.15,136.5
X$18435 125 614 126 644 645 cell_1rw
* cell instance $18436 m0 *1 21.15,139.23
X$18436 125 617 126 644 645 cell_1rw
* cell instance $18437 r0 *1 21.15,139.23
X$18437 125 616 126 644 645 cell_1rw
* cell instance $18438 m0 *1 21.15,141.96
X$18438 125 618 126 644 645 cell_1rw
* cell instance $18439 r0 *1 21.15,141.96
X$18439 125 619 126 644 645 cell_1rw
* cell instance $18440 m0 *1 21.15,144.69
X$18440 125 620 126 644 645 cell_1rw
* cell instance $18441 r0 *1 21.15,144.69
X$18441 125 621 126 644 645 cell_1rw
* cell instance $18442 m0 *1 21.15,147.42
X$18442 125 622 126 644 645 cell_1rw
* cell instance $18443 m0 *1 21.15,150.15
X$18443 125 624 126 644 645 cell_1rw
* cell instance $18444 r0 *1 21.15,147.42
X$18444 125 623 126 644 645 cell_1rw
* cell instance $18445 r0 *1 21.15,150.15
X$18445 125 625 126 644 645 cell_1rw
* cell instance $18446 m0 *1 21.15,152.88
X$18446 125 626 126 644 645 cell_1rw
* cell instance $18447 r0 *1 21.15,152.88
X$18447 125 627 126 644 645 cell_1rw
* cell instance $18448 m0 *1 21.15,155.61
X$18448 125 628 126 644 645 cell_1rw
* cell instance $18449 r0 *1 21.15,155.61
X$18449 125 629 126 644 645 cell_1rw
* cell instance $18450 m0 *1 21.15,158.34
X$18450 125 630 126 644 645 cell_1rw
* cell instance $18451 r0 *1 21.15,158.34
X$18451 125 631 126 644 645 cell_1rw
* cell instance $18452 m0 *1 21.15,161.07
X$18452 125 632 126 644 645 cell_1rw
* cell instance $18453 r0 *1 21.15,161.07
X$18453 125 633 126 644 645 cell_1rw
* cell instance $18454 m0 *1 21.15,163.8
X$18454 125 634 126 644 645 cell_1rw
* cell instance $18455 r0 *1 21.15,163.8
X$18455 125 635 126 644 645 cell_1rw
* cell instance $18456 m0 *1 21.15,166.53
X$18456 125 637 126 644 645 cell_1rw
* cell instance $18457 m0 *1 21.15,169.26
X$18457 125 639 126 644 645 cell_1rw
* cell instance $18458 r0 *1 21.15,166.53
X$18458 125 636 126 644 645 cell_1rw
* cell instance $18459 m0 *1 21.15,171.99
X$18459 125 640 126 644 645 cell_1rw
* cell instance $18460 r0 *1 21.15,169.26
X$18460 125 638 126 644 645 cell_1rw
* cell instance $18461 r0 *1 21.15,171.99
X$18461 125 641 126 644 645 cell_1rw
* cell instance $18462 m0 *1 21.15,174.72
X$18462 125 642 126 644 645 cell_1rw
* cell instance $18463 r0 *1 21.15,174.72
X$18463 125 643 126 644 645 cell_1rw
* cell instance $18464 r0 *1 21.855,87.36
X$18464 127 322 128 644 645 cell_1rw
* cell instance $18465 m0 *1 21.855,90.09
X$18465 127 581 128 644 645 cell_1rw
* cell instance $18466 m0 *1 21.855,92.82
X$18466 127 583 128 644 645 cell_1rw
* cell instance $18467 r0 *1 21.855,90.09
X$18467 127 580 128 644 645 cell_1rw
* cell instance $18468 r0 *1 21.855,92.82
X$18468 127 582 128 644 645 cell_1rw
* cell instance $18469 m0 *1 21.855,95.55
X$18469 127 584 128 644 645 cell_1rw
* cell instance $18470 r0 *1 21.855,95.55
X$18470 127 585 128 644 645 cell_1rw
* cell instance $18471 m0 *1 21.855,98.28
X$18471 127 586 128 644 645 cell_1rw
* cell instance $18472 r0 *1 21.855,98.28
X$18472 127 587 128 644 645 cell_1rw
* cell instance $18473 m0 *1 21.855,101.01
X$18473 127 588 128 644 645 cell_1rw
* cell instance $18474 r0 *1 21.855,101.01
X$18474 127 589 128 644 645 cell_1rw
* cell instance $18475 m0 *1 21.855,103.74
X$18475 127 590 128 644 645 cell_1rw
* cell instance $18476 r0 *1 21.855,103.74
X$18476 127 591 128 644 645 cell_1rw
* cell instance $18477 m0 *1 21.855,106.47
X$18477 127 593 128 644 645 cell_1rw
* cell instance $18478 r0 *1 21.855,106.47
X$18478 127 592 128 644 645 cell_1rw
* cell instance $18479 m0 *1 21.855,109.2
X$18479 127 594 128 644 645 cell_1rw
* cell instance $18480 r0 *1 21.855,109.2
X$18480 127 595 128 644 645 cell_1rw
* cell instance $18481 m0 *1 21.855,111.93
X$18481 127 597 128 644 645 cell_1rw
* cell instance $18482 r0 *1 21.855,111.93
X$18482 127 596 128 644 645 cell_1rw
* cell instance $18483 m0 *1 21.855,114.66
X$18483 127 598 128 644 645 cell_1rw
* cell instance $18484 r0 *1 21.855,114.66
X$18484 127 599 128 644 645 cell_1rw
* cell instance $18485 m0 *1 21.855,117.39
X$18485 127 600 128 644 645 cell_1rw
* cell instance $18486 r0 *1 21.855,117.39
X$18486 127 601 128 644 645 cell_1rw
* cell instance $18487 m0 *1 21.855,120.12
X$18487 127 602 128 644 645 cell_1rw
* cell instance $18488 r0 *1 21.855,120.12
X$18488 127 603 128 644 645 cell_1rw
* cell instance $18489 m0 *1 21.855,122.85
X$18489 127 604 128 644 645 cell_1rw
* cell instance $18490 r0 *1 21.855,122.85
X$18490 127 605 128 644 645 cell_1rw
* cell instance $18491 m0 *1 21.855,125.58
X$18491 127 606 128 644 645 cell_1rw
* cell instance $18492 r0 *1 21.855,125.58
X$18492 127 607 128 644 645 cell_1rw
* cell instance $18493 m0 *1 21.855,128.31
X$18493 127 609 128 644 645 cell_1rw
* cell instance $18494 r0 *1 21.855,128.31
X$18494 127 608 128 644 645 cell_1rw
* cell instance $18495 m0 *1 21.855,131.04
X$18495 127 610 128 644 645 cell_1rw
* cell instance $18496 r0 *1 21.855,131.04
X$18496 127 611 128 644 645 cell_1rw
* cell instance $18497 m0 *1 21.855,133.77
X$18497 127 612 128 644 645 cell_1rw
* cell instance $18498 r0 *1 21.855,133.77
X$18498 127 613 128 644 645 cell_1rw
* cell instance $18499 m0 *1 21.855,136.5
X$18499 127 615 128 644 645 cell_1rw
* cell instance $18500 r0 *1 21.855,136.5
X$18500 127 614 128 644 645 cell_1rw
* cell instance $18501 m0 *1 21.855,139.23
X$18501 127 617 128 644 645 cell_1rw
* cell instance $18502 r0 *1 21.855,139.23
X$18502 127 616 128 644 645 cell_1rw
* cell instance $18503 m0 *1 21.855,141.96
X$18503 127 618 128 644 645 cell_1rw
* cell instance $18504 r0 *1 21.855,141.96
X$18504 127 619 128 644 645 cell_1rw
* cell instance $18505 m0 *1 21.855,144.69
X$18505 127 620 128 644 645 cell_1rw
* cell instance $18506 r0 *1 21.855,144.69
X$18506 127 621 128 644 645 cell_1rw
* cell instance $18507 m0 *1 21.855,147.42
X$18507 127 622 128 644 645 cell_1rw
* cell instance $18508 r0 *1 21.855,147.42
X$18508 127 623 128 644 645 cell_1rw
* cell instance $18509 m0 *1 21.855,150.15
X$18509 127 624 128 644 645 cell_1rw
* cell instance $18510 r0 *1 21.855,150.15
X$18510 127 625 128 644 645 cell_1rw
* cell instance $18511 m0 *1 21.855,152.88
X$18511 127 626 128 644 645 cell_1rw
* cell instance $18512 r0 *1 21.855,152.88
X$18512 127 627 128 644 645 cell_1rw
* cell instance $18513 m0 *1 21.855,155.61
X$18513 127 628 128 644 645 cell_1rw
* cell instance $18514 r0 *1 21.855,155.61
X$18514 127 629 128 644 645 cell_1rw
* cell instance $18515 m0 *1 21.855,158.34
X$18515 127 630 128 644 645 cell_1rw
* cell instance $18516 r0 *1 21.855,158.34
X$18516 127 631 128 644 645 cell_1rw
* cell instance $18517 m0 *1 21.855,161.07
X$18517 127 632 128 644 645 cell_1rw
* cell instance $18518 r0 *1 21.855,161.07
X$18518 127 633 128 644 645 cell_1rw
* cell instance $18519 m0 *1 21.855,163.8
X$18519 127 634 128 644 645 cell_1rw
* cell instance $18520 m0 *1 21.855,166.53
X$18520 127 637 128 644 645 cell_1rw
* cell instance $18521 r0 *1 21.855,163.8
X$18521 127 635 128 644 645 cell_1rw
* cell instance $18522 r0 *1 21.855,166.53
X$18522 127 636 128 644 645 cell_1rw
* cell instance $18523 m0 *1 21.855,169.26
X$18523 127 639 128 644 645 cell_1rw
* cell instance $18524 r0 *1 21.855,169.26
X$18524 127 638 128 644 645 cell_1rw
* cell instance $18525 m0 *1 21.855,171.99
X$18525 127 640 128 644 645 cell_1rw
* cell instance $18526 r0 *1 21.855,171.99
X$18526 127 641 128 644 645 cell_1rw
* cell instance $18527 m0 *1 21.855,174.72
X$18527 127 642 128 644 645 cell_1rw
* cell instance $18528 r0 *1 21.855,174.72
X$18528 127 643 128 644 645 cell_1rw
* cell instance $18529 r0 *1 22.56,87.36
X$18529 129 322 130 644 645 cell_1rw
* cell instance $18530 m0 *1 22.56,90.09
X$18530 129 581 130 644 645 cell_1rw
* cell instance $18531 m0 *1 22.56,92.82
X$18531 129 583 130 644 645 cell_1rw
* cell instance $18532 r0 *1 22.56,90.09
X$18532 129 580 130 644 645 cell_1rw
* cell instance $18533 r0 *1 22.56,92.82
X$18533 129 582 130 644 645 cell_1rw
* cell instance $18534 m0 *1 22.56,95.55
X$18534 129 584 130 644 645 cell_1rw
* cell instance $18535 r0 *1 22.56,95.55
X$18535 129 585 130 644 645 cell_1rw
* cell instance $18536 m0 *1 22.56,98.28
X$18536 129 586 130 644 645 cell_1rw
* cell instance $18537 r0 *1 22.56,98.28
X$18537 129 587 130 644 645 cell_1rw
* cell instance $18538 m0 *1 22.56,101.01
X$18538 129 588 130 644 645 cell_1rw
* cell instance $18539 m0 *1 22.56,103.74
X$18539 129 590 130 644 645 cell_1rw
* cell instance $18540 r0 *1 22.56,101.01
X$18540 129 589 130 644 645 cell_1rw
* cell instance $18541 r0 *1 22.56,103.74
X$18541 129 591 130 644 645 cell_1rw
* cell instance $18542 m0 *1 22.56,106.47
X$18542 129 593 130 644 645 cell_1rw
* cell instance $18543 r0 *1 22.56,106.47
X$18543 129 592 130 644 645 cell_1rw
* cell instance $18544 m0 *1 22.56,109.2
X$18544 129 594 130 644 645 cell_1rw
* cell instance $18545 r0 *1 22.56,109.2
X$18545 129 595 130 644 645 cell_1rw
* cell instance $18546 m0 *1 22.56,111.93
X$18546 129 597 130 644 645 cell_1rw
* cell instance $18547 r0 *1 22.56,111.93
X$18547 129 596 130 644 645 cell_1rw
* cell instance $18548 m0 *1 22.56,114.66
X$18548 129 598 130 644 645 cell_1rw
* cell instance $18549 r0 *1 22.56,114.66
X$18549 129 599 130 644 645 cell_1rw
* cell instance $18550 m0 *1 22.56,117.39
X$18550 129 600 130 644 645 cell_1rw
* cell instance $18551 m0 *1 22.56,120.12
X$18551 129 602 130 644 645 cell_1rw
* cell instance $18552 r0 *1 22.56,117.39
X$18552 129 601 130 644 645 cell_1rw
* cell instance $18553 r0 *1 22.56,120.12
X$18553 129 603 130 644 645 cell_1rw
* cell instance $18554 m0 *1 22.56,122.85
X$18554 129 604 130 644 645 cell_1rw
* cell instance $18555 r0 *1 22.56,122.85
X$18555 129 605 130 644 645 cell_1rw
* cell instance $18556 m0 *1 22.56,125.58
X$18556 129 606 130 644 645 cell_1rw
* cell instance $18557 m0 *1 22.56,128.31
X$18557 129 609 130 644 645 cell_1rw
* cell instance $18558 r0 *1 22.56,125.58
X$18558 129 607 130 644 645 cell_1rw
* cell instance $18559 m0 *1 22.56,131.04
X$18559 129 610 130 644 645 cell_1rw
* cell instance $18560 r0 *1 22.56,128.31
X$18560 129 608 130 644 645 cell_1rw
* cell instance $18561 r0 *1 22.56,131.04
X$18561 129 611 130 644 645 cell_1rw
* cell instance $18562 m0 *1 22.56,133.77
X$18562 129 612 130 644 645 cell_1rw
* cell instance $18563 r0 *1 22.56,133.77
X$18563 129 613 130 644 645 cell_1rw
* cell instance $18564 m0 *1 22.56,136.5
X$18564 129 615 130 644 645 cell_1rw
* cell instance $18565 r0 *1 22.56,136.5
X$18565 129 614 130 644 645 cell_1rw
* cell instance $18566 m0 *1 22.56,139.23
X$18566 129 617 130 644 645 cell_1rw
* cell instance $18567 r0 *1 22.56,139.23
X$18567 129 616 130 644 645 cell_1rw
* cell instance $18568 m0 *1 22.56,141.96
X$18568 129 618 130 644 645 cell_1rw
* cell instance $18569 r0 *1 22.56,141.96
X$18569 129 619 130 644 645 cell_1rw
* cell instance $18570 m0 *1 22.56,144.69
X$18570 129 620 130 644 645 cell_1rw
* cell instance $18571 r0 *1 22.56,144.69
X$18571 129 621 130 644 645 cell_1rw
* cell instance $18572 m0 *1 22.56,147.42
X$18572 129 622 130 644 645 cell_1rw
* cell instance $18573 r0 *1 22.56,147.42
X$18573 129 623 130 644 645 cell_1rw
* cell instance $18574 m0 *1 22.56,150.15
X$18574 129 624 130 644 645 cell_1rw
* cell instance $18575 r0 *1 22.56,150.15
X$18575 129 625 130 644 645 cell_1rw
* cell instance $18576 m0 *1 22.56,152.88
X$18576 129 626 130 644 645 cell_1rw
* cell instance $18577 r0 *1 22.56,152.88
X$18577 129 627 130 644 645 cell_1rw
* cell instance $18578 m0 *1 22.56,155.61
X$18578 129 628 130 644 645 cell_1rw
* cell instance $18579 m0 *1 22.56,158.34
X$18579 129 630 130 644 645 cell_1rw
* cell instance $18580 r0 *1 22.56,155.61
X$18580 129 629 130 644 645 cell_1rw
* cell instance $18581 r0 *1 22.56,158.34
X$18581 129 631 130 644 645 cell_1rw
* cell instance $18582 m0 *1 22.56,161.07
X$18582 129 632 130 644 645 cell_1rw
* cell instance $18583 r0 *1 22.56,161.07
X$18583 129 633 130 644 645 cell_1rw
* cell instance $18584 m0 *1 22.56,163.8
X$18584 129 634 130 644 645 cell_1rw
* cell instance $18585 r0 *1 22.56,163.8
X$18585 129 635 130 644 645 cell_1rw
* cell instance $18586 m0 *1 22.56,166.53
X$18586 129 637 130 644 645 cell_1rw
* cell instance $18587 r0 *1 22.56,166.53
X$18587 129 636 130 644 645 cell_1rw
* cell instance $18588 m0 *1 22.56,169.26
X$18588 129 639 130 644 645 cell_1rw
* cell instance $18589 r0 *1 22.56,169.26
X$18589 129 638 130 644 645 cell_1rw
* cell instance $18590 m0 *1 22.56,171.99
X$18590 129 640 130 644 645 cell_1rw
* cell instance $18591 m0 *1 22.56,174.72
X$18591 129 642 130 644 645 cell_1rw
* cell instance $18592 r0 *1 22.56,171.99
X$18592 129 641 130 644 645 cell_1rw
* cell instance $18593 r0 *1 22.56,174.72
X$18593 129 643 130 644 645 cell_1rw
* cell instance $18594 m0 *1 23.265,90.09
X$18594 131 581 132 644 645 cell_1rw
* cell instance $18595 r0 *1 23.265,87.36
X$18595 131 322 132 644 645 cell_1rw
* cell instance $18596 r0 *1 23.265,90.09
X$18596 131 580 132 644 645 cell_1rw
* cell instance $18597 m0 *1 23.265,92.82
X$18597 131 583 132 644 645 cell_1rw
* cell instance $18598 r0 *1 23.265,92.82
X$18598 131 582 132 644 645 cell_1rw
* cell instance $18599 m0 *1 23.265,95.55
X$18599 131 584 132 644 645 cell_1rw
* cell instance $18600 m0 *1 23.265,98.28
X$18600 131 586 132 644 645 cell_1rw
* cell instance $18601 r0 *1 23.265,95.55
X$18601 131 585 132 644 645 cell_1rw
* cell instance $18602 r0 *1 23.265,98.28
X$18602 131 587 132 644 645 cell_1rw
* cell instance $18603 m0 *1 23.265,101.01
X$18603 131 588 132 644 645 cell_1rw
* cell instance $18604 r0 *1 23.265,101.01
X$18604 131 589 132 644 645 cell_1rw
* cell instance $18605 m0 *1 23.265,103.74
X$18605 131 590 132 644 645 cell_1rw
* cell instance $18606 r0 *1 23.265,103.74
X$18606 131 591 132 644 645 cell_1rw
* cell instance $18607 m0 *1 23.265,106.47
X$18607 131 593 132 644 645 cell_1rw
* cell instance $18608 r0 *1 23.265,106.47
X$18608 131 592 132 644 645 cell_1rw
* cell instance $18609 m0 *1 23.265,109.2
X$18609 131 594 132 644 645 cell_1rw
* cell instance $18610 m0 *1 23.265,111.93
X$18610 131 597 132 644 645 cell_1rw
* cell instance $18611 r0 *1 23.265,109.2
X$18611 131 595 132 644 645 cell_1rw
* cell instance $18612 r0 *1 23.265,111.93
X$18612 131 596 132 644 645 cell_1rw
* cell instance $18613 m0 *1 23.265,114.66
X$18613 131 598 132 644 645 cell_1rw
* cell instance $18614 m0 *1 23.265,117.39
X$18614 131 600 132 644 645 cell_1rw
* cell instance $18615 r0 *1 23.265,114.66
X$18615 131 599 132 644 645 cell_1rw
* cell instance $18616 r0 *1 23.265,117.39
X$18616 131 601 132 644 645 cell_1rw
* cell instance $18617 m0 *1 23.265,120.12
X$18617 131 602 132 644 645 cell_1rw
* cell instance $18618 r0 *1 23.265,120.12
X$18618 131 603 132 644 645 cell_1rw
* cell instance $18619 m0 *1 23.265,122.85
X$18619 131 604 132 644 645 cell_1rw
* cell instance $18620 r0 *1 23.265,122.85
X$18620 131 605 132 644 645 cell_1rw
* cell instance $18621 m0 *1 23.265,125.58
X$18621 131 606 132 644 645 cell_1rw
* cell instance $18622 r0 *1 23.265,125.58
X$18622 131 607 132 644 645 cell_1rw
* cell instance $18623 m0 *1 23.265,128.31
X$18623 131 609 132 644 645 cell_1rw
* cell instance $18624 r0 *1 23.265,128.31
X$18624 131 608 132 644 645 cell_1rw
* cell instance $18625 m0 *1 23.265,131.04
X$18625 131 610 132 644 645 cell_1rw
* cell instance $18626 r0 *1 23.265,131.04
X$18626 131 611 132 644 645 cell_1rw
* cell instance $18627 m0 *1 23.265,133.77
X$18627 131 612 132 644 645 cell_1rw
* cell instance $18628 m0 *1 23.265,136.5
X$18628 131 615 132 644 645 cell_1rw
* cell instance $18629 r0 *1 23.265,133.77
X$18629 131 613 132 644 645 cell_1rw
* cell instance $18630 r0 *1 23.265,136.5
X$18630 131 614 132 644 645 cell_1rw
* cell instance $18631 m0 *1 23.265,139.23
X$18631 131 617 132 644 645 cell_1rw
* cell instance $18632 r0 *1 23.265,139.23
X$18632 131 616 132 644 645 cell_1rw
* cell instance $18633 m0 *1 23.265,141.96
X$18633 131 618 132 644 645 cell_1rw
* cell instance $18634 m0 *1 23.265,144.69
X$18634 131 620 132 644 645 cell_1rw
* cell instance $18635 r0 *1 23.265,141.96
X$18635 131 619 132 644 645 cell_1rw
* cell instance $18636 m0 *1 23.265,147.42
X$18636 131 622 132 644 645 cell_1rw
* cell instance $18637 r0 *1 23.265,144.69
X$18637 131 621 132 644 645 cell_1rw
* cell instance $18638 r0 *1 23.265,147.42
X$18638 131 623 132 644 645 cell_1rw
* cell instance $18639 m0 *1 23.265,150.15
X$18639 131 624 132 644 645 cell_1rw
* cell instance $18640 r0 *1 23.265,150.15
X$18640 131 625 132 644 645 cell_1rw
* cell instance $18641 m0 *1 23.265,152.88
X$18641 131 626 132 644 645 cell_1rw
* cell instance $18642 r0 *1 23.265,152.88
X$18642 131 627 132 644 645 cell_1rw
* cell instance $18643 m0 *1 23.265,155.61
X$18643 131 628 132 644 645 cell_1rw
* cell instance $18644 r0 *1 23.265,155.61
X$18644 131 629 132 644 645 cell_1rw
* cell instance $18645 m0 *1 23.265,158.34
X$18645 131 630 132 644 645 cell_1rw
* cell instance $18646 r0 *1 23.265,158.34
X$18646 131 631 132 644 645 cell_1rw
* cell instance $18647 m0 *1 23.265,161.07
X$18647 131 632 132 644 645 cell_1rw
* cell instance $18648 r0 *1 23.265,161.07
X$18648 131 633 132 644 645 cell_1rw
* cell instance $18649 m0 *1 23.265,163.8
X$18649 131 634 132 644 645 cell_1rw
* cell instance $18650 r0 *1 23.265,163.8
X$18650 131 635 132 644 645 cell_1rw
* cell instance $18651 m0 *1 23.265,166.53
X$18651 131 637 132 644 645 cell_1rw
* cell instance $18652 r0 *1 23.265,166.53
X$18652 131 636 132 644 645 cell_1rw
* cell instance $18653 m0 *1 23.265,169.26
X$18653 131 639 132 644 645 cell_1rw
* cell instance $18654 r0 *1 23.265,169.26
X$18654 131 638 132 644 645 cell_1rw
* cell instance $18655 m0 *1 23.265,171.99
X$18655 131 640 132 644 645 cell_1rw
* cell instance $18656 r0 *1 23.265,171.99
X$18656 131 641 132 644 645 cell_1rw
* cell instance $18657 m0 *1 23.265,174.72
X$18657 131 642 132 644 645 cell_1rw
* cell instance $18658 r0 *1 23.265,174.72
X$18658 131 643 132 644 645 cell_1rw
* cell instance $18659 m0 *1 23.97,90.09
X$18659 133 581 134 644 645 cell_1rw
* cell instance $18660 r0 *1 23.97,87.36
X$18660 133 322 134 644 645 cell_1rw
* cell instance $18661 r0 *1 23.97,90.09
X$18661 133 580 134 644 645 cell_1rw
* cell instance $18662 m0 *1 23.97,92.82
X$18662 133 583 134 644 645 cell_1rw
* cell instance $18663 r0 *1 23.97,92.82
X$18663 133 582 134 644 645 cell_1rw
* cell instance $18664 m0 *1 23.97,95.55
X$18664 133 584 134 644 645 cell_1rw
* cell instance $18665 r0 *1 23.97,95.55
X$18665 133 585 134 644 645 cell_1rw
* cell instance $18666 m0 *1 23.97,98.28
X$18666 133 586 134 644 645 cell_1rw
* cell instance $18667 r0 *1 23.97,98.28
X$18667 133 587 134 644 645 cell_1rw
* cell instance $18668 m0 *1 23.97,101.01
X$18668 133 588 134 644 645 cell_1rw
* cell instance $18669 m0 *1 23.97,103.74
X$18669 133 590 134 644 645 cell_1rw
* cell instance $18670 r0 *1 23.97,101.01
X$18670 133 589 134 644 645 cell_1rw
* cell instance $18671 r0 *1 23.97,103.74
X$18671 133 591 134 644 645 cell_1rw
* cell instance $18672 m0 *1 23.97,106.47
X$18672 133 593 134 644 645 cell_1rw
* cell instance $18673 m0 *1 23.97,109.2
X$18673 133 594 134 644 645 cell_1rw
* cell instance $18674 r0 *1 23.97,106.47
X$18674 133 592 134 644 645 cell_1rw
* cell instance $18675 r0 *1 23.97,109.2
X$18675 133 595 134 644 645 cell_1rw
* cell instance $18676 m0 *1 23.97,111.93
X$18676 133 597 134 644 645 cell_1rw
* cell instance $18677 r0 *1 23.97,111.93
X$18677 133 596 134 644 645 cell_1rw
* cell instance $18678 m0 *1 23.97,114.66
X$18678 133 598 134 644 645 cell_1rw
* cell instance $18679 r0 *1 23.97,114.66
X$18679 133 599 134 644 645 cell_1rw
* cell instance $18680 m0 *1 23.97,117.39
X$18680 133 600 134 644 645 cell_1rw
* cell instance $18681 r0 *1 23.97,117.39
X$18681 133 601 134 644 645 cell_1rw
* cell instance $18682 m0 *1 23.97,120.12
X$18682 133 602 134 644 645 cell_1rw
* cell instance $18683 m0 *1 23.97,122.85
X$18683 133 604 134 644 645 cell_1rw
* cell instance $18684 r0 *1 23.97,120.12
X$18684 133 603 134 644 645 cell_1rw
* cell instance $18685 m0 *1 23.97,125.58
X$18685 133 606 134 644 645 cell_1rw
* cell instance $18686 r0 *1 23.97,122.85
X$18686 133 605 134 644 645 cell_1rw
* cell instance $18687 r0 *1 23.97,125.58
X$18687 133 607 134 644 645 cell_1rw
* cell instance $18688 m0 *1 23.97,128.31
X$18688 133 609 134 644 645 cell_1rw
* cell instance $18689 r0 *1 23.97,128.31
X$18689 133 608 134 644 645 cell_1rw
* cell instance $18690 m0 *1 23.97,131.04
X$18690 133 610 134 644 645 cell_1rw
* cell instance $18691 r0 *1 23.97,131.04
X$18691 133 611 134 644 645 cell_1rw
* cell instance $18692 m0 *1 23.97,133.77
X$18692 133 612 134 644 645 cell_1rw
* cell instance $18693 r0 *1 23.97,133.77
X$18693 133 613 134 644 645 cell_1rw
* cell instance $18694 m0 *1 23.97,136.5
X$18694 133 615 134 644 645 cell_1rw
* cell instance $18695 r0 *1 23.97,136.5
X$18695 133 614 134 644 645 cell_1rw
* cell instance $18696 m0 *1 23.97,139.23
X$18696 133 617 134 644 645 cell_1rw
* cell instance $18697 r0 *1 23.97,139.23
X$18697 133 616 134 644 645 cell_1rw
* cell instance $18698 m0 *1 23.97,141.96
X$18698 133 618 134 644 645 cell_1rw
* cell instance $18699 r0 *1 23.97,141.96
X$18699 133 619 134 644 645 cell_1rw
* cell instance $18700 m0 *1 23.97,144.69
X$18700 133 620 134 644 645 cell_1rw
* cell instance $18701 r0 *1 23.97,144.69
X$18701 133 621 134 644 645 cell_1rw
* cell instance $18702 m0 *1 23.97,147.42
X$18702 133 622 134 644 645 cell_1rw
* cell instance $18703 m0 *1 23.97,150.15
X$18703 133 624 134 644 645 cell_1rw
* cell instance $18704 r0 *1 23.97,147.42
X$18704 133 623 134 644 645 cell_1rw
* cell instance $18705 r0 *1 23.97,150.15
X$18705 133 625 134 644 645 cell_1rw
* cell instance $18706 m0 *1 23.97,152.88
X$18706 133 626 134 644 645 cell_1rw
* cell instance $18707 r0 *1 23.97,152.88
X$18707 133 627 134 644 645 cell_1rw
* cell instance $18708 m0 *1 23.97,155.61
X$18708 133 628 134 644 645 cell_1rw
* cell instance $18709 r0 *1 23.97,155.61
X$18709 133 629 134 644 645 cell_1rw
* cell instance $18710 m0 *1 23.97,158.34
X$18710 133 630 134 644 645 cell_1rw
* cell instance $18711 m0 *1 23.97,161.07
X$18711 133 632 134 644 645 cell_1rw
* cell instance $18712 r0 *1 23.97,158.34
X$18712 133 631 134 644 645 cell_1rw
* cell instance $18713 r0 *1 23.97,161.07
X$18713 133 633 134 644 645 cell_1rw
* cell instance $18714 m0 *1 23.97,163.8
X$18714 133 634 134 644 645 cell_1rw
* cell instance $18715 r0 *1 23.97,163.8
X$18715 133 635 134 644 645 cell_1rw
* cell instance $18716 m0 *1 23.97,166.53
X$18716 133 637 134 644 645 cell_1rw
* cell instance $18717 r0 *1 23.97,166.53
X$18717 133 636 134 644 645 cell_1rw
* cell instance $18718 m0 *1 23.97,169.26
X$18718 133 639 134 644 645 cell_1rw
* cell instance $18719 r0 *1 23.97,169.26
X$18719 133 638 134 644 645 cell_1rw
* cell instance $18720 m0 *1 23.97,171.99
X$18720 133 640 134 644 645 cell_1rw
* cell instance $18721 r0 *1 23.97,171.99
X$18721 133 641 134 644 645 cell_1rw
* cell instance $18722 m0 *1 23.97,174.72
X$18722 133 642 134 644 645 cell_1rw
* cell instance $18723 r0 *1 23.97,174.72
X$18723 133 643 134 644 645 cell_1rw
* cell instance $18724 r0 *1 24.675,87.36
X$18724 135 322 136 644 645 cell_1rw
* cell instance $18725 m0 *1 24.675,90.09
X$18725 135 581 136 644 645 cell_1rw
* cell instance $18726 r0 *1 24.675,90.09
X$18726 135 580 136 644 645 cell_1rw
* cell instance $18727 m0 *1 24.675,92.82
X$18727 135 583 136 644 645 cell_1rw
* cell instance $18728 r0 *1 24.675,92.82
X$18728 135 582 136 644 645 cell_1rw
* cell instance $18729 m0 *1 24.675,95.55
X$18729 135 584 136 644 645 cell_1rw
* cell instance $18730 r0 *1 24.675,95.55
X$18730 135 585 136 644 645 cell_1rw
* cell instance $18731 m0 *1 24.675,98.28
X$18731 135 586 136 644 645 cell_1rw
* cell instance $18732 m0 *1 24.675,101.01
X$18732 135 588 136 644 645 cell_1rw
* cell instance $18733 r0 *1 24.675,98.28
X$18733 135 587 136 644 645 cell_1rw
* cell instance $18734 r0 *1 24.675,101.01
X$18734 135 589 136 644 645 cell_1rw
* cell instance $18735 m0 *1 24.675,103.74
X$18735 135 590 136 644 645 cell_1rw
* cell instance $18736 r0 *1 24.675,103.74
X$18736 135 591 136 644 645 cell_1rw
* cell instance $18737 m0 *1 24.675,106.47
X$18737 135 593 136 644 645 cell_1rw
* cell instance $18738 r0 *1 24.675,106.47
X$18738 135 592 136 644 645 cell_1rw
* cell instance $18739 m0 *1 24.675,109.2
X$18739 135 594 136 644 645 cell_1rw
* cell instance $18740 r0 *1 24.675,109.2
X$18740 135 595 136 644 645 cell_1rw
* cell instance $18741 m0 *1 24.675,111.93
X$18741 135 597 136 644 645 cell_1rw
* cell instance $18742 r0 *1 24.675,111.93
X$18742 135 596 136 644 645 cell_1rw
* cell instance $18743 m0 *1 24.675,114.66
X$18743 135 598 136 644 645 cell_1rw
* cell instance $18744 r0 *1 24.675,114.66
X$18744 135 599 136 644 645 cell_1rw
* cell instance $18745 m0 *1 24.675,117.39
X$18745 135 600 136 644 645 cell_1rw
* cell instance $18746 r0 *1 24.675,117.39
X$18746 135 601 136 644 645 cell_1rw
* cell instance $18747 m0 *1 24.675,120.12
X$18747 135 602 136 644 645 cell_1rw
* cell instance $18748 m0 *1 24.675,122.85
X$18748 135 604 136 644 645 cell_1rw
* cell instance $18749 r0 *1 24.675,120.12
X$18749 135 603 136 644 645 cell_1rw
* cell instance $18750 r0 *1 24.675,122.85
X$18750 135 605 136 644 645 cell_1rw
* cell instance $18751 m0 *1 24.675,125.58
X$18751 135 606 136 644 645 cell_1rw
* cell instance $18752 r0 *1 24.675,125.58
X$18752 135 607 136 644 645 cell_1rw
* cell instance $18753 m0 *1 24.675,128.31
X$18753 135 609 136 644 645 cell_1rw
* cell instance $18754 r0 *1 24.675,128.31
X$18754 135 608 136 644 645 cell_1rw
* cell instance $18755 m0 *1 24.675,131.04
X$18755 135 610 136 644 645 cell_1rw
* cell instance $18756 r0 *1 24.675,131.04
X$18756 135 611 136 644 645 cell_1rw
* cell instance $18757 m0 *1 24.675,133.77
X$18757 135 612 136 644 645 cell_1rw
* cell instance $18758 r0 *1 24.675,133.77
X$18758 135 613 136 644 645 cell_1rw
* cell instance $18759 m0 *1 24.675,136.5
X$18759 135 615 136 644 645 cell_1rw
* cell instance $18760 r0 *1 24.675,136.5
X$18760 135 614 136 644 645 cell_1rw
* cell instance $18761 m0 *1 24.675,139.23
X$18761 135 617 136 644 645 cell_1rw
* cell instance $18762 r0 *1 24.675,139.23
X$18762 135 616 136 644 645 cell_1rw
* cell instance $18763 m0 *1 24.675,141.96
X$18763 135 618 136 644 645 cell_1rw
* cell instance $18764 m0 *1 24.675,144.69
X$18764 135 620 136 644 645 cell_1rw
* cell instance $18765 r0 *1 24.675,141.96
X$18765 135 619 136 644 645 cell_1rw
* cell instance $18766 m0 *1 24.675,147.42
X$18766 135 622 136 644 645 cell_1rw
* cell instance $18767 r0 *1 24.675,144.69
X$18767 135 621 136 644 645 cell_1rw
* cell instance $18768 m0 *1 24.675,150.15
X$18768 135 624 136 644 645 cell_1rw
* cell instance $18769 r0 *1 24.675,147.42
X$18769 135 623 136 644 645 cell_1rw
* cell instance $18770 r0 *1 24.675,150.15
X$18770 135 625 136 644 645 cell_1rw
* cell instance $18771 m0 *1 24.675,152.88
X$18771 135 626 136 644 645 cell_1rw
* cell instance $18772 r0 *1 24.675,152.88
X$18772 135 627 136 644 645 cell_1rw
* cell instance $18773 m0 *1 24.675,155.61
X$18773 135 628 136 644 645 cell_1rw
* cell instance $18774 r0 *1 24.675,155.61
X$18774 135 629 136 644 645 cell_1rw
* cell instance $18775 m0 *1 24.675,158.34
X$18775 135 630 136 644 645 cell_1rw
* cell instance $18776 r0 *1 24.675,158.34
X$18776 135 631 136 644 645 cell_1rw
* cell instance $18777 m0 *1 24.675,161.07
X$18777 135 632 136 644 645 cell_1rw
* cell instance $18778 r0 *1 24.675,161.07
X$18778 135 633 136 644 645 cell_1rw
* cell instance $18779 m0 *1 24.675,163.8
X$18779 135 634 136 644 645 cell_1rw
* cell instance $18780 r0 *1 24.675,163.8
X$18780 135 635 136 644 645 cell_1rw
* cell instance $18781 m0 *1 24.675,166.53
X$18781 135 637 136 644 645 cell_1rw
* cell instance $18782 m0 *1 24.675,169.26
X$18782 135 639 136 644 645 cell_1rw
* cell instance $18783 r0 *1 24.675,166.53
X$18783 135 636 136 644 645 cell_1rw
* cell instance $18784 m0 *1 24.675,171.99
X$18784 135 640 136 644 645 cell_1rw
* cell instance $18785 r0 *1 24.675,169.26
X$18785 135 638 136 644 645 cell_1rw
* cell instance $18786 r0 *1 24.675,171.99
X$18786 135 641 136 644 645 cell_1rw
* cell instance $18787 m0 *1 24.675,174.72
X$18787 135 642 136 644 645 cell_1rw
* cell instance $18788 r0 *1 24.675,174.72
X$18788 135 643 136 644 645 cell_1rw
* cell instance $18789 r0 *1 25.38,87.36
X$18789 137 322 138 644 645 cell_1rw
* cell instance $18790 m0 *1 25.38,90.09
X$18790 137 581 138 644 645 cell_1rw
* cell instance $18791 r0 *1 25.38,90.09
X$18791 137 580 138 644 645 cell_1rw
* cell instance $18792 m0 *1 25.38,92.82
X$18792 137 583 138 644 645 cell_1rw
* cell instance $18793 r0 *1 25.38,92.82
X$18793 137 582 138 644 645 cell_1rw
* cell instance $18794 m0 *1 25.38,95.55
X$18794 137 584 138 644 645 cell_1rw
* cell instance $18795 r0 *1 25.38,95.55
X$18795 137 585 138 644 645 cell_1rw
* cell instance $18796 m0 *1 25.38,98.28
X$18796 137 586 138 644 645 cell_1rw
* cell instance $18797 r0 *1 25.38,98.28
X$18797 137 587 138 644 645 cell_1rw
* cell instance $18798 m0 *1 25.38,101.01
X$18798 137 588 138 644 645 cell_1rw
* cell instance $18799 r0 *1 25.38,101.01
X$18799 137 589 138 644 645 cell_1rw
* cell instance $18800 m0 *1 25.38,103.74
X$18800 137 590 138 644 645 cell_1rw
* cell instance $18801 r0 *1 25.38,103.74
X$18801 137 591 138 644 645 cell_1rw
* cell instance $18802 m0 *1 25.38,106.47
X$18802 137 593 138 644 645 cell_1rw
* cell instance $18803 r0 *1 25.38,106.47
X$18803 137 592 138 644 645 cell_1rw
* cell instance $18804 m0 *1 25.38,109.2
X$18804 137 594 138 644 645 cell_1rw
* cell instance $18805 r0 *1 25.38,109.2
X$18805 137 595 138 644 645 cell_1rw
* cell instance $18806 m0 *1 25.38,111.93
X$18806 137 597 138 644 645 cell_1rw
* cell instance $18807 r0 *1 25.38,111.93
X$18807 137 596 138 644 645 cell_1rw
* cell instance $18808 m0 *1 25.38,114.66
X$18808 137 598 138 644 645 cell_1rw
* cell instance $18809 r0 *1 25.38,114.66
X$18809 137 599 138 644 645 cell_1rw
* cell instance $18810 m0 *1 25.38,117.39
X$18810 137 600 138 644 645 cell_1rw
* cell instance $18811 r0 *1 25.38,117.39
X$18811 137 601 138 644 645 cell_1rw
* cell instance $18812 m0 *1 25.38,120.12
X$18812 137 602 138 644 645 cell_1rw
* cell instance $18813 r0 *1 25.38,120.12
X$18813 137 603 138 644 645 cell_1rw
* cell instance $18814 m0 *1 25.38,122.85
X$18814 137 604 138 644 645 cell_1rw
* cell instance $18815 r0 *1 25.38,122.85
X$18815 137 605 138 644 645 cell_1rw
* cell instance $18816 m0 *1 25.38,125.58
X$18816 137 606 138 644 645 cell_1rw
* cell instance $18817 r0 *1 25.38,125.58
X$18817 137 607 138 644 645 cell_1rw
* cell instance $18818 m0 *1 25.38,128.31
X$18818 137 609 138 644 645 cell_1rw
* cell instance $18819 r0 *1 25.38,128.31
X$18819 137 608 138 644 645 cell_1rw
* cell instance $18820 m0 *1 25.38,131.04
X$18820 137 610 138 644 645 cell_1rw
* cell instance $18821 r0 *1 25.38,131.04
X$18821 137 611 138 644 645 cell_1rw
* cell instance $18822 m0 *1 25.38,133.77
X$18822 137 612 138 644 645 cell_1rw
* cell instance $18823 r0 *1 25.38,133.77
X$18823 137 613 138 644 645 cell_1rw
* cell instance $18824 m0 *1 25.38,136.5
X$18824 137 615 138 644 645 cell_1rw
* cell instance $18825 r0 *1 25.38,136.5
X$18825 137 614 138 644 645 cell_1rw
* cell instance $18826 m0 *1 25.38,139.23
X$18826 137 617 138 644 645 cell_1rw
* cell instance $18827 r0 *1 25.38,139.23
X$18827 137 616 138 644 645 cell_1rw
* cell instance $18828 m0 *1 25.38,141.96
X$18828 137 618 138 644 645 cell_1rw
* cell instance $18829 r0 *1 25.38,141.96
X$18829 137 619 138 644 645 cell_1rw
* cell instance $18830 m0 *1 25.38,144.69
X$18830 137 620 138 644 645 cell_1rw
* cell instance $18831 r0 *1 25.38,144.69
X$18831 137 621 138 644 645 cell_1rw
* cell instance $18832 m0 *1 25.38,147.42
X$18832 137 622 138 644 645 cell_1rw
* cell instance $18833 r0 *1 25.38,147.42
X$18833 137 623 138 644 645 cell_1rw
* cell instance $18834 m0 *1 25.38,150.15
X$18834 137 624 138 644 645 cell_1rw
* cell instance $18835 r0 *1 25.38,150.15
X$18835 137 625 138 644 645 cell_1rw
* cell instance $18836 m0 *1 25.38,152.88
X$18836 137 626 138 644 645 cell_1rw
* cell instance $18837 r0 *1 25.38,152.88
X$18837 137 627 138 644 645 cell_1rw
* cell instance $18838 m0 *1 25.38,155.61
X$18838 137 628 138 644 645 cell_1rw
* cell instance $18839 r0 *1 25.38,155.61
X$18839 137 629 138 644 645 cell_1rw
* cell instance $18840 m0 *1 25.38,158.34
X$18840 137 630 138 644 645 cell_1rw
* cell instance $18841 r0 *1 25.38,158.34
X$18841 137 631 138 644 645 cell_1rw
* cell instance $18842 m0 *1 25.38,161.07
X$18842 137 632 138 644 645 cell_1rw
* cell instance $18843 r0 *1 25.38,161.07
X$18843 137 633 138 644 645 cell_1rw
* cell instance $18844 m0 *1 25.38,163.8
X$18844 137 634 138 644 645 cell_1rw
* cell instance $18845 r0 *1 25.38,163.8
X$18845 137 635 138 644 645 cell_1rw
* cell instance $18846 m0 *1 25.38,166.53
X$18846 137 637 138 644 645 cell_1rw
* cell instance $18847 r0 *1 25.38,166.53
X$18847 137 636 138 644 645 cell_1rw
* cell instance $18848 m0 *1 25.38,169.26
X$18848 137 639 138 644 645 cell_1rw
* cell instance $18849 m0 *1 25.38,171.99
X$18849 137 640 138 644 645 cell_1rw
* cell instance $18850 r0 *1 25.38,169.26
X$18850 137 638 138 644 645 cell_1rw
* cell instance $18851 r0 *1 25.38,171.99
X$18851 137 641 138 644 645 cell_1rw
* cell instance $18852 m0 *1 25.38,174.72
X$18852 137 642 138 644 645 cell_1rw
* cell instance $18853 r0 *1 25.38,174.72
X$18853 137 643 138 644 645 cell_1rw
* cell instance $18854 r0 *1 26.085,87.36
X$18854 139 322 140 644 645 cell_1rw
* cell instance $18855 m0 *1 26.085,90.09
X$18855 139 581 140 644 645 cell_1rw
* cell instance $18856 r0 *1 26.085,90.09
X$18856 139 580 140 644 645 cell_1rw
* cell instance $18857 m0 *1 26.085,92.82
X$18857 139 583 140 644 645 cell_1rw
* cell instance $18858 r0 *1 26.085,92.82
X$18858 139 582 140 644 645 cell_1rw
* cell instance $18859 m0 *1 26.085,95.55
X$18859 139 584 140 644 645 cell_1rw
* cell instance $18860 m0 *1 26.085,98.28
X$18860 139 586 140 644 645 cell_1rw
* cell instance $18861 r0 *1 26.085,95.55
X$18861 139 585 140 644 645 cell_1rw
* cell instance $18862 m0 *1 26.085,101.01
X$18862 139 588 140 644 645 cell_1rw
* cell instance $18863 r0 *1 26.085,98.28
X$18863 139 587 140 644 645 cell_1rw
* cell instance $18864 r0 *1 26.085,101.01
X$18864 139 589 140 644 645 cell_1rw
* cell instance $18865 m0 *1 26.085,103.74
X$18865 139 590 140 644 645 cell_1rw
* cell instance $18866 r0 *1 26.085,103.74
X$18866 139 591 140 644 645 cell_1rw
* cell instance $18867 m0 *1 26.085,106.47
X$18867 139 593 140 644 645 cell_1rw
* cell instance $18868 r0 *1 26.085,106.47
X$18868 139 592 140 644 645 cell_1rw
* cell instance $18869 m0 *1 26.085,109.2
X$18869 139 594 140 644 645 cell_1rw
* cell instance $18870 r0 *1 26.085,109.2
X$18870 139 595 140 644 645 cell_1rw
* cell instance $18871 m0 *1 26.085,111.93
X$18871 139 597 140 644 645 cell_1rw
* cell instance $18872 r0 *1 26.085,111.93
X$18872 139 596 140 644 645 cell_1rw
* cell instance $18873 m0 *1 26.085,114.66
X$18873 139 598 140 644 645 cell_1rw
* cell instance $18874 r0 *1 26.085,114.66
X$18874 139 599 140 644 645 cell_1rw
* cell instance $18875 m0 *1 26.085,117.39
X$18875 139 600 140 644 645 cell_1rw
* cell instance $18876 r0 *1 26.085,117.39
X$18876 139 601 140 644 645 cell_1rw
* cell instance $18877 m0 *1 26.085,120.12
X$18877 139 602 140 644 645 cell_1rw
* cell instance $18878 r0 *1 26.085,120.12
X$18878 139 603 140 644 645 cell_1rw
* cell instance $18879 m0 *1 26.085,122.85
X$18879 139 604 140 644 645 cell_1rw
* cell instance $18880 r0 *1 26.085,122.85
X$18880 139 605 140 644 645 cell_1rw
* cell instance $18881 m0 *1 26.085,125.58
X$18881 139 606 140 644 645 cell_1rw
* cell instance $18882 r0 *1 26.085,125.58
X$18882 139 607 140 644 645 cell_1rw
* cell instance $18883 m0 *1 26.085,128.31
X$18883 139 609 140 644 645 cell_1rw
* cell instance $18884 r0 *1 26.085,128.31
X$18884 139 608 140 644 645 cell_1rw
* cell instance $18885 m0 *1 26.085,131.04
X$18885 139 610 140 644 645 cell_1rw
* cell instance $18886 r0 *1 26.085,131.04
X$18886 139 611 140 644 645 cell_1rw
* cell instance $18887 m0 *1 26.085,133.77
X$18887 139 612 140 644 645 cell_1rw
* cell instance $18888 m0 *1 26.085,136.5
X$18888 139 615 140 644 645 cell_1rw
* cell instance $18889 r0 *1 26.085,133.77
X$18889 139 613 140 644 645 cell_1rw
* cell instance $18890 r0 *1 26.085,136.5
X$18890 139 614 140 644 645 cell_1rw
* cell instance $18891 m0 *1 26.085,139.23
X$18891 139 617 140 644 645 cell_1rw
* cell instance $18892 r0 *1 26.085,139.23
X$18892 139 616 140 644 645 cell_1rw
* cell instance $18893 m0 *1 26.085,141.96
X$18893 139 618 140 644 645 cell_1rw
* cell instance $18894 r0 *1 26.085,141.96
X$18894 139 619 140 644 645 cell_1rw
* cell instance $18895 m0 *1 26.085,144.69
X$18895 139 620 140 644 645 cell_1rw
* cell instance $18896 r0 *1 26.085,144.69
X$18896 139 621 140 644 645 cell_1rw
* cell instance $18897 m0 *1 26.085,147.42
X$18897 139 622 140 644 645 cell_1rw
* cell instance $18898 r0 *1 26.085,147.42
X$18898 139 623 140 644 645 cell_1rw
* cell instance $18899 m0 *1 26.085,150.15
X$18899 139 624 140 644 645 cell_1rw
* cell instance $18900 r0 *1 26.085,150.15
X$18900 139 625 140 644 645 cell_1rw
* cell instance $18901 m0 *1 26.085,152.88
X$18901 139 626 140 644 645 cell_1rw
* cell instance $18902 r0 *1 26.085,152.88
X$18902 139 627 140 644 645 cell_1rw
* cell instance $18903 m0 *1 26.085,155.61
X$18903 139 628 140 644 645 cell_1rw
* cell instance $18904 m0 *1 26.085,158.34
X$18904 139 630 140 644 645 cell_1rw
* cell instance $18905 r0 *1 26.085,155.61
X$18905 139 629 140 644 645 cell_1rw
* cell instance $18906 r0 *1 26.085,158.34
X$18906 139 631 140 644 645 cell_1rw
* cell instance $18907 m0 *1 26.085,161.07
X$18907 139 632 140 644 645 cell_1rw
* cell instance $18908 r0 *1 26.085,161.07
X$18908 139 633 140 644 645 cell_1rw
* cell instance $18909 m0 *1 26.085,163.8
X$18909 139 634 140 644 645 cell_1rw
* cell instance $18910 r0 *1 26.085,163.8
X$18910 139 635 140 644 645 cell_1rw
* cell instance $18911 m0 *1 26.085,166.53
X$18911 139 637 140 644 645 cell_1rw
* cell instance $18912 r0 *1 26.085,166.53
X$18912 139 636 140 644 645 cell_1rw
* cell instance $18913 m0 *1 26.085,169.26
X$18913 139 639 140 644 645 cell_1rw
* cell instance $18914 r0 *1 26.085,169.26
X$18914 139 638 140 644 645 cell_1rw
* cell instance $18915 m0 *1 26.085,171.99
X$18915 139 640 140 644 645 cell_1rw
* cell instance $18916 r0 *1 26.085,171.99
X$18916 139 641 140 644 645 cell_1rw
* cell instance $18917 m0 *1 26.085,174.72
X$18917 139 642 140 644 645 cell_1rw
* cell instance $18918 r0 *1 26.085,174.72
X$18918 139 643 140 644 645 cell_1rw
* cell instance $18919 r0 *1 26.79,87.36
X$18919 141 322 142 644 645 cell_1rw
* cell instance $18920 m0 *1 26.79,90.09
X$18920 141 581 142 644 645 cell_1rw
* cell instance $18921 r0 *1 26.79,90.09
X$18921 141 580 142 644 645 cell_1rw
* cell instance $18922 m0 *1 26.79,92.82
X$18922 141 583 142 644 645 cell_1rw
* cell instance $18923 r0 *1 26.79,92.82
X$18923 141 582 142 644 645 cell_1rw
* cell instance $18924 m0 *1 26.79,95.55
X$18924 141 584 142 644 645 cell_1rw
* cell instance $18925 r0 *1 26.79,95.55
X$18925 141 585 142 644 645 cell_1rw
* cell instance $18926 m0 *1 26.79,98.28
X$18926 141 586 142 644 645 cell_1rw
* cell instance $18927 r0 *1 26.79,98.28
X$18927 141 587 142 644 645 cell_1rw
* cell instance $18928 m0 *1 26.79,101.01
X$18928 141 588 142 644 645 cell_1rw
* cell instance $18929 r0 *1 26.79,101.01
X$18929 141 589 142 644 645 cell_1rw
* cell instance $18930 m0 *1 26.79,103.74
X$18930 141 590 142 644 645 cell_1rw
* cell instance $18931 r0 *1 26.79,103.74
X$18931 141 591 142 644 645 cell_1rw
* cell instance $18932 m0 *1 26.79,106.47
X$18932 141 593 142 644 645 cell_1rw
* cell instance $18933 r0 *1 26.79,106.47
X$18933 141 592 142 644 645 cell_1rw
* cell instance $18934 m0 *1 26.79,109.2
X$18934 141 594 142 644 645 cell_1rw
* cell instance $18935 r0 *1 26.79,109.2
X$18935 141 595 142 644 645 cell_1rw
* cell instance $18936 m0 *1 26.79,111.93
X$18936 141 597 142 644 645 cell_1rw
* cell instance $18937 r0 *1 26.79,111.93
X$18937 141 596 142 644 645 cell_1rw
* cell instance $18938 m0 *1 26.79,114.66
X$18938 141 598 142 644 645 cell_1rw
* cell instance $18939 m0 *1 26.79,117.39
X$18939 141 600 142 644 645 cell_1rw
* cell instance $18940 r0 *1 26.79,114.66
X$18940 141 599 142 644 645 cell_1rw
* cell instance $18941 r0 *1 26.79,117.39
X$18941 141 601 142 644 645 cell_1rw
* cell instance $18942 m0 *1 26.79,120.12
X$18942 141 602 142 644 645 cell_1rw
* cell instance $18943 r0 *1 26.79,120.12
X$18943 141 603 142 644 645 cell_1rw
* cell instance $18944 m0 *1 26.79,122.85
X$18944 141 604 142 644 645 cell_1rw
* cell instance $18945 r0 *1 26.79,122.85
X$18945 141 605 142 644 645 cell_1rw
* cell instance $18946 m0 *1 26.79,125.58
X$18946 141 606 142 644 645 cell_1rw
* cell instance $18947 r0 *1 26.79,125.58
X$18947 141 607 142 644 645 cell_1rw
* cell instance $18948 m0 *1 26.79,128.31
X$18948 141 609 142 644 645 cell_1rw
* cell instance $18949 r0 *1 26.79,128.31
X$18949 141 608 142 644 645 cell_1rw
* cell instance $18950 m0 *1 26.79,131.04
X$18950 141 610 142 644 645 cell_1rw
* cell instance $18951 m0 *1 26.79,133.77
X$18951 141 612 142 644 645 cell_1rw
* cell instance $18952 r0 *1 26.79,131.04
X$18952 141 611 142 644 645 cell_1rw
* cell instance $18953 r0 *1 26.79,133.77
X$18953 141 613 142 644 645 cell_1rw
* cell instance $18954 m0 *1 26.79,136.5
X$18954 141 615 142 644 645 cell_1rw
* cell instance $18955 m0 *1 26.79,139.23
X$18955 141 617 142 644 645 cell_1rw
* cell instance $18956 r0 *1 26.79,136.5
X$18956 141 614 142 644 645 cell_1rw
* cell instance $18957 r0 *1 26.79,139.23
X$18957 141 616 142 644 645 cell_1rw
* cell instance $18958 m0 *1 26.79,141.96
X$18958 141 618 142 644 645 cell_1rw
* cell instance $18959 m0 *1 26.79,144.69
X$18959 141 620 142 644 645 cell_1rw
* cell instance $18960 r0 *1 26.79,141.96
X$18960 141 619 142 644 645 cell_1rw
* cell instance $18961 r0 *1 26.79,144.69
X$18961 141 621 142 644 645 cell_1rw
* cell instance $18962 m0 *1 26.79,147.42
X$18962 141 622 142 644 645 cell_1rw
* cell instance $18963 r0 *1 26.79,147.42
X$18963 141 623 142 644 645 cell_1rw
* cell instance $18964 m0 *1 26.79,150.15
X$18964 141 624 142 644 645 cell_1rw
* cell instance $18965 r0 *1 26.79,150.15
X$18965 141 625 142 644 645 cell_1rw
* cell instance $18966 m0 *1 26.79,152.88
X$18966 141 626 142 644 645 cell_1rw
* cell instance $18967 r0 *1 26.79,152.88
X$18967 141 627 142 644 645 cell_1rw
* cell instance $18968 m0 *1 26.79,155.61
X$18968 141 628 142 644 645 cell_1rw
* cell instance $18969 r0 *1 26.79,155.61
X$18969 141 629 142 644 645 cell_1rw
* cell instance $18970 m0 *1 26.79,158.34
X$18970 141 630 142 644 645 cell_1rw
* cell instance $18971 r0 *1 26.79,158.34
X$18971 141 631 142 644 645 cell_1rw
* cell instance $18972 m0 *1 26.79,161.07
X$18972 141 632 142 644 645 cell_1rw
* cell instance $18973 m0 *1 26.79,163.8
X$18973 141 634 142 644 645 cell_1rw
* cell instance $18974 r0 *1 26.79,161.07
X$18974 141 633 142 644 645 cell_1rw
* cell instance $18975 r0 *1 26.79,163.8
X$18975 141 635 142 644 645 cell_1rw
* cell instance $18976 m0 *1 26.79,166.53
X$18976 141 637 142 644 645 cell_1rw
* cell instance $18977 r0 *1 26.79,166.53
X$18977 141 636 142 644 645 cell_1rw
* cell instance $18978 m0 *1 26.79,169.26
X$18978 141 639 142 644 645 cell_1rw
* cell instance $18979 r0 *1 26.79,169.26
X$18979 141 638 142 644 645 cell_1rw
* cell instance $18980 m0 *1 26.79,171.99
X$18980 141 640 142 644 645 cell_1rw
* cell instance $18981 r0 *1 26.79,171.99
X$18981 141 641 142 644 645 cell_1rw
* cell instance $18982 m0 *1 26.79,174.72
X$18982 141 642 142 644 645 cell_1rw
* cell instance $18983 r0 *1 26.79,174.72
X$18983 141 643 142 644 645 cell_1rw
* cell instance $18984 r0 *1 27.495,87.36
X$18984 143 322 144 644 645 cell_1rw
* cell instance $18985 m0 *1 27.495,90.09
X$18985 143 581 144 644 645 cell_1rw
* cell instance $18986 r0 *1 27.495,90.09
X$18986 143 580 144 644 645 cell_1rw
* cell instance $18987 m0 *1 27.495,92.82
X$18987 143 583 144 644 645 cell_1rw
* cell instance $18988 r0 *1 27.495,92.82
X$18988 143 582 144 644 645 cell_1rw
* cell instance $18989 m0 *1 27.495,95.55
X$18989 143 584 144 644 645 cell_1rw
* cell instance $18990 r0 *1 27.495,95.55
X$18990 143 585 144 644 645 cell_1rw
* cell instance $18991 m0 *1 27.495,98.28
X$18991 143 586 144 644 645 cell_1rw
* cell instance $18992 r0 *1 27.495,98.28
X$18992 143 587 144 644 645 cell_1rw
* cell instance $18993 m0 *1 27.495,101.01
X$18993 143 588 144 644 645 cell_1rw
* cell instance $18994 r0 *1 27.495,101.01
X$18994 143 589 144 644 645 cell_1rw
* cell instance $18995 m0 *1 27.495,103.74
X$18995 143 590 144 644 645 cell_1rw
* cell instance $18996 r0 *1 27.495,103.74
X$18996 143 591 144 644 645 cell_1rw
* cell instance $18997 m0 *1 27.495,106.47
X$18997 143 593 144 644 645 cell_1rw
* cell instance $18998 r0 *1 27.495,106.47
X$18998 143 592 144 644 645 cell_1rw
* cell instance $18999 m0 *1 27.495,109.2
X$18999 143 594 144 644 645 cell_1rw
* cell instance $19000 m0 *1 27.495,111.93
X$19000 143 597 144 644 645 cell_1rw
* cell instance $19001 r0 *1 27.495,109.2
X$19001 143 595 144 644 645 cell_1rw
* cell instance $19002 m0 *1 27.495,114.66
X$19002 143 598 144 644 645 cell_1rw
* cell instance $19003 r0 *1 27.495,111.93
X$19003 143 596 144 644 645 cell_1rw
* cell instance $19004 r0 *1 27.495,114.66
X$19004 143 599 144 644 645 cell_1rw
* cell instance $19005 m0 *1 27.495,117.39
X$19005 143 600 144 644 645 cell_1rw
* cell instance $19006 r0 *1 27.495,117.39
X$19006 143 601 144 644 645 cell_1rw
* cell instance $19007 m0 *1 27.495,120.12
X$19007 143 602 144 644 645 cell_1rw
* cell instance $19008 r0 *1 27.495,120.12
X$19008 143 603 144 644 645 cell_1rw
* cell instance $19009 m0 *1 27.495,122.85
X$19009 143 604 144 644 645 cell_1rw
* cell instance $19010 r0 *1 27.495,122.85
X$19010 143 605 144 644 645 cell_1rw
* cell instance $19011 m0 *1 27.495,125.58
X$19011 143 606 144 644 645 cell_1rw
* cell instance $19012 r0 *1 27.495,125.58
X$19012 143 607 144 644 645 cell_1rw
* cell instance $19013 m0 *1 27.495,128.31
X$19013 143 609 144 644 645 cell_1rw
* cell instance $19014 m0 *1 27.495,131.04
X$19014 143 610 144 644 645 cell_1rw
* cell instance $19015 r0 *1 27.495,128.31
X$19015 143 608 144 644 645 cell_1rw
* cell instance $19016 r0 *1 27.495,131.04
X$19016 143 611 144 644 645 cell_1rw
* cell instance $19017 m0 *1 27.495,133.77
X$19017 143 612 144 644 645 cell_1rw
* cell instance $19018 r0 *1 27.495,133.77
X$19018 143 613 144 644 645 cell_1rw
* cell instance $19019 m0 *1 27.495,136.5
X$19019 143 615 144 644 645 cell_1rw
* cell instance $19020 r0 *1 27.495,136.5
X$19020 143 614 144 644 645 cell_1rw
* cell instance $19021 m0 *1 27.495,139.23
X$19021 143 617 144 644 645 cell_1rw
* cell instance $19022 r0 *1 27.495,139.23
X$19022 143 616 144 644 645 cell_1rw
* cell instance $19023 m0 *1 27.495,141.96
X$19023 143 618 144 644 645 cell_1rw
* cell instance $19024 m0 *1 27.495,144.69
X$19024 143 620 144 644 645 cell_1rw
* cell instance $19025 r0 *1 27.495,141.96
X$19025 143 619 144 644 645 cell_1rw
* cell instance $19026 r0 *1 27.495,144.69
X$19026 143 621 144 644 645 cell_1rw
* cell instance $19027 m0 *1 27.495,147.42
X$19027 143 622 144 644 645 cell_1rw
* cell instance $19028 r0 *1 27.495,147.42
X$19028 143 623 144 644 645 cell_1rw
* cell instance $19029 m0 *1 27.495,150.15
X$19029 143 624 144 644 645 cell_1rw
* cell instance $19030 r0 *1 27.495,150.15
X$19030 143 625 144 644 645 cell_1rw
* cell instance $19031 m0 *1 27.495,152.88
X$19031 143 626 144 644 645 cell_1rw
* cell instance $19032 r0 *1 27.495,152.88
X$19032 143 627 144 644 645 cell_1rw
* cell instance $19033 m0 *1 27.495,155.61
X$19033 143 628 144 644 645 cell_1rw
* cell instance $19034 m0 *1 27.495,158.34
X$19034 143 630 144 644 645 cell_1rw
* cell instance $19035 r0 *1 27.495,155.61
X$19035 143 629 144 644 645 cell_1rw
* cell instance $19036 r0 *1 27.495,158.34
X$19036 143 631 144 644 645 cell_1rw
* cell instance $19037 m0 *1 27.495,161.07
X$19037 143 632 144 644 645 cell_1rw
* cell instance $19038 r0 *1 27.495,161.07
X$19038 143 633 144 644 645 cell_1rw
* cell instance $19039 m0 *1 27.495,163.8
X$19039 143 634 144 644 645 cell_1rw
* cell instance $19040 r0 *1 27.495,163.8
X$19040 143 635 144 644 645 cell_1rw
* cell instance $19041 m0 *1 27.495,166.53
X$19041 143 637 144 644 645 cell_1rw
* cell instance $19042 r0 *1 27.495,166.53
X$19042 143 636 144 644 645 cell_1rw
* cell instance $19043 m0 *1 27.495,169.26
X$19043 143 639 144 644 645 cell_1rw
* cell instance $19044 r0 *1 27.495,169.26
X$19044 143 638 144 644 645 cell_1rw
* cell instance $19045 m0 *1 27.495,171.99
X$19045 143 640 144 644 645 cell_1rw
* cell instance $19046 r0 *1 27.495,171.99
X$19046 143 641 144 644 645 cell_1rw
* cell instance $19047 m0 *1 27.495,174.72
X$19047 143 642 144 644 645 cell_1rw
* cell instance $19048 r0 *1 27.495,174.72
X$19048 143 643 144 644 645 cell_1rw
* cell instance $19049 r0 *1 28.2,87.36
X$19049 145 322 146 644 645 cell_1rw
* cell instance $19050 m0 *1 28.2,90.09
X$19050 145 581 146 644 645 cell_1rw
* cell instance $19051 m0 *1 28.2,92.82
X$19051 145 583 146 644 645 cell_1rw
* cell instance $19052 r0 *1 28.2,90.09
X$19052 145 580 146 644 645 cell_1rw
* cell instance $19053 r0 *1 28.2,92.82
X$19053 145 582 146 644 645 cell_1rw
* cell instance $19054 m0 *1 28.2,95.55
X$19054 145 584 146 644 645 cell_1rw
* cell instance $19055 r0 *1 28.2,95.55
X$19055 145 585 146 644 645 cell_1rw
* cell instance $19056 m0 *1 28.2,98.28
X$19056 145 586 146 644 645 cell_1rw
* cell instance $19057 r0 *1 28.2,98.28
X$19057 145 587 146 644 645 cell_1rw
* cell instance $19058 m0 *1 28.2,101.01
X$19058 145 588 146 644 645 cell_1rw
* cell instance $19059 m0 *1 28.2,103.74
X$19059 145 590 146 644 645 cell_1rw
* cell instance $19060 r0 *1 28.2,101.01
X$19060 145 589 146 644 645 cell_1rw
* cell instance $19061 r0 *1 28.2,103.74
X$19061 145 591 146 644 645 cell_1rw
* cell instance $19062 m0 *1 28.2,106.47
X$19062 145 593 146 644 645 cell_1rw
* cell instance $19063 m0 *1 28.2,109.2
X$19063 145 594 146 644 645 cell_1rw
* cell instance $19064 r0 *1 28.2,106.47
X$19064 145 592 146 644 645 cell_1rw
* cell instance $19065 m0 *1 28.2,111.93
X$19065 145 597 146 644 645 cell_1rw
* cell instance $19066 r0 *1 28.2,109.2
X$19066 145 595 146 644 645 cell_1rw
* cell instance $19067 m0 *1 28.2,114.66
X$19067 145 598 146 644 645 cell_1rw
* cell instance $19068 r0 *1 28.2,111.93
X$19068 145 596 146 644 645 cell_1rw
* cell instance $19069 r0 *1 28.2,114.66
X$19069 145 599 146 644 645 cell_1rw
* cell instance $19070 m0 *1 28.2,117.39
X$19070 145 600 146 644 645 cell_1rw
* cell instance $19071 r0 *1 28.2,117.39
X$19071 145 601 146 644 645 cell_1rw
* cell instance $19072 m0 *1 28.2,120.12
X$19072 145 602 146 644 645 cell_1rw
* cell instance $19073 r0 *1 28.2,120.12
X$19073 145 603 146 644 645 cell_1rw
* cell instance $19074 m0 *1 28.2,122.85
X$19074 145 604 146 644 645 cell_1rw
* cell instance $19075 r0 *1 28.2,122.85
X$19075 145 605 146 644 645 cell_1rw
* cell instance $19076 m0 *1 28.2,125.58
X$19076 145 606 146 644 645 cell_1rw
* cell instance $19077 r0 *1 28.2,125.58
X$19077 145 607 146 644 645 cell_1rw
* cell instance $19078 m0 *1 28.2,128.31
X$19078 145 609 146 644 645 cell_1rw
* cell instance $19079 r0 *1 28.2,128.31
X$19079 145 608 146 644 645 cell_1rw
* cell instance $19080 m0 *1 28.2,131.04
X$19080 145 610 146 644 645 cell_1rw
* cell instance $19081 r0 *1 28.2,131.04
X$19081 145 611 146 644 645 cell_1rw
* cell instance $19082 m0 *1 28.2,133.77
X$19082 145 612 146 644 645 cell_1rw
* cell instance $19083 r0 *1 28.2,133.77
X$19083 145 613 146 644 645 cell_1rw
* cell instance $19084 m0 *1 28.2,136.5
X$19084 145 615 146 644 645 cell_1rw
* cell instance $19085 r0 *1 28.2,136.5
X$19085 145 614 146 644 645 cell_1rw
* cell instance $19086 m0 *1 28.2,139.23
X$19086 145 617 146 644 645 cell_1rw
* cell instance $19087 r0 *1 28.2,139.23
X$19087 145 616 146 644 645 cell_1rw
* cell instance $19088 m0 *1 28.2,141.96
X$19088 145 618 146 644 645 cell_1rw
* cell instance $19089 r0 *1 28.2,141.96
X$19089 145 619 146 644 645 cell_1rw
* cell instance $19090 m0 *1 28.2,144.69
X$19090 145 620 146 644 645 cell_1rw
* cell instance $19091 r0 *1 28.2,144.69
X$19091 145 621 146 644 645 cell_1rw
* cell instance $19092 m0 *1 28.2,147.42
X$19092 145 622 146 644 645 cell_1rw
* cell instance $19093 r0 *1 28.2,147.42
X$19093 145 623 146 644 645 cell_1rw
* cell instance $19094 m0 *1 28.2,150.15
X$19094 145 624 146 644 645 cell_1rw
* cell instance $19095 r0 *1 28.2,150.15
X$19095 145 625 146 644 645 cell_1rw
* cell instance $19096 m0 *1 28.2,152.88
X$19096 145 626 146 644 645 cell_1rw
* cell instance $19097 r0 *1 28.2,152.88
X$19097 145 627 146 644 645 cell_1rw
* cell instance $19098 m0 *1 28.2,155.61
X$19098 145 628 146 644 645 cell_1rw
* cell instance $19099 r0 *1 28.2,155.61
X$19099 145 629 146 644 645 cell_1rw
* cell instance $19100 m0 *1 28.2,158.34
X$19100 145 630 146 644 645 cell_1rw
* cell instance $19101 r0 *1 28.2,158.34
X$19101 145 631 146 644 645 cell_1rw
* cell instance $19102 m0 *1 28.2,161.07
X$19102 145 632 146 644 645 cell_1rw
* cell instance $19103 r0 *1 28.2,161.07
X$19103 145 633 146 644 645 cell_1rw
* cell instance $19104 m0 *1 28.2,163.8
X$19104 145 634 146 644 645 cell_1rw
* cell instance $19105 r0 *1 28.2,163.8
X$19105 145 635 146 644 645 cell_1rw
* cell instance $19106 m0 *1 28.2,166.53
X$19106 145 637 146 644 645 cell_1rw
* cell instance $19107 r0 *1 28.2,166.53
X$19107 145 636 146 644 645 cell_1rw
* cell instance $19108 m0 *1 28.2,169.26
X$19108 145 639 146 644 645 cell_1rw
* cell instance $19109 r0 *1 28.2,169.26
X$19109 145 638 146 644 645 cell_1rw
* cell instance $19110 m0 *1 28.2,171.99
X$19110 145 640 146 644 645 cell_1rw
* cell instance $19111 r0 *1 28.2,171.99
X$19111 145 641 146 644 645 cell_1rw
* cell instance $19112 m0 *1 28.2,174.72
X$19112 145 642 146 644 645 cell_1rw
* cell instance $19113 r0 *1 28.2,174.72
X$19113 145 643 146 644 645 cell_1rw
* cell instance $19114 r0 *1 28.905,87.36
X$19114 147 322 148 644 645 cell_1rw
* cell instance $19115 m0 *1 28.905,90.09
X$19115 147 581 148 644 645 cell_1rw
* cell instance $19116 r0 *1 28.905,90.09
X$19116 147 580 148 644 645 cell_1rw
* cell instance $19117 m0 *1 28.905,92.82
X$19117 147 583 148 644 645 cell_1rw
* cell instance $19118 r0 *1 28.905,92.82
X$19118 147 582 148 644 645 cell_1rw
* cell instance $19119 m0 *1 28.905,95.55
X$19119 147 584 148 644 645 cell_1rw
* cell instance $19120 r0 *1 28.905,95.55
X$19120 147 585 148 644 645 cell_1rw
* cell instance $19121 m0 *1 28.905,98.28
X$19121 147 586 148 644 645 cell_1rw
* cell instance $19122 m0 *1 28.905,101.01
X$19122 147 588 148 644 645 cell_1rw
* cell instance $19123 r0 *1 28.905,98.28
X$19123 147 587 148 644 645 cell_1rw
* cell instance $19124 m0 *1 28.905,103.74
X$19124 147 590 148 644 645 cell_1rw
* cell instance $19125 r0 *1 28.905,101.01
X$19125 147 589 148 644 645 cell_1rw
* cell instance $19126 r0 *1 28.905,103.74
X$19126 147 591 148 644 645 cell_1rw
* cell instance $19127 m0 *1 28.905,106.47
X$19127 147 593 148 644 645 cell_1rw
* cell instance $19128 r0 *1 28.905,106.47
X$19128 147 592 148 644 645 cell_1rw
* cell instance $19129 m0 *1 28.905,109.2
X$19129 147 594 148 644 645 cell_1rw
* cell instance $19130 r0 *1 28.905,109.2
X$19130 147 595 148 644 645 cell_1rw
* cell instance $19131 m0 *1 28.905,111.93
X$19131 147 597 148 644 645 cell_1rw
* cell instance $19132 m0 *1 28.905,114.66
X$19132 147 598 148 644 645 cell_1rw
* cell instance $19133 r0 *1 28.905,111.93
X$19133 147 596 148 644 645 cell_1rw
* cell instance $19134 r0 *1 28.905,114.66
X$19134 147 599 148 644 645 cell_1rw
* cell instance $19135 m0 *1 28.905,117.39
X$19135 147 600 148 644 645 cell_1rw
* cell instance $19136 r0 *1 28.905,117.39
X$19136 147 601 148 644 645 cell_1rw
* cell instance $19137 m0 *1 28.905,120.12
X$19137 147 602 148 644 645 cell_1rw
* cell instance $19138 r0 *1 28.905,120.12
X$19138 147 603 148 644 645 cell_1rw
* cell instance $19139 m0 *1 28.905,122.85
X$19139 147 604 148 644 645 cell_1rw
* cell instance $19140 r0 *1 28.905,122.85
X$19140 147 605 148 644 645 cell_1rw
* cell instance $19141 m0 *1 28.905,125.58
X$19141 147 606 148 644 645 cell_1rw
* cell instance $19142 m0 *1 28.905,128.31
X$19142 147 609 148 644 645 cell_1rw
* cell instance $19143 r0 *1 28.905,125.58
X$19143 147 607 148 644 645 cell_1rw
* cell instance $19144 r0 *1 28.905,128.31
X$19144 147 608 148 644 645 cell_1rw
* cell instance $19145 m0 *1 28.905,131.04
X$19145 147 610 148 644 645 cell_1rw
* cell instance $19146 r0 *1 28.905,131.04
X$19146 147 611 148 644 645 cell_1rw
* cell instance $19147 m0 *1 28.905,133.77
X$19147 147 612 148 644 645 cell_1rw
* cell instance $19148 r0 *1 28.905,133.77
X$19148 147 613 148 644 645 cell_1rw
* cell instance $19149 m0 *1 28.905,136.5
X$19149 147 615 148 644 645 cell_1rw
* cell instance $19150 m0 *1 28.905,139.23
X$19150 147 617 148 644 645 cell_1rw
* cell instance $19151 r0 *1 28.905,136.5
X$19151 147 614 148 644 645 cell_1rw
* cell instance $19152 r0 *1 28.905,139.23
X$19152 147 616 148 644 645 cell_1rw
* cell instance $19153 m0 *1 28.905,141.96
X$19153 147 618 148 644 645 cell_1rw
* cell instance $19154 r0 *1 28.905,141.96
X$19154 147 619 148 644 645 cell_1rw
* cell instance $19155 m0 *1 28.905,144.69
X$19155 147 620 148 644 645 cell_1rw
* cell instance $19156 r0 *1 28.905,144.69
X$19156 147 621 148 644 645 cell_1rw
* cell instance $19157 m0 *1 28.905,147.42
X$19157 147 622 148 644 645 cell_1rw
* cell instance $19158 r0 *1 28.905,147.42
X$19158 147 623 148 644 645 cell_1rw
* cell instance $19159 m0 *1 28.905,150.15
X$19159 147 624 148 644 645 cell_1rw
* cell instance $19160 r0 *1 28.905,150.15
X$19160 147 625 148 644 645 cell_1rw
* cell instance $19161 m0 *1 28.905,152.88
X$19161 147 626 148 644 645 cell_1rw
* cell instance $19162 r0 *1 28.905,152.88
X$19162 147 627 148 644 645 cell_1rw
* cell instance $19163 m0 *1 28.905,155.61
X$19163 147 628 148 644 645 cell_1rw
* cell instance $19164 r0 *1 28.905,155.61
X$19164 147 629 148 644 645 cell_1rw
* cell instance $19165 m0 *1 28.905,158.34
X$19165 147 630 148 644 645 cell_1rw
* cell instance $19166 r0 *1 28.905,158.34
X$19166 147 631 148 644 645 cell_1rw
* cell instance $19167 m0 *1 28.905,161.07
X$19167 147 632 148 644 645 cell_1rw
* cell instance $19168 r0 *1 28.905,161.07
X$19168 147 633 148 644 645 cell_1rw
* cell instance $19169 m0 *1 28.905,163.8
X$19169 147 634 148 644 645 cell_1rw
* cell instance $19170 r0 *1 28.905,163.8
X$19170 147 635 148 644 645 cell_1rw
* cell instance $19171 m0 *1 28.905,166.53
X$19171 147 637 148 644 645 cell_1rw
* cell instance $19172 r0 *1 28.905,166.53
X$19172 147 636 148 644 645 cell_1rw
* cell instance $19173 m0 *1 28.905,169.26
X$19173 147 639 148 644 645 cell_1rw
* cell instance $19174 r0 *1 28.905,169.26
X$19174 147 638 148 644 645 cell_1rw
* cell instance $19175 m0 *1 28.905,171.99
X$19175 147 640 148 644 645 cell_1rw
* cell instance $19176 r0 *1 28.905,171.99
X$19176 147 641 148 644 645 cell_1rw
* cell instance $19177 m0 *1 28.905,174.72
X$19177 147 642 148 644 645 cell_1rw
* cell instance $19178 r0 *1 28.905,174.72
X$19178 147 643 148 644 645 cell_1rw
* cell instance $19179 r0 *1 29.61,87.36
X$19179 149 322 150 644 645 cell_1rw
* cell instance $19180 m0 *1 29.61,90.09
X$19180 149 581 150 644 645 cell_1rw
* cell instance $19181 r0 *1 29.61,90.09
X$19181 149 580 150 644 645 cell_1rw
* cell instance $19182 m0 *1 29.61,92.82
X$19182 149 583 150 644 645 cell_1rw
* cell instance $19183 m0 *1 29.61,95.55
X$19183 149 584 150 644 645 cell_1rw
* cell instance $19184 r0 *1 29.61,92.82
X$19184 149 582 150 644 645 cell_1rw
* cell instance $19185 r0 *1 29.61,95.55
X$19185 149 585 150 644 645 cell_1rw
* cell instance $19186 m0 *1 29.61,98.28
X$19186 149 586 150 644 645 cell_1rw
* cell instance $19187 m0 *1 29.61,101.01
X$19187 149 588 150 644 645 cell_1rw
* cell instance $19188 r0 *1 29.61,98.28
X$19188 149 587 150 644 645 cell_1rw
* cell instance $19189 r0 *1 29.61,101.01
X$19189 149 589 150 644 645 cell_1rw
* cell instance $19190 m0 *1 29.61,103.74
X$19190 149 590 150 644 645 cell_1rw
* cell instance $19191 r0 *1 29.61,103.74
X$19191 149 591 150 644 645 cell_1rw
* cell instance $19192 m0 *1 29.61,106.47
X$19192 149 593 150 644 645 cell_1rw
* cell instance $19193 m0 *1 29.61,109.2
X$19193 149 594 150 644 645 cell_1rw
* cell instance $19194 r0 *1 29.61,106.47
X$19194 149 592 150 644 645 cell_1rw
* cell instance $19195 r0 *1 29.61,109.2
X$19195 149 595 150 644 645 cell_1rw
* cell instance $19196 m0 *1 29.61,111.93
X$19196 149 597 150 644 645 cell_1rw
* cell instance $19197 r0 *1 29.61,111.93
X$19197 149 596 150 644 645 cell_1rw
* cell instance $19198 m0 *1 29.61,114.66
X$19198 149 598 150 644 645 cell_1rw
* cell instance $19199 r0 *1 29.61,114.66
X$19199 149 599 150 644 645 cell_1rw
* cell instance $19200 m0 *1 29.61,117.39
X$19200 149 600 150 644 645 cell_1rw
* cell instance $19201 m0 *1 29.61,120.12
X$19201 149 602 150 644 645 cell_1rw
* cell instance $19202 r0 *1 29.61,117.39
X$19202 149 601 150 644 645 cell_1rw
* cell instance $19203 r0 *1 29.61,120.12
X$19203 149 603 150 644 645 cell_1rw
* cell instance $19204 m0 *1 29.61,122.85
X$19204 149 604 150 644 645 cell_1rw
* cell instance $19205 r0 *1 29.61,122.85
X$19205 149 605 150 644 645 cell_1rw
* cell instance $19206 m0 *1 29.61,125.58
X$19206 149 606 150 644 645 cell_1rw
* cell instance $19207 m0 *1 29.61,128.31
X$19207 149 609 150 644 645 cell_1rw
* cell instance $19208 r0 *1 29.61,125.58
X$19208 149 607 150 644 645 cell_1rw
* cell instance $19209 r0 *1 29.61,128.31
X$19209 149 608 150 644 645 cell_1rw
* cell instance $19210 m0 *1 29.61,131.04
X$19210 149 610 150 644 645 cell_1rw
* cell instance $19211 r0 *1 29.61,131.04
X$19211 149 611 150 644 645 cell_1rw
* cell instance $19212 m0 *1 29.61,133.77
X$19212 149 612 150 644 645 cell_1rw
* cell instance $19213 r0 *1 29.61,133.77
X$19213 149 613 150 644 645 cell_1rw
* cell instance $19214 m0 *1 29.61,136.5
X$19214 149 615 150 644 645 cell_1rw
* cell instance $19215 m0 *1 29.61,139.23
X$19215 149 617 150 644 645 cell_1rw
* cell instance $19216 r0 *1 29.61,136.5
X$19216 149 614 150 644 645 cell_1rw
* cell instance $19217 r0 *1 29.61,139.23
X$19217 149 616 150 644 645 cell_1rw
* cell instance $19218 m0 *1 29.61,141.96
X$19218 149 618 150 644 645 cell_1rw
* cell instance $19219 r0 *1 29.61,141.96
X$19219 149 619 150 644 645 cell_1rw
* cell instance $19220 m0 *1 29.61,144.69
X$19220 149 620 150 644 645 cell_1rw
* cell instance $19221 r0 *1 29.61,144.69
X$19221 149 621 150 644 645 cell_1rw
* cell instance $19222 m0 *1 29.61,147.42
X$19222 149 622 150 644 645 cell_1rw
* cell instance $19223 r0 *1 29.61,147.42
X$19223 149 623 150 644 645 cell_1rw
* cell instance $19224 m0 *1 29.61,150.15
X$19224 149 624 150 644 645 cell_1rw
* cell instance $19225 m0 *1 29.61,152.88
X$19225 149 626 150 644 645 cell_1rw
* cell instance $19226 r0 *1 29.61,150.15
X$19226 149 625 150 644 645 cell_1rw
* cell instance $19227 r0 *1 29.61,152.88
X$19227 149 627 150 644 645 cell_1rw
* cell instance $19228 m0 *1 29.61,155.61
X$19228 149 628 150 644 645 cell_1rw
* cell instance $19229 r0 *1 29.61,155.61
X$19229 149 629 150 644 645 cell_1rw
* cell instance $19230 m0 *1 29.61,158.34
X$19230 149 630 150 644 645 cell_1rw
* cell instance $19231 r0 *1 29.61,158.34
X$19231 149 631 150 644 645 cell_1rw
* cell instance $19232 m0 *1 29.61,161.07
X$19232 149 632 150 644 645 cell_1rw
* cell instance $19233 m0 *1 29.61,163.8
X$19233 149 634 150 644 645 cell_1rw
* cell instance $19234 r0 *1 29.61,161.07
X$19234 149 633 150 644 645 cell_1rw
* cell instance $19235 r0 *1 29.61,163.8
X$19235 149 635 150 644 645 cell_1rw
* cell instance $19236 m0 *1 29.61,166.53
X$19236 149 637 150 644 645 cell_1rw
* cell instance $19237 r0 *1 29.61,166.53
X$19237 149 636 150 644 645 cell_1rw
* cell instance $19238 m0 *1 29.61,169.26
X$19238 149 639 150 644 645 cell_1rw
* cell instance $19239 r0 *1 29.61,169.26
X$19239 149 638 150 644 645 cell_1rw
* cell instance $19240 m0 *1 29.61,171.99
X$19240 149 640 150 644 645 cell_1rw
* cell instance $19241 r0 *1 29.61,171.99
X$19241 149 641 150 644 645 cell_1rw
* cell instance $19242 m0 *1 29.61,174.72
X$19242 149 642 150 644 645 cell_1rw
* cell instance $19243 r0 *1 29.61,174.72
X$19243 149 643 150 644 645 cell_1rw
* cell instance $19244 r0 *1 30.315,87.36
X$19244 151 322 152 644 645 cell_1rw
* cell instance $19245 m0 *1 30.315,90.09
X$19245 151 581 152 644 645 cell_1rw
* cell instance $19246 r0 *1 30.315,90.09
X$19246 151 580 152 644 645 cell_1rw
* cell instance $19247 m0 *1 30.315,92.82
X$19247 151 583 152 644 645 cell_1rw
* cell instance $19248 r0 *1 30.315,92.82
X$19248 151 582 152 644 645 cell_1rw
* cell instance $19249 m0 *1 30.315,95.55
X$19249 151 584 152 644 645 cell_1rw
* cell instance $19250 r0 *1 30.315,95.55
X$19250 151 585 152 644 645 cell_1rw
* cell instance $19251 m0 *1 30.315,98.28
X$19251 151 586 152 644 645 cell_1rw
* cell instance $19252 r0 *1 30.315,98.28
X$19252 151 587 152 644 645 cell_1rw
* cell instance $19253 m0 *1 30.315,101.01
X$19253 151 588 152 644 645 cell_1rw
* cell instance $19254 r0 *1 30.315,101.01
X$19254 151 589 152 644 645 cell_1rw
* cell instance $19255 m0 *1 30.315,103.74
X$19255 151 590 152 644 645 cell_1rw
* cell instance $19256 r0 *1 30.315,103.74
X$19256 151 591 152 644 645 cell_1rw
* cell instance $19257 m0 *1 30.315,106.47
X$19257 151 593 152 644 645 cell_1rw
* cell instance $19258 r0 *1 30.315,106.47
X$19258 151 592 152 644 645 cell_1rw
* cell instance $19259 m0 *1 30.315,109.2
X$19259 151 594 152 644 645 cell_1rw
* cell instance $19260 m0 *1 30.315,111.93
X$19260 151 597 152 644 645 cell_1rw
* cell instance $19261 r0 *1 30.315,109.2
X$19261 151 595 152 644 645 cell_1rw
* cell instance $19262 r0 *1 30.315,111.93
X$19262 151 596 152 644 645 cell_1rw
* cell instance $19263 m0 *1 30.315,114.66
X$19263 151 598 152 644 645 cell_1rw
* cell instance $19264 m0 *1 30.315,117.39
X$19264 151 600 152 644 645 cell_1rw
* cell instance $19265 r0 *1 30.315,114.66
X$19265 151 599 152 644 645 cell_1rw
* cell instance $19266 r0 *1 30.315,117.39
X$19266 151 601 152 644 645 cell_1rw
* cell instance $19267 m0 *1 30.315,120.12
X$19267 151 602 152 644 645 cell_1rw
* cell instance $19268 r0 *1 30.315,120.12
X$19268 151 603 152 644 645 cell_1rw
* cell instance $19269 m0 *1 30.315,122.85
X$19269 151 604 152 644 645 cell_1rw
* cell instance $19270 r0 *1 30.315,122.85
X$19270 151 605 152 644 645 cell_1rw
* cell instance $19271 m0 *1 30.315,125.58
X$19271 151 606 152 644 645 cell_1rw
* cell instance $19272 r0 *1 30.315,125.58
X$19272 151 607 152 644 645 cell_1rw
* cell instance $19273 m0 *1 30.315,128.31
X$19273 151 609 152 644 645 cell_1rw
* cell instance $19274 r0 *1 30.315,128.31
X$19274 151 608 152 644 645 cell_1rw
* cell instance $19275 m0 *1 30.315,131.04
X$19275 151 610 152 644 645 cell_1rw
* cell instance $19276 r0 *1 30.315,131.04
X$19276 151 611 152 644 645 cell_1rw
* cell instance $19277 m0 *1 30.315,133.77
X$19277 151 612 152 644 645 cell_1rw
* cell instance $19278 r0 *1 30.315,133.77
X$19278 151 613 152 644 645 cell_1rw
* cell instance $19279 m0 *1 30.315,136.5
X$19279 151 615 152 644 645 cell_1rw
* cell instance $19280 r0 *1 30.315,136.5
X$19280 151 614 152 644 645 cell_1rw
* cell instance $19281 m0 *1 30.315,139.23
X$19281 151 617 152 644 645 cell_1rw
* cell instance $19282 r0 *1 30.315,139.23
X$19282 151 616 152 644 645 cell_1rw
* cell instance $19283 m0 *1 30.315,141.96
X$19283 151 618 152 644 645 cell_1rw
* cell instance $19284 r0 *1 30.315,141.96
X$19284 151 619 152 644 645 cell_1rw
* cell instance $19285 m0 *1 30.315,144.69
X$19285 151 620 152 644 645 cell_1rw
* cell instance $19286 r0 *1 30.315,144.69
X$19286 151 621 152 644 645 cell_1rw
* cell instance $19287 m0 *1 30.315,147.42
X$19287 151 622 152 644 645 cell_1rw
* cell instance $19288 m0 *1 30.315,150.15
X$19288 151 624 152 644 645 cell_1rw
* cell instance $19289 r0 *1 30.315,147.42
X$19289 151 623 152 644 645 cell_1rw
* cell instance $19290 m0 *1 30.315,152.88
X$19290 151 626 152 644 645 cell_1rw
* cell instance $19291 r0 *1 30.315,150.15
X$19291 151 625 152 644 645 cell_1rw
* cell instance $19292 r0 *1 30.315,152.88
X$19292 151 627 152 644 645 cell_1rw
* cell instance $19293 m0 *1 30.315,155.61
X$19293 151 628 152 644 645 cell_1rw
* cell instance $19294 r0 *1 30.315,155.61
X$19294 151 629 152 644 645 cell_1rw
* cell instance $19295 m0 *1 30.315,158.34
X$19295 151 630 152 644 645 cell_1rw
* cell instance $19296 r0 *1 30.315,158.34
X$19296 151 631 152 644 645 cell_1rw
* cell instance $19297 m0 *1 30.315,161.07
X$19297 151 632 152 644 645 cell_1rw
* cell instance $19298 m0 *1 30.315,163.8
X$19298 151 634 152 644 645 cell_1rw
* cell instance $19299 r0 *1 30.315,161.07
X$19299 151 633 152 644 645 cell_1rw
* cell instance $19300 r0 *1 30.315,163.8
X$19300 151 635 152 644 645 cell_1rw
* cell instance $19301 m0 *1 30.315,166.53
X$19301 151 637 152 644 645 cell_1rw
* cell instance $19302 r0 *1 30.315,166.53
X$19302 151 636 152 644 645 cell_1rw
* cell instance $19303 m0 *1 30.315,169.26
X$19303 151 639 152 644 645 cell_1rw
* cell instance $19304 m0 *1 30.315,171.99
X$19304 151 640 152 644 645 cell_1rw
* cell instance $19305 r0 *1 30.315,169.26
X$19305 151 638 152 644 645 cell_1rw
* cell instance $19306 r0 *1 30.315,171.99
X$19306 151 641 152 644 645 cell_1rw
* cell instance $19307 m0 *1 30.315,174.72
X$19307 151 642 152 644 645 cell_1rw
* cell instance $19308 r0 *1 30.315,174.72
X$19308 151 643 152 644 645 cell_1rw
* cell instance $19309 r0 *1 31.02,87.36
X$19309 153 322 154 644 645 cell_1rw
* cell instance $19310 m0 *1 31.02,90.09
X$19310 153 581 154 644 645 cell_1rw
* cell instance $19311 r0 *1 31.02,90.09
X$19311 153 580 154 644 645 cell_1rw
* cell instance $19312 m0 *1 31.02,92.82
X$19312 153 583 154 644 645 cell_1rw
* cell instance $19313 r0 *1 31.02,92.82
X$19313 153 582 154 644 645 cell_1rw
* cell instance $19314 m0 *1 31.02,95.55
X$19314 153 584 154 644 645 cell_1rw
* cell instance $19315 r0 *1 31.02,95.55
X$19315 153 585 154 644 645 cell_1rw
* cell instance $19316 m0 *1 31.02,98.28
X$19316 153 586 154 644 645 cell_1rw
* cell instance $19317 r0 *1 31.02,98.28
X$19317 153 587 154 644 645 cell_1rw
* cell instance $19318 m0 *1 31.02,101.01
X$19318 153 588 154 644 645 cell_1rw
* cell instance $19319 r0 *1 31.02,101.01
X$19319 153 589 154 644 645 cell_1rw
* cell instance $19320 m0 *1 31.02,103.74
X$19320 153 590 154 644 645 cell_1rw
* cell instance $19321 r0 *1 31.02,103.74
X$19321 153 591 154 644 645 cell_1rw
* cell instance $19322 m0 *1 31.02,106.47
X$19322 153 593 154 644 645 cell_1rw
* cell instance $19323 r0 *1 31.02,106.47
X$19323 153 592 154 644 645 cell_1rw
* cell instance $19324 m0 *1 31.02,109.2
X$19324 153 594 154 644 645 cell_1rw
* cell instance $19325 r0 *1 31.02,109.2
X$19325 153 595 154 644 645 cell_1rw
* cell instance $19326 m0 *1 31.02,111.93
X$19326 153 597 154 644 645 cell_1rw
* cell instance $19327 r0 *1 31.02,111.93
X$19327 153 596 154 644 645 cell_1rw
* cell instance $19328 m0 *1 31.02,114.66
X$19328 153 598 154 644 645 cell_1rw
* cell instance $19329 r0 *1 31.02,114.66
X$19329 153 599 154 644 645 cell_1rw
* cell instance $19330 m0 *1 31.02,117.39
X$19330 153 600 154 644 645 cell_1rw
* cell instance $19331 r0 *1 31.02,117.39
X$19331 153 601 154 644 645 cell_1rw
* cell instance $19332 m0 *1 31.02,120.12
X$19332 153 602 154 644 645 cell_1rw
* cell instance $19333 r0 *1 31.02,120.12
X$19333 153 603 154 644 645 cell_1rw
* cell instance $19334 m0 *1 31.02,122.85
X$19334 153 604 154 644 645 cell_1rw
* cell instance $19335 r0 *1 31.02,122.85
X$19335 153 605 154 644 645 cell_1rw
* cell instance $19336 m0 *1 31.02,125.58
X$19336 153 606 154 644 645 cell_1rw
* cell instance $19337 r0 *1 31.02,125.58
X$19337 153 607 154 644 645 cell_1rw
* cell instance $19338 m0 *1 31.02,128.31
X$19338 153 609 154 644 645 cell_1rw
* cell instance $19339 r0 *1 31.02,128.31
X$19339 153 608 154 644 645 cell_1rw
* cell instance $19340 m0 *1 31.02,131.04
X$19340 153 610 154 644 645 cell_1rw
* cell instance $19341 r0 *1 31.02,131.04
X$19341 153 611 154 644 645 cell_1rw
* cell instance $19342 m0 *1 31.02,133.77
X$19342 153 612 154 644 645 cell_1rw
* cell instance $19343 r0 *1 31.02,133.77
X$19343 153 613 154 644 645 cell_1rw
* cell instance $19344 m0 *1 31.02,136.5
X$19344 153 615 154 644 645 cell_1rw
* cell instance $19345 r0 *1 31.02,136.5
X$19345 153 614 154 644 645 cell_1rw
* cell instance $19346 m0 *1 31.02,139.23
X$19346 153 617 154 644 645 cell_1rw
* cell instance $19347 r0 *1 31.02,139.23
X$19347 153 616 154 644 645 cell_1rw
* cell instance $19348 m0 *1 31.02,141.96
X$19348 153 618 154 644 645 cell_1rw
* cell instance $19349 r0 *1 31.02,141.96
X$19349 153 619 154 644 645 cell_1rw
* cell instance $19350 m0 *1 31.02,144.69
X$19350 153 620 154 644 645 cell_1rw
* cell instance $19351 r0 *1 31.02,144.69
X$19351 153 621 154 644 645 cell_1rw
* cell instance $19352 m0 *1 31.02,147.42
X$19352 153 622 154 644 645 cell_1rw
* cell instance $19353 r0 *1 31.02,147.42
X$19353 153 623 154 644 645 cell_1rw
* cell instance $19354 m0 *1 31.02,150.15
X$19354 153 624 154 644 645 cell_1rw
* cell instance $19355 r0 *1 31.02,150.15
X$19355 153 625 154 644 645 cell_1rw
* cell instance $19356 m0 *1 31.02,152.88
X$19356 153 626 154 644 645 cell_1rw
* cell instance $19357 r0 *1 31.02,152.88
X$19357 153 627 154 644 645 cell_1rw
* cell instance $19358 m0 *1 31.02,155.61
X$19358 153 628 154 644 645 cell_1rw
* cell instance $19359 r0 *1 31.02,155.61
X$19359 153 629 154 644 645 cell_1rw
* cell instance $19360 m0 *1 31.02,158.34
X$19360 153 630 154 644 645 cell_1rw
* cell instance $19361 r0 *1 31.02,158.34
X$19361 153 631 154 644 645 cell_1rw
* cell instance $19362 m0 *1 31.02,161.07
X$19362 153 632 154 644 645 cell_1rw
* cell instance $19363 r0 *1 31.02,161.07
X$19363 153 633 154 644 645 cell_1rw
* cell instance $19364 m0 *1 31.02,163.8
X$19364 153 634 154 644 645 cell_1rw
* cell instance $19365 r0 *1 31.02,163.8
X$19365 153 635 154 644 645 cell_1rw
* cell instance $19366 m0 *1 31.02,166.53
X$19366 153 637 154 644 645 cell_1rw
* cell instance $19367 r0 *1 31.02,166.53
X$19367 153 636 154 644 645 cell_1rw
* cell instance $19368 m0 *1 31.02,169.26
X$19368 153 639 154 644 645 cell_1rw
* cell instance $19369 r0 *1 31.02,169.26
X$19369 153 638 154 644 645 cell_1rw
* cell instance $19370 m0 *1 31.02,171.99
X$19370 153 640 154 644 645 cell_1rw
* cell instance $19371 r0 *1 31.02,171.99
X$19371 153 641 154 644 645 cell_1rw
* cell instance $19372 m0 *1 31.02,174.72
X$19372 153 642 154 644 645 cell_1rw
* cell instance $19373 r0 *1 31.02,174.72
X$19373 153 643 154 644 645 cell_1rw
* cell instance $19374 m0 *1 31.725,90.09
X$19374 155 581 156 644 645 cell_1rw
* cell instance $19375 r0 *1 31.725,87.36
X$19375 155 322 156 644 645 cell_1rw
* cell instance $19376 r0 *1 31.725,90.09
X$19376 155 580 156 644 645 cell_1rw
* cell instance $19377 m0 *1 31.725,92.82
X$19377 155 583 156 644 645 cell_1rw
* cell instance $19378 r0 *1 31.725,92.82
X$19378 155 582 156 644 645 cell_1rw
* cell instance $19379 m0 *1 31.725,95.55
X$19379 155 584 156 644 645 cell_1rw
* cell instance $19380 r0 *1 31.725,95.55
X$19380 155 585 156 644 645 cell_1rw
* cell instance $19381 m0 *1 31.725,98.28
X$19381 155 586 156 644 645 cell_1rw
* cell instance $19382 r0 *1 31.725,98.28
X$19382 155 587 156 644 645 cell_1rw
* cell instance $19383 m0 *1 31.725,101.01
X$19383 155 588 156 644 645 cell_1rw
* cell instance $19384 r0 *1 31.725,101.01
X$19384 155 589 156 644 645 cell_1rw
* cell instance $19385 m0 *1 31.725,103.74
X$19385 155 590 156 644 645 cell_1rw
* cell instance $19386 r0 *1 31.725,103.74
X$19386 155 591 156 644 645 cell_1rw
* cell instance $19387 m0 *1 31.725,106.47
X$19387 155 593 156 644 645 cell_1rw
* cell instance $19388 r0 *1 31.725,106.47
X$19388 155 592 156 644 645 cell_1rw
* cell instance $19389 m0 *1 31.725,109.2
X$19389 155 594 156 644 645 cell_1rw
* cell instance $19390 m0 *1 31.725,111.93
X$19390 155 597 156 644 645 cell_1rw
* cell instance $19391 r0 *1 31.725,109.2
X$19391 155 595 156 644 645 cell_1rw
* cell instance $19392 r0 *1 31.725,111.93
X$19392 155 596 156 644 645 cell_1rw
* cell instance $19393 m0 *1 31.725,114.66
X$19393 155 598 156 644 645 cell_1rw
* cell instance $19394 r0 *1 31.725,114.66
X$19394 155 599 156 644 645 cell_1rw
* cell instance $19395 m0 *1 31.725,117.39
X$19395 155 600 156 644 645 cell_1rw
* cell instance $19396 r0 *1 31.725,117.39
X$19396 155 601 156 644 645 cell_1rw
* cell instance $19397 m0 *1 31.725,120.12
X$19397 155 602 156 644 645 cell_1rw
* cell instance $19398 r0 *1 31.725,120.12
X$19398 155 603 156 644 645 cell_1rw
* cell instance $19399 m0 *1 31.725,122.85
X$19399 155 604 156 644 645 cell_1rw
* cell instance $19400 r0 *1 31.725,122.85
X$19400 155 605 156 644 645 cell_1rw
* cell instance $19401 m0 *1 31.725,125.58
X$19401 155 606 156 644 645 cell_1rw
* cell instance $19402 r0 *1 31.725,125.58
X$19402 155 607 156 644 645 cell_1rw
* cell instance $19403 m0 *1 31.725,128.31
X$19403 155 609 156 644 645 cell_1rw
* cell instance $19404 r0 *1 31.725,128.31
X$19404 155 608 156 644 645 cell_1rw
* cell instance $19405 m0 *1 31.725,131.04
X$19405 155 610 156 644 645 cell_1rw
* cell instance $19406 m0 *1 31.725,133.77
X$19406 155 612 156 644 645 cell_1rw
* cell instance $19407 r0 *1 31.725,131.04
X$19407 155 611 156 644 645 cell_1rw
* cell instance $19408 r0 *1 31.725,133.77
X$19408 155 613 156 644 645 cell_1rw
* cell instance $19409 m0 *1 31.725,136.5
X$19409 155 615 156 644 645 cell_1rw
* cell instance $19410 m0 *1 31.725,139.23
X$19410 155 617 156 644 645 cell_1rw
* cell instance $19411 r0 *1 31.725,136.5
X$19411 155 614 156 644 645 cell_1rw
* cell instance $19412 r0 *1 31.725,139.23
X$19412 155 616 156 644 645 cell_1rw
* cell instance $19413 m0 *1 31.725,141.96
X$19413 155 618 156 644 645 cell_1rw
* cell instance $19414 r0 *1 31.725,141.96
X$19414 155 619 156 644 645 cell_1rw
* cell instance $19415 m0 *1 31.725,144.69
X$19415 155 620 156 644 645 cell_1rw
* cell instance $19416 r0 *1 31.725,144.69
X$19416 155 621 156 644 645 cell_1rw
* cell instance $19417 m0 *1 31.725,147.42
X$19417 155 622 156 644 645 cell_1rw
* cell instance $19418 r0 *1 31.725,147.42
X$19418 155 623 156 644 645 cell_1rw
* cell instance $19419 m0 *1 31.725,150.15
X$19419 155 624 156 644 645 cell_1rw
* cell instance $19420 r0 *1 31.725,150.15
X$19420 155 625 156 644 645 cell_1rw
* cell instance $19421 m0 *1 31.725,152.88
X$19421 155 626 156 644 645 cell_1rw
* cell instance $19422 r0 *1 31.725,152.88
X$19422 155 627 156 644 645 cell_1rw
* cell instance $19423 m0 *1 31.725,155.61
X$19423 155 628 156 644 645 cell_1rw
* cell instance $19424 r0 *1 31.725,155.61
X$19424 155 629 156 644 645 cell_1rw
* cell instance $19425 m0 *1 31.725,158.34
X$19425 155 630 156 644 645 cell_1rw
* cell instance $19426 r0 *1 31.725,158.34
X$19426 155 631 156 644 645 cell_1rw
* cell instance $19427 m0 *1 31.725,161.07
X$19427 155 632 156 644 645 cell_1rw
* cell instance $19428 r0 *1 31.725,161.07
X$19428 155 633 156 644 645 cell_1rw
* cell instance $19429 m0 *1 31.725,163.8
X$19429 155 634 156 644 645 cell_1rw
* cell instance $19430 r0 *1 31.725,163.8
X$19430 155 635 156 644 645 cell_1rw
* cell instance $19431 m0 *1 31.725,166.53
X$19431 155 637 156 644 645 cell_1rw
* cell instance $19432 r0 *1 31.725,166.53
X$19432 155 636 156 644 645 cell_1rw
* cell instance $19433 m0 *1 31.725,169.26
X$19433 155 639 156 644 645 cell_1rw
* cell instance $19434 r0 *1 31.725,169.26
X$19434 155 638 156 644 645 cell_1rw
* cell instance $19435 m0 *1 31.725,171.99
X$19435 155 640 156 644 645 cell_1rw
* cell instance $19436 r0 *1 31.725,171.99
X$19436 155 641 156 644 645 cell_1rw
* cell instance $19437 m0 *1 31.725,174.72
X$19437 155 642 156 644 645 cell_1rw
* cell instance $19438 r0 *1 31.725,174.72
X$19438 155 643 156 644 645 cell_1rw
* cell instance $19439 m0 *1 32.43,90.09
X$19439 157 581 158 644 645 cell_1rw
* cell instance $19440 r0 *1 32.43,87.36
X$19440 157 322 158 644 645 cell_1rw
* cell instance $19441 r0 *1 32.43,90.09
X$19441 157 580 158 644 645 cell_1rw
* cell instance $19442 m0 *1 32.43,92.82
X$19442 157 583 158 644 645 cell_1rw
* cell instance $19443 r0 *1 32.43,92.82
X$19443 157 582 158 644 645 cell_1rw
* cell instance $19444 m0 *1 32.43,95.55
X$19444 157 584 158 644 645 cell_1rw
* cell instance $19445 r0 *1 32.43,95.55
X$19445 157 585 158 644 645 cell_1rw
* cell instance $19446 m0 *1 32.43,98.28
X$19446 157 586 158 644 645 cell_1rw
* cell instance $19447 r0 *1 32.43,98.28
X$19447 157 587 158 644 645 cell_1rw
* cell instance $19448 m0 *1 32.43,101.01
X$19448 157 588 158 644 645 cell_1rw
* cell instance $19449 r0 *1 32.43,101.01
X$19449 157 589 158 644 645 cell_1rw
* cell instance $19450 m0 *1 32.43,103.74
X$19450 157 590 158 644 645 cell_1rw
* cell instance $19451 r0 *1 32.43,103.74
X$19451 157 591 158 644 645 cell_1rw
* cell instance $19452 m0 *1 32.43,106.47
X$19452 157 593 158 644 645 cell_1rw
* cell instance $19453 r0 *1 32.43,106.47
X$19453 157 592 158 644 645 cell_1rw
* cell instance $19454 m0 *1 32.43,109.2
X$19454 157 594 158 644 645 cell_1rw
* cell instance $19455 r0 *1 32.43,109.2
X$19455 157 595 158 644 645 cell_1rw
* cell instance $19456 m0 *1 32.43,111.93
X$19456 157 597 158 644 645 cell_1rw
* cell instance $19457 r0 *1 32.43,111.93
X$19457 157 596 158 644 645 cell_1rw
* cell instance $19458 m0 *1 32.43,114.66
X$19458 157 598 158 644 645 cell_1rw
* cell instance $19459 r0 *1 32.43,114.66
X$19459 157 599 158 644 645 cell_1rw
* cell instance $19460 m0 *1 32.43,117.39
X$19460 157 600 158 644 645 cell_1rw
* cell instance $19461 r0 *1 32.43,117.39
X$19461 157 601 158 644 645 cell_1rw
* cell instance $19462 m0 *1 32.43,120.12
X$19462 157 602 158 644 645 cell_1rw
* cell instance $19463 r0 *1 32.43,120.12
X$19463 157 603 158 644 645 cell_1rw
* cell instance $19464 m0 *1 32.43,122.85
X$19464 157 604 158 644 645 cell_1rw
* cell instance $19465 r0 *1 32.43,122.85
X$19465 157 605 158 644 645 cell_1rw
* cell instance $19466 m0 *1 32.43,125.58
X$19466 157 606 158 644 645 cell_1rw
* cell instance $19467 r0 *1 32.43,125.58
X$19467 157 607 158 644 645 cell_1rw
* cell instance $19468 m0 *1 32.43,128.31
X$19468 157 609 158 644 645 cell_1rw
* cell instance $19469 r0 *1 32.43,128.31
X$19469 157 608 158 644 645 cell_1rw
* cell instance $19470 m0 *1 32.43,131.04
X$19470 157 610 158 644 645 cell_1rw
* cell instance $19471 r0 *1 32.43,131.04
X$19471 157 611 158 644 645 cell_1rw
* cell instance $19472 m0 *1 32.43,133.77
X$19472 157 612 158 644 645 cell_1rw
* cell instance $19473 r0 *1 32.43,133.77
X$19473 157 613 158 644 645 cell_1rw
* cell instance $19474 m0 *1 32.43,136.5
X$19474 157 615 158 644 645 cell_1rw
* cell instance $19475 r0 *1 32.43,136.5
X$19475 157 614 158 644 645 cell_1rw
* cell instance $19476 m0 *1 32.43,139.23
X$19476 157 617 158 644 645 cell_1rw
* cell instance $19477 r0 *1 32.43,139.23
X$19477 157 616 158 644 645 cell_1rw
* cell instance $19478 m0 *1 32.43,141.96
X$19478 157 618 158 644 645 cell_1rw
* cell instance $19479 r0 *1 32.43,141.96
X$19479 157 619 158 644 645 cell_1rw
* cell instance $19480 m0 *1 32.43,144.69
X$19480 157 620 158 644 645 cell_1rw
* cell instance $19481 r0 *1 32.43,144.69
X$19481 157 621 158 644 645 cell_1rw
* cell instance $19482 m0 *1 32.43,147.42
X$19482 157 622 158 644 645 cell_1rw
* cell instance $19483 r0 *1 32.43,147.42
X$19483 157 623 158 644 645 cell_1rw
* cell instance $19484 m0 *1 32.43,150.15
X$19484 157 624 158 644 645 cell_1rw
* cell instance $19485 r0 *1 32.43,150.15
X$19485 157 625 158 644 645 cell_1rw
* cell instance $19486 m0 *1 32.43,152.88
X$19486 157 626 158 644 645 cell_1rw
* cell instance $19487 r0 *1 32.43,152.88
X$19487 157 627 158 644 645 cell_1rw
* cell instance $19488 m0 *1 32.43,155.61
X$19488 157 628 158 644 645 cell_1rw
* cell instance $19489 r0 *1 32.43,155.61
X$19489 157 629 158 644 645 cell_1rw
* cell instance $19490 m0 *1 32.43,158.34
X$19490 157 630 158 644 645 cell_1rw
* cell instance $19491 r0 *1 32.43,158.34
X$19491 157 631 158 644 645 cell_1rw
* cell instance $19492 m0 *1 32.43,161.07
X$19492 157 632 158 644 645 cell_1rw
* cell instance $19493 r0 *1 32.43,161.07
X$19493 157 633 158 644 645 cell_1rw
* cell instance $19494 m0 *1 32.43,163.8
X$19494 157 634 158 644 645 cell_1rw
* cell instance $19495 r0 *1 32.43,163.8
X$19495 157 635 158 644 645 cell_1rw
* cell instance $19496 m0 *1 32.43,166.53
X$19496 157 637 158 644 645 cell_1rw
* cell instance $19497 r0 *1 32.43,166.53
X$19497 157 636 158 644 645 cell_1rw
* cell instance $19498 m0 *1 32.43,169.26
X$19498 157 639 158 644 645 cell_1rw
* cell instance $19499 r0 *1 32.43,169.26
X$19499 157 638 158 644 645 cell_1rw
* cell instance $19500 m0 *1 32.43,171.99
X$19500 157 640 158 644 645 cell_1rw
* cell instance $19501 r0 *1 32.43,171.99
X$19501 157 641 158 644 645 cell_1rw
* cell instance $19502 m0 *1 32.43,174.72
X$19502 157 642 158 644 645 cell_1rw
* cell instance $19503 r0 *1 32.43,174.72
X$19503 157 643 158 644 645 cell_1rw
* cell instance $19504 r0 *1 33.135,87.36
X$19504 159 322 160 644 645 cell_1rw
* cell instance $19505 m0 *1 33.135,90.09
X$19505 159 581 160 644 645 cell_1rw
* cell instance $19506 r0 *1 33.135,90.09
X$19506 159 580 160 644 645 cell_1rw
* cell instance $19507 m0 *1 33.135,92.82
X$19507 159 583 160 644 645 cell_1rw
* cell instance $19508 r0 *1 33.135,92.82
X$19508 159 582 160 644 645 cell_1rw
* cell instance $19509 m0 *1 33.135,95.55
X$19509 159 584 160 644 645 cell_1rw
* cell instance $19510 r0 *1 33.135,95.55
X$19510 159 585 160 644 645 cell_1rw
* cell instance $19511 m0 *1 33.135,98.28
X$19511 159 586 160 644 645 cell_1rw
* cell instance $19512 r0 *1 33.135,98.28
X$19512 159 587 160 644 645 cell_1rw
* cell instance $19513 m0 *1 33.135,101.01
X$19513 159 588 160 644 645 cell_1rw
* cell instance $19514 r0 *1 33.135,101.01
X$19514 159 589 160 644 645 cell_1rw
* cell instance $19515 m0 *1 33.135,103.74
X$19515 159 590 160 644 645 cell_1rw
* cell instance $19516 r0 *1 33.135,103.74
X$19516 159 591 160 644 645 cell_1rw
* cell instance $19517 m0 *1 33.135,106.47
X$19517 159 593 160 644 645 cell_1rw
* cell instance $19518 m0 *1 33.135,109.2
X$19518 159 594 160 644 645 cell_1rw
* cell instance $19519 r0 *1 33.135,106.47
X$19519 159 592 160 644 645 cell_1rw
* cell instance $19520 r0 *1 33.135,109.2
X$19520 159 595 160 644 645 cell_1rw
* cell instance $19521 m0 *1 33.135,111.93
X$19521 159 597 160 644 645 cell_1rw
* cell instance $19522 r0 *1 33.135,111.93
X$19522 159 596 160 644 645 cell_1rw
* cell instance $19523 m0 *1 33.135,114.66
X$19523 159 598 160 644 645 cell_1rw
* cell instance $19524 r0 *1 33.135,114.66
X$19524 159 599 160 644 645 cell_1rw
* cell instance $19525 m0 *1 33.135,117.39
X$19525 159 600 160 644 645 cell_1rw
* cell instance $19526 r0 *1 33.135,117.39
X$19526 159 601 160 644 645 cell_1rw
* cell instance $19527 m0 *1 33.135,120.12
X$19527 159 602 160 644 645 cell_1rw
* cell instance $19528 r0 *1 33.135,120.12
X$19528 159 603 160 644 645 cell_1rw
* cell instance $19529 m0 *1 33.135,122.85
X$19529 159 604 160 644 645 cell_1rw
* cell instance $19530 r0 *1 33.135,122.85
X$19530 159 605 160 644 645 cell_1rw
* cell instance $19531 m0 *1 33.135,125.58
X$19531 159 606 160 644 645 cell_1rw
* cell instance $19532 r0 *1 33.135,125.58
X$19532 159 607 160 644 645 cell_1rw
* cell instance $19533 m0 *1 33.135,128.31
X$19533 159 609 160 644 645 cell_1rw
* cell instance $19534 r0 *1 33.135,128.31
X$19534 159 608 160 644 645 cell_1rw
* cell instance $19535 m0 *1 33.135,131.04
X$19535 159 610 160 644 645 cell_1rw
* cell instance $19536 r0 *1 33.135,131.04
X$19536 159 611 160 644 645 cell_1rw
* cell instance $19537 m0 *1 33.135,133.77
X$19537 159 612 160 644 645 cell_1rw
* cell instance $19538 r0 *1 33.135,133.77
X$19538 159 613 160 644 645 cell_1rw
* cell instance $19539 m0 *1 33.135,136.5
X$19539 159 615 160 644 645 cell_1rw
* cell instance $19540 r0 *1 33.135,136.5
X$19540 159 614 160 644 645 cell_1rw
* cell instance $19541 m0 *1 33.135,139.23
X$19541 159 617 160 644 645 cell_1rw
* cell instance $19542 r0 *1 33.135,139.23
X$19542 159 616 160 644 645 cell_1rw
* cell instance $19543 m0 *1 33.135,141.96
X$19543 159 618 160 644 645 cell_1rw
* cell instance $19544 r0 *1 33.135,141.96
X$19544 159 619 160 644 645 cell_1rw
* cell instance $19545 m0 *1 33.135,144.69
X$19545 159 620 160 644 645 cell_1rw
* cell instance $19546 r0 *1 33.135,144.69
X$19546 159 621 160 644 645 cell_1rw
* cell instance $19547 m0 *1 33.135,147.42
X$19547 159 622 160 644 645 cell_1rw
* cell instance $19548 r0 *1 33.135,147.42
X$19548 159 623 160 644 645 cell_1rw
* cell instance $19549 m0 *1 33.135,150.15
X$19549 159 624 160 644 645 cell_1rw
* cell instance $19550 r0 *1 33.135,150.15
X$19550 159 625 160 644 645 cell_1rw
* cell instance $19551 m0 *1 33.135,152.88
X$19551 159 626 160 644 645 cell_1rw
* cell instance $19552 r0 *1 33.135,152.88
X$19552 159 627 160 644 645 cell_1rw
* cell instance $19553 m0 *1 33.135,155.61
X$19553 159 628 160 644 645 cell_1rw
* cell instance $19554 r0 *1 33.135,155.61
X$19554 159 629 160 644 645 cell_1rw
* cell instance $19555 m0 *1 33.135,158.34
X$19555 159 630 160 644 645 cell_1rw
* cell instance $19556 r0 *1 33.135,158.34
X$19556 159 631 160 644 645 cell_1rw
* cell instance $19557 m0 *1 33.135,161.07
X$19557 159 632 160 644 645 cell_1rw
* cell instance $19558 r0 *1 33.135,161.07
X$19558 159 633 160 644 645 cell_1rw
* cell instance $19559 m0 *1 33.135,163.8
X$19559 159 634 160 644 645 cell_1rw
* cell instance $19560 m0 *1 33.135,166.53
X$19560 159 637 160 644 645 cell_1rw
* cell instance $19561 r0 *1 33.135,163.8
X$19561 159 635 160 644 645 cell_1rw
* cell instance $19562 r0 *1 33.135,166.53
X$19562 159 636 160 644 645 cell_1rw
* cell instance $19563 m0 *1 33.135,169.26
X$19563 159 639 160 644 645 cell_1rw
* cell instance $19564 r0 *1 33.135,169.26
X$19564 159 638 160 644 645 cell_1rw
* cell instance $19565 m0 *1 33.135,171.99
X$19565 159 640 160 644 645 cell_1rw
* cell instance $19566 r0 *1 33.135,171.99
X$19566 159 641 160 644 645 cell_1rw
* cell instance $19567 m0 *1 33.135,174.72
X$19567 159 642 160 644 645 cell_1rw
* cell instance $19568 r0 *1 33.135,174.72
X$19568 159 643 160 644 645 cell_1rw
* cell instance $19569 r0 *1 33.84,87.36
X$19569 161 322 162 644 645 cell_1rw
* cell instance $19570 m0 *1 33.84,90.09
X$19570 161 581 162 644 645 cell_1rw
* cell instance $19571 r0 *1 33.84,90.09
X$19571 161 580 162 644 645 cell_1rw
* cell instance $19572 m0 *1 33.84,92.82
X$19572 161 583 162 644 645 cell_1rw
* cell instance $19573 r0 *1 33.84,92.82
X$19573 161 582 162 644 645 cell_1rw
* cell instance $19574 m0 *1 33.84,95.55
X$19574 161 584 162 644 645 cell_1rw
* cell instance $19575 r0 *1 33.84,95.55
X$19575 161 585 162 644 645 cell_1rw
* cell instance $19576 m0 *1 33.84,98.28
X$19576 161 586 162 644 645 cell_1rw
* cell instance $19577 r0 *1 33.84,98.28
X$19577 161 587 162 644 645 cell_1rw
* cell instance $19578 m0 *1 33.84,101.01
X$19578 161 588 162 644 645 cell_1rw
* cell instance $19579 r0 *1 33.84,101.01
X$19579 161 589 162 644 645 cell_1rw
* cell instance $19580 m0 *1 33.84,103.74
X$19580 161 590 162 644 645 cell_1rw
* cell instance $19581 r0 *1 33.84,103.74
X$19581 161 591 162 644 645 cell_1rw
* cell instance $19582 m0 *1 33.84,106.47
X$19582 161 593 162 644 645 cell_1rw
* cell instance $19583 r0 *1 33.84,106.47
X$19583 161 592 162 644 645 cell_1rw
* cell instance $19584 m0 *1 33.84,109.2
X$19584 161 594 162 644 645 cell_1rw
* cell instance $19585 r0 *1 33.84,109.2
X$19585 161 595 162 644 645 cell_1rw
* cell instance $19586 m0 *1 33.84,111.93
X$19586 161 597 162 644 645 cell_1rw
* cell instance $19587 m0 *1 33.84,114.66
X$19587 161 598 162 644 645 cell_1rw
* cell instance $19588 r0 *1 33.84,111.93
X$19588 161 596 162 644 645 cell_1rw
* cell instance $19589 m0 *1 33.84,117.39
X$19589 161 600 162 644 645 cell_1rw
* cell instance $19590 r0 *1 33.84,114.66
X$19590 161 599 162 644 645 cell_1rw
* cell instance $19591 r0 *1 33.84,117.39
X$19591 161 601 162 644 645 cell_1rw
* cell instance $19592 m0 *1 33.84,120.12
X$19592 161 602 162 644 645 cell_1rw
* cell instance $19593 r0 *1 33.84,120.12
X$19593 161 603 162 644 645 cell_1rw
* cell instance $19594 m0 *1 33.84,122.85
X$19594 161 604 162 644 645 cell_1rw
* cell instance $19595 r0 *1 33.84,122.85
X$19595 161 605 162 644 645 cell_1rw
* cell instance $19596 m0 *1 33.84,125.58
X$19596 161 606 162 644 645 cell_1rw
* cell instance $19597 m0 *1 33.84,128.31
X$19597 161 609 162 644 645 cell_1rw
* cell instance $19598 r0 *1 33.84,125.58
X$19598 161 607 162 644 645 cell_1rw
* cell instance $19599 r0 *1 33.84,128.31
X$19599 161 608 162 644 645 cell_1rw
* cell instance $19600 m0 *1 33.84,131.04
X$19600 161 610 162 644 645 cell_1rw
* cell instance $19601 r0 *1 33.84,131.04
X$19601 161 611 162 644 645 cell_1rw
* cell instance $19602 m0 *1 33.84,133.77
X$19602 161 612 162 644 645 cell_1rw
* cell instance $19603 r0 *1 33.84,133.77
X$19603 161 613 162 644 645 cell_1rw
* cell instance $19604 m0 *1 33.84,136.5
X$19604 161 615 162 644 645 cell_1rw
* cell instance $19605 r0 *1 33.84,136.5
X$19605 161 614 162 644 645 cell_1rw
* cell instance $19606 m0 *1 33.84,139.23
X$19606 161 617 162 644 645 cell_1rw
* cell instance $19607 r0 *1 33.84,139.23
X$19607 161 616 162 644 645 cell_1rw
* cell instance $19608 m0 *1 33.84,141.96
X$19608 161 618 162 644 645 cell_1rw
* cell instance $19609 r0 *1 33.84,141.96
X$19609 161 619 162 644 645 cell_1rw
* cell instance $19610 m0 *1 33.84,144.69
X$19610 161 620 162 644 645 cell_1rw
* cell instance $19611 r0 *1 33.84,144.69
X$19611 161 621 162 644 645 cell_1rw
* cell instance $19612 m0 *1 33.84,147.42
X$19612 161 622 162 644 645 cell_1rw
* cell instance $19613 m0 *1 33.84,150.15
X$19613 161 624 162 644 645 cell_1rw
* cell instance $19614 r0 *1 33.84,147.42
X$19614 161 623 162 644 645 cell_1rw
* cell instance $19615 r0 *1 33.84,150.15
X$19615 161 625 162 644 645 cell_1rw
* cell instance $19616 m0 *1 33.84,152.88
X$19616 161 626 162 644 645 cell_1rw
* cell instance $19617 r0 *1 33.84,152.88
X$19617 161 627 162 644 645 cell_1rw
* cell instance $19618 m0 *1 33.84,155.61
X$19618 161 628 162 644 645 cell_1rw
* cell instance $19619 m0 *1 33.84,158.34
X$19619 161 630 162 644 645 cell_1rw
* cell instance $19620 r0 *1 33.84,155.61
X$19620 161 629 162 644 645 cell_1rw
* cell instance $19621 r0 *1 33.84,158.34
X$19621 161 631 162 644 645 cell_1rw
* cell instance $19622 m0 *1 33.84,161.07
X$19622 161 632 162 644 645 cell_1rw
* cell instance $19623 r0 *1 33.84,161.07
X$19623 161 633 162 644 645 cell_1rw
* cell instance $19624 m0 *1 33.84,163.8
X$19624 161 634 162 644 645 cell_1rw
* cell instance $19625 m0 *1 33.84,166.53
X$19625 161 637 162 644 645 cell_1rw
* cell instance $19626 r0 *1 33.84,163.8
X$19626 161 635 162 644 645 cell_1rw
* cell instance $19627 r0 *1 33.84,166.53
X$19627 161 636 162 644 645 cell_1rw
* cell instance $19628 m0 *1 33.84,169.26
X$19628 161 639 162 644 645 cell_1rw
* cell instance $19629 r0 *1 33.84,169.26
X$19629 161 638 162 644 645 cell_1rw
* cell instance $19630 m0 *1 33.84,171.99
X$19630 161 640 162 644 645 cell_1rw
* cell instance $19631 m0 *1 33.84,174.72
X$19631 161 642 162 644 645 cell_1rw
* cell instance $19632 r0 *1 33.84,171.99
X$19632 161 641 162 644 645 cell_1rw
* cell instance $19633 r0 *1 33.84,174.72
X$19633 161 643 162 644 645 cell_1rw
* cell instance $19634 r0 *1 34.545,87.36
X$19634 163 322 164 644 645 cell_1rw
* cell instance $19635 m0 *1 34.545,90.09
X$19635 163 581 164 644 645 cell_1rw
* cell instance $19636 r0 *1 34.545,90.09
X$19636 163 580 164 644 645 cell_1rw
* cell instance $19637 m0 *1 34.545,92.82
X$19637 163 583 164 644 645 cell_1rw
* cell instance $19638 r0 *1 34.545,92.82
X$19638 163 582 164 644 645 cell_1rw
* cell instance $19639 m0 *1 34.545,95.55
X$19639 163 584 164 644 645 cell_1rw
* cell instance $19640 r0 *1 34.545,95.55
X$19640 163 585 164 644 645 cell_1rw
* cell instance $19641 m0 *1 34.545,98.28
X$19641 163 586 164 644 645 cell_1rw
* cell instance $19642 r0 *1 34.545,98.28
X$19642 163 587 164 644 645 cell_1rw
* cell instance $19643 m0 *1 34.545,101.01
X$19643 163 588 164 644 645 cell_1rw
* cell instance $19644 r0 *1 34.545,101.01
X$19644 163 589 164 644 645 cell_1rw
* cell instance $19645 m0 *1 34.545,103.74
X$19645 163 590 164 644 645 cell_1rw
* cell instance $19646 m0 *1 34.545,106.47
X$19646 163 593 164 644 645 cell_1rw
* cell instance $19647 r0 *1 34.545,103.74
X$19647 163 591 164 644 645 cell_1rw
* cell instance $19648 r0 *1 34.545,106.47
X$19648 163 592 164 644 645 cell_1rw
* cell instance $19649 m0 *1 34.545,109.2
X$19649 163 594 164 644 645 cell_1rw
* cell instance $19650 r0 *1 34.545,109.2
X$19650 163 595 164 644 645 cell_1rw
* cell instance $19651 m0 *1 34.545,111.93
X$19651 163 597 164 644 645 cell_1rw
* cell instance $19652 r0 *1 34.545,111.93
X$19652 163 596 164 644 645 cell_1rw
* cell instance $19653 m0 *1 34.545,114.66
X$19653 163 598 164 644 645 cell_1rw
* cell instance $19654 r0 *1 34.545,114.66
X$19654 163 599 164 644 645 cell_1rw
* cell instance $19655 m0 *1 34.545,117.39
X$19655 163 600 164 644 645 cell_1rw
* cell instance $19656 r0 *1 34.545,117.39
X$19656 163 601 164 644 645 cell_1rw
* cell instance $19657 m0 *1 34.545,120.12
X$19657 163 602 164 644 645 cell_1rw
* cell instance $19658 m0 *1 34.545,122.85
X$19658 163 604 164 644 645 cell_1rw
* cell instance $19659 r0 *1 34.545,120.12
X$19659 163 603 164 644 645 cell_1rw
* cell instance $19660 r0 *1 34.545,122.85
X$19660 163 605 164 644 645 cell_1rw
* cell instance $19661 m0 *1 34.545,125.58
X$19661 163 606 164 644 645 cell_1rw
* cell instance $19662 m0 *1 34.545,128.31
X$19662 163 609 164 644 645 cell_1rw
* cell instance $19663 r0 *1 34.545,125.58
X$19663 163 607 164 644 645 cell_1rw
* cell instance $19664 r0 *1 34.545,128.31
X$19664 163 608 164 644 645 cell_1rw
* cell instance $19665 m0 *1 34.545,131.04
X$19665 163 610 164 644 645 cell_1rw
* cell instance $19666 r0 *1 34.545,131.04
X$19666 163 611 164 644 645 cell_1rw
* cell instance $19667 m0 *1 34.545,133.77
X$19667 163 612 164 644 645 cell_1rw
* cell instance $19668 r0 *1 34.545,133.77
X$19668 163 613 164 644 645 cell_1rw
* cell instance $19669 m0 *1 34.545,136.5
X$19669 163 615 164 644 645 cell_1rw
* cell instance $19670 r0 *1 34.545,136.5
X$19670 163 614 164 644 645 cell_1rw
* cell instance $19671 m0 *1 34.545,139.23
X$19671 163 617 164 644 645 cell_1rw
* cell instance $19672 r0 *1 34.545,139.23
X$19672 163 616 164 644 645 cell_1rw
* cell instance $19673 m0 *1 34.545,141.96
X$19673 163 618 164 644 645 cell_1rw
* cell instance $19674 r0 *1 34.545,141.96
X$19674 163 619 164 644 645 cell_1rw
* cell instance $19675 m0 *1 34.545,144.69
X$19675 163 620 164 644 645 cell_1rw
* cell instance $19676 r0 *1 34.545,144.69
X$19676 163 621 164 644 645 cell_1rw
* cell instance $19677 m0 *1 34.545,147.42
X$19677 163 622 164 644 645 cell_1rw
* cell instance $19678 r0 *1 34.545,147.42
X$19678 163 623 164 644 645 cell_1rw
* cell instance $19679 m0 *1 34.545,150.15
X$19679 163 624 164 644 645 cell_1rw
* cell instance $19680 r0 *1 34.545,150.15
X$19680 163 625 164 644 645 cell_1rw
* cell instance $19681 m0 *1 34.545,152.88
X$19681 163 626 164 644 645 cell_1rw
* cell instance $19682 r0 *1 34.545,152.88
X$19682 163 627 164 644 645 cell_1rw
* cell instance $19683 m0 *1 34.545,155.61
X$19683 163 628 164 644 645 cell_1rw
* cell instance $19684 m0 *1 34.545,158.34
X$19684 163 630 164 644 645 cell_1rw
* cell instance $19685 r0 *1 34.545,155.61
X$19685 163 629 164 644 645 cell_1rw
* cell instance $19686 r0 *1 34.545,158.34
X$19686 163 631 164 644 645 cell_1rw
* cell instance $19687 m0 *1 34.545,161.07
X$19687 163 632 164 644 645 cell_1rw
* cell instance $19688 r0 *1 34.545,161.07
X$19688 163 633 164 644 645 cell_1rw
* cell instance $19689 m0 *1 34.545,163.8
X$19689 163 634 164 644 645 cell_1rw
* cell instance $19690 r0 *1 34.545,163.8
X$19690 163 635 164 644 645 cell_1rw
* cell instance $19691 m0 *1 34.545,166.53
X$19691 163 637 164 644 645 cell_1rw
* cell instance $19692 m0 *1 34.545,169.26
X$19692 163 639 164 644 645 cell_1rw
* cell instance $19693 r0 *1 34.545,166.53
X$19693 163 636 164 644 645 cell_1rw
* cell instance $19694 r0 *1 34.545,169.26
X$19694 163 638 164 644 645 cell_1rw
* cell instance $19695 m0 *1 34.545,171.99
X$19695 163 640 164 644 645 cell_1rw
* cell instance $19696 r0 *1 34.545,171.99
X$19696 163 641 164 644 645 cell_1rw
* cell instance $19697 m0 *1 34.545,174.72
X$19697 163 642 164 644 645 cell_1rw
* cell instance $19698 r0 *1 34.545,174.72
X$19698 163 643 164 644 645 cell_1rw
* cell instance $19699 m0 *1 35.25,90.09
X$19699 165 581 166 644 645 cell_1rw
* cell instance $19700 r0 *1 35.25,87.36
X$19700 165 322 166 644 645 cell_1rw
* cell instance $19701 m0 *1 35.25,92.82
X$19701 165 583 166 644 645 cell_1rw
* cell instance $19702 r0 *1 35.25,90.09
X$19702 165 580 166 644 645 cell_1rw
* cell instance $19703 r0 *1 35.25,92.82
X$19703 165 582 166 644 645 cell_1rw
* cell instance $19704 m0 *1 35.25,95.55
X$19704 165 584 166 644 645 cell_1rw
* cell instance $19705 r0 *1 35.25,95.55
X$19705 165 585 166 644 645 cell_1rw
* cell instance $19706 m0 *1 35.25,98.28
X$19706 165 586 166 644 645 cell_1rw
* cell instance $19707 r0 *1 35.25,98.28
X$19707 165 587 166 644 645 cell_1rw
* cell instance $19708 m0 *1 35.25,101.01
X$19708 165 588 166 644 645 cell_1rw
* cell instance $19709 r0 *1 35.25,101.01
X$19709 165 589 166 644 645 cell_1rw
* cell instance $19710 m0 *1 35.25,103.74
X$19710 165 590 166 644 645 cell_1rw
* cell instance $19711 r0 *1 35.25,103.74
X$19711 165 591 166 644 645 cell_1rw
* cell instance $19712 m0 *1 35.25,106.47
X$19712 165 593 166 644 645 cell_1rw
* cell instance $19713 r0 *1 35.25,106.47
X$19713 165 592 166 644 645 cell_1rw
* cell instance $19714 m0 *1 35.25,109.2
X$19714 165 594 166 644 645 cell_1rw
* cell instance $19715 m0 *1 35.25,111.93
X$19715 165 597 166 644 645 cell_1rw
* cell instance $19716 r0 *1 35.25,109.2
X$19716 165 595 166 644 645 cell_1rw
* cell instance $19717 r0 *1 35.25,111.93
X$19717 165 596 166 644 645 cell_1rw
* cell instance $19718 m0 *1 35.25,114.66
X$19718 165 598 166 644 645 cell_1rw
* cell instance $19719 r0 *1 35.25,114.66
X$19719 165 599 166 644 645 cell_1rw
* cell instance $19720 m0 *1 35.25,117.39
X$19720 165 600 166 644 645 cell_1rw
* cell instance $19721 r0 *1 35.25,117.39
X$19721 165 601 166 644 645 cell_1rw
* cell instance $19722 m0 *1 35.25,120.12
X$19722 165 602 166 644 645 cell_1rw
* cell instance $19723 r0 *1 35.25,120.12
X$19723 165 603 166 644 645 cell_1rw
* cell instance $19724 m0 *1 35.25,122.85
X$19724 165 604 166 644 645 cell_1rw
* cell instance $19725 m0 *1 35.25,125.58
X$19725 165 606 166 644 645 cell_1rw
* cell instance $19726 r0 *1 35.25,122.85
X$19726 165 605 166 644 645 cell_1rw
* cell instance $19727 r0 *1 35.25,125.58
X$19727 165 607 166 644 645 cell_1rw
* cell instance $19728 m0 *1 35.25,128.31
X$19728 165 609 166 644 645 cell_1rw
* cell instance $19729 r0 *1 35.25,128.31
X$19729 165 608 166 644 645 cell_1rw
* cell instance $19730 m0 *1 35.25,131.04
X$19730 165 610 166 644 645 cell_1rw
* cell instance $19731 r0 *1 35.25,131.04
X$19731 165 611 166 644 645 cell_1rw
* cell instance $19732 m0 *1 35.25,133.77
X$19732 165 612 166 644 645 cell_1rw
* cell instance $19733 r0 *1 35.25,133.77
X$19733 165 613 166 644 645 cell_1rw
* cell instance $19734 m0 *1 35.25,136.5
X$19734 165 615 166 644 645 cell_1rw
* cell instance $19735 r0 *1 35.25,136.5
X$19735 165 614 166 644 645 cell_1rw
* cell instance $19736 m0 *1 35.25,139.23
X$19736 165 617 166 644 645 cell_1rw
* cell instance $19737 r0 *1 35.25,139.23
X$19737 165 616 166 644 645 cell_1rw
* cell instance $19738 m0 *1 35.25,141.96
X$19738 165 618 166 644 645 cell_1rw
* cell instance $19739 r0 *1 35.25,141.96
X$19739 165 619 166 644 645 cell_1rw
* cell instance $19740 m0 *1 35.25,144.69
X$19740 165 620 166 644 645 cell_1rw
* cell instance $19741 r0 *1 35.25,144.69
X$19741 165 621 166 644 645 cell_1rw
* cell instance $19742 m0 *1 35.25,147.42
X$19742 165 622 166 644 645 cell_1rw
* cell instance $19743 r0 *1 35.25,147.42
X$19743 165 623 166 644 645 cell_1rw
* cell instance $19744 m0 *1 35.25,150.15
X$19744 165 624 166 644 645 cell_1rw
* cell instance $19745 r0 *1 35.25,150.15
X$19745 165 625 166 644 645 cell_1rw
* cell instance $19746 m0 *1 35.25,152.88
X$19746 165 626 166 644 645 cell_1rw
* cell instance $19747 m0 *1 35.25,155.61
X$19747 165 628 166 644 645 cell_1rw
* cell instance $19748 r0 *1 35.25,152.88
X$19748 165 627 166 644 645 cell_1rw
* cell instance $19749 r0 *1 35.25,155.61
X$19749 165 629 166 644 645 cell_1rw
* cell instance $19750 m0 *1 35.25,158.34
X$19750 165 630 166 644 645 cell_1rw
* cell instance $19751 r0 *1 35.25,158.34
X$19751 165 631 166 644 645 cell_1rw
* cell instance $19752 m0 *1 35.25,161.07
X$19752 165 632 166 644 645 cell_1rw
* cell instance $19753 r0 *1 35.25,161.07
X$19753 165 633 166 644 645 cell_1rw
* cell instance $19754 m0 *1 35.25,163.8
X$19754 165 634 166 644 645 cell_1rw
* cell instance $19755 m0 *1 35.25,166.53
X$19755 165 637 166 644 645 cell_1rw
* cell instance $19756 r0 *1 35.25,163.8
X$19756 165 635 166 644 645 cell_1rw
* cell instance $19757 r0 *1 35.25,166.53
X$19757 165 636 166 644 645 cell_1rw
* cell instance $19758 m0 *1 35.25,169.26
X$19758 165 639 166 644 645 cell_1rw
* cell instance $19759 r0 *1 35.25,169.26
X$19759 165 638 166 644 645 cell_1rw
* cell instance $19760 m0 *1 35.25,171.99
X$19760 165 640 166 644 645 cell_1rw
* cell instance $19761 r0 *1 35.25,171.99
X$19761 165 641 166 644 645 cell_1rw
* cell instance $19762 m0 *1 35.25,174.72
X$19762 165 642 166 644 645 cell_1rw
* cell instance $19763 r0 *1 35.25,174.72
X$19763 165 643 166 644 645 cell_1rw
* cell instance $19764 m0 *1 35.955,90.09
X$19764 167 581 168 644 645 cell_1rw
* cell instance $19765 r0 *1 35.955,87.36
X$19765 167 322 168 644 645 cell_1rw
* cell instance $19766 r0 *1 35.955,90.09
X$19766 167 580 168 644 645 cell_1rw
* cell instance $19767 m0 *1 35.955,92.82
X$19767 167 583 168 644 645 cell_1rw
* cell instance $19768 r0 *1 35.955,92.82
X$19768 167 582 168 644 645 cell_1rw
* cell instance $19769 m0 *1 35.955,95.55
X$19769 167 584 168 644 645 cell_1rw
* cell instance $19770 r0 *1 35.955,95.55
X$19770 167 585 168 644 645 cell_1rw
* cell instance $19771 m0 *1 35.955,98.28
X$19771 167 586 168 644 645 cell_1rw
* cell instance $19772 r0 *1 35.955,98.28
X$19772 167 587 168 644 645 cell_1rw
* cell instance $19773 m0 *1 35.955,101.01
X$19773 167 588 168 644 645 cell_1rw
* cell instance $19774 r0 *1 35.955,101.01
X$19774 167 589 168 644 645 cell_1rw
* cell instance $19775 m0 *1 35.955,103.74
X$19775 167 590 168 644 645 cell_1rw
* cell instance $19776 m0 *1 35.955,106.47
X$19776 167 593 168 644 645 cell_1rw
* cell instance $19777 r0 *1 35.955,103.74
X$19777 167 591 168 644 645 cell_1rw
* cell instance $19778 r0 *1 35.955,106.47
X$19778 167 592 168 644 645 cell_1rw
* cell instance $19779 m0 *1 35.955,109.2
X$19779 167 594 168 644 645 cell_1rw
* cell instance $19780 r0 *1 35.955,109.2
X$19780 167 595 168 644 645 cell_1rw
* cell instance $19781 m0 *1 35.955,111.93
X$19781 167 597 168 644 645 cell_1rw
* cell instance $19782 r0 *1 35.955,111.93
X$19782 167 596 168 644 645 cell_1rw
* cell instance $19783 m0 *1 35.955,114.66
X$19783 167 598 168 644 645 cell_1rw
* cell instance $19784 m0 *1 35.955,117.39
X$19784 167 600 168 644 645 cell_1rw
* cell instance $19785 r0 *1 35.955,114.66
X$19785 167 599 168 644 645 cell_1rw
* cell instance $19786 r0 *1 35.955,117.39
X$19786 167 601 168 644 645 cell_1rw
* cell instance $19787 m0 *1 35.955,120.12
X$19787 167 602 168 644 645 cell_1rw
* cell instance $19788 r0 *1 35.955,120.12
X$19788 167 603 168 644 645 cell_1rw
* cell instance $19789 m0 *1 35.955,122.85
X$19789 167 604 168 644 645 cell_1rw
* cell instance $19790 r0 *1 35.955,122.85
X$19790 167 605 168 644 645 cell_1rw
* cell instance $19791 m0 *1 35.955,125.58
X$19791 167 606 168 644 645 cell_1rw
* cell instance $19792 r0 *1 35.955,125.58
X$19792 167 607 168 644 645 cell_1rw
* cell instance $19793 m0 *1 35.955,128.31
X$19793 167 609 168 644 645 cell_1rw
* cell instance $19794 r0 *1 35.955,128.31
X$19794 167 608 168 644 645 cell_1rw
* cell instance $19795 m0 *1 35.955,131.04
X$19795 167 610 168 644 645 cell_1rw
* cell instance $19796 r0 *1 35.955,131.04
X$19796 167 611 168 644 645 cell_1rw
* cell instance $19797 m0 *1 35.955,133.77
X$19797 167 612 168 644 645 cell_1rw
* cell instance $19798 r0 *1 35.955,133.77
X$19798 167 613 168 644 645 cell_1rw
* cell instance $19799 m0 *1 35.955,136.5
X$19799 167 615 168 644 645 cell_1rw
* cell instance $19800 r0 *1 35.955,136.5
X$19800 167 614 168 644 645 cell_1rw
* cell instance $19801 m0 *1 35.955,139.23
X$19801 167 617 168 644 645 cell_1rw
* cell instance $19802 r0 *1 35.955,139.23
X$19802 167 616 168 644 645 cell_1rw
* cell instance $19803 m0 *1 35.955,141.96
X$19803 167 618 168 644 645 cell_1rw
* cell instance $19804 r0 *1 35.955,141.96
X$19804 167 619 168 644 645 cell_1rw
* cell instance $19805 m0 *1 35.955,144.69
X$19805 167 620 168 644 645 cell_1rw
* cell instance $19806 r0 *1 35.955,144.69
X$19806 167 621 168 644 645 cell_1rw
* cell instance $19807 m0 *1 35.955,147.42
X$19807 167 622 168 644 645 cell_1rw
* cell instance $19808 r0 *1 35.955,147.42
X$19808 167 623 168 644 645 cell_1rw
* cell instance $19809 m0 *1 35.955,150.15
X$19809 167 624 168 644 645 cell_1rw
* cell instance $19810 r0 *1 35.955,150.15
X$19810 167 625 168 644 645 cell_1rw
* cell instance $19811 m0 *1 35.955,152.88
X$19811 167 626 168 644 645 cell_1rw
* cell instance $19812 r0 *1 35.955,152.88
X$19812 167 627 168 644 645 cell_1rw
* cell instance $19813 m0 *1 35.955,155.61
X$19813 167 628 168 644 645 cell_1rw
* cell instance $19814 m0 *1 35.955,158.34
X$19814 167 630 168 644 645 cell_1rw
* cell instance $19815 r0 *1 35.955,155.61
X$19815 167 629 168 644 645 cell_1rw
* cell instance $19816 r0 *1 35.955,158.34
X$19816 167 631 168 644 645 cell_1rw
* cell instance $19817 m0 *1 35.955,161.07
X$19817 167 632 168 644 645 cell_1rw
* cell instance $19818 r0 *1 35.955,161.07
X$19818 167 633 168 644 645 cell_1rw
* cell instance $19819 m0 *1 35.955,163.8
X$19819 167 634 168 644 645 cell_1rw
* cell instance $19820 r0 *1 35.955,163.8
X$19820 167 635 168 644 645 cell_1rw
* cell instance $19821 m0 *1 35.955,166.53
X$19821 167 637 168 644 645 cell_1rw
* cell instance $19822 r0 *1 35.955,166.53
X$19822 167 636 168 644 645 cell_1rw
* cell instance $19823 m0 *1 35.955,169.26
X$19823 167 639 168 644 645 cell_1rw
* cell instance $19824 r0 *1 35.955,169.26
X$19824 167 638 168 644 645 cell_1rw
* cell instance $19825 m0 *1 35.955,171.99
X$19825 167 640 168 644 645 cell_1rw
* cell instance $19826 r0 *1 35.955,171.99
X$19826 167 641 168 644 645 cell_1rw
* cell instance $19827 m0 *1 35.955,174.72
X$19827 167 642 168 644 645 cell_1rw
* cell instance $19828 r0 *1 35.955,174.72
X$19828 167 643 168 644 645 cell_1rw
* cell instance $19829 m0 *1 36.66,90.09
X$19829 169 581 170 644 645 cell_1rw
* cell instance $19830 r0 *1 36.66,87.36
X$19830 169 322 170 644 645 cell_1rw
* cell instance $19831 r0 *1 36.66,90.09
X$19831 169 580 170 644 645 cell_1rw
* cell instance $19832 m0 *1 36.66,92.82
X$19832 169 583 170 644 645 cell_1rw
* cell instance $19833 m0 *1 36.66,95.55
X$19833 169 584 170 644 645 cell_1rw
* cell instance $19834 r0 *1 36.66,92.82
X$19834 169 582 170 644 645 cell_1rw
* cell instance $19835 r0 *1 36.66,95.55
X$19835 169 585 170 644 645 cell_1rw
* cell instance $19836 m0 *1 36.66,98.28
X$19836 169 586 170 644 645 cell_1rw
* cell instance $19837 m0 *1 36.66,101.01
X$19837 169 588 170 644 645 cell_1rw
* cell instance $19838 r0 *1 36.66,98.28
X$19838 169 587 170 644 645 cell_1rw
* cell instance $19839 r0 *1 36.66,101.01
X$19839 169 589 170 644 645 cell_1rw
* cell instance $19840 m0 *1 36.66,103.74
X$19840 169 590 170 644 645 cell_1rw
* cell instance $19841 r0 *1 36.66,103.74
X$19841 169 591 170 644 645 cell_1rw
* cell instance $19842 m0 *1 36.66,106.47
X$19842 169 593 170 644 645 cell_1rw
* cell instance $19843 r0 *1 36.66,106.47
X$19843 169 592 170 644 645 cell_1rw
* cell instance $19844 m0 *1 36.66,109.2
X$19844 169 594 170 644 645 cell_1rw
* cell instance $19845 r0 *1 36.66,109.2
X$19845 169 595 170 644 645 cell_1rw
* cell instance $19846 m0 *1 36.66,111.93
X$19846 169 597 170 644 645 cell_1rw
* cell instance $19847 r0 *1 36.66,111.93
X$19847 169 596 170 644 645 cell_1rw
* cell instance $19848 m0 *1 36.66,114.66
X$19848 169 598 170 644 645 cell_1rw
* cell instance $19849 r0 *1 36.66,114.66
X$19849 169 599 170 644 645 cell_1rw
* cell instance $19850 m0 *1 36.66,117.39
X$19850 169 600 170 644 645 cell_1rw
* cell instance $19851 r0 *1 36.66,117.39
X$19851 169 601 170 644 645 cell_1rw
* cell instance $19852 m0 *1 36.66,120.12
X$19852 169 602 170 644 645 cell_1rw
* cell instance $19853 m0 *1 36.66,122.85
X$19853 169 604 170 644 645 cell_1rw
* cell instance $19854 r0 *1 36.66,120.12
X$19854 169 603 170 644 645 cell_1rw
* cell instance $19855 r0 *1 36.66,122.85
X$19855 169 605 170 644 645 cell_1rw
* cell instance $19856 m0 *1 36.66,125.58
X$19856 169 606 170 644 645 cell_1rw
* cell instance $19857 m0 *1 36.66,128.31
X$19857 169 609 170 644 645 cell_1rw
* cell instance $19858 r0 *1 36.66,125.58
X$19858 169 607 170 644 645 cell_1rw
* cell instance $19859 r0 *1 36.66,128.31
X$19859 169 608 170 644 645 cell_1rw
* cell instance $19860 m0 *1 36.66,131.04
X$19860 169 610 170 644 645 cell_1rw
* cell instance $19861 m0 *1 36.66,133.77
X$19861 169 612 170 644 645 cell_1rw
* cell instance $19862 r0 *1 36.66,131.04
X$19862 169 611 170 644 645 cell_1rw
* cell instance $19863 r0 *1 36.66,133.77
X$19863 169 613 170 644 645 cell_1rw
* cell instance $19864 m0 *1 36.66,136.5
X$19864 169 615 170 644 645 cell_1rw
* cell instance $19865 r0 *1 36.66,136.5
X$19865 169 614 170 644 645 cell_1rw
* cell instance $19866 m0 *1 36.66,139.23
X$19866 169 617 170 644 645 cell_1rw
* cell instance $19867 r0 *1 36.66,139.23
X$19867 169 616 170 644 645 cell_1rw
* cell instance $19868 m0 *1 36.66,141.96
X$19868 169 618 170 644 645 cell_1rw
* cell instance $19869 r0 *1 36.66,141.96
X$19869 169 619 170 644 645 cell_1rw
* cell instance $19870 m0 *1 36.66,144.69
X$19870 169 620 170 644 645 cell_1rw
* cell instance $19871 r0 *1 36.66,144.69
X$19871 169 621 170 644 645 cell_1rw
* cell instance $19872 m0 *1 36.66,147.42
X$19872 169 622 170 644 645 cell_1rw
* cell instance $19873 r0 *1 36.66,147.42
X$19873 169 623 170 644 645 cell_1rw
* cell instance $19874 m0 *1 36.66,150.15
X$19874 169 624 170 644 645 cell_1rw
* cell instance $19875 r0 *1 36.66,150.15
X$19875 169 625 170 644 645 cell_1rw
* cell instance $19876 m0 *1 36.66,152.88
X$19876 169 626 170 644 645 cell_1rw
* cell instance $19877 r0 *1 36.66,152.88
X$19877 169 627 170 644 645 cell_1rw
* cell instance $19878 m0 *1 36.66,155.61
X$19878 169 628 170 644 645 cell_1rw
* cell instance $19879 r0 *1 36.66,155.61
X$19879 169 629 170 644 645 cell_1rw
* cell instance $19880 m0 *1 36.66,158.34
X$19880 169 630 170 644 645 cell_1rw
* cell instance $19881 r0 *1 36.66,158.34
X$19881 169 631 170 644 645 cell_1rw
* cell instance $19882 m0 *1 36.66,161.07
X$19882 169 632 170 644 645 cell_1rw
* cell instance $19883 r0 *1 36.66,161.07
X$19883 169 633 170 644 645 cell_1rw
* cell instance $19884 m0 *1 36.66,163.8
X$19884 169 634 170 644 645 cell_1rw
* cell instance $19885 r0 *1 36.66,163.8
X$19885 169 635 170 644 645 cell_1rw
* cell instance $19886 m0 *1 36.66,166.53
X$19886 169 637 170 644 645 cell_1rw
* cell instance $19887 r0 *1 36.66,166.53
X$19887 169 636 170 644 645 cell_1rw
* cell instance $19888 m0 *1 36.66,169.26
X$19888 169 639 170 644 645 cell_1rw
* cell instance $19889 r0 *1 36.66,169.26
X$19889 169 638 170 644 645 cell_1rw
* cell instance $19890 m0 *1 36.66,171.99
X$19890 169 640 170 644 645 cell_1rw
* cell instance $19891 r0 *1 36.66,171.99
X$19891 169 641 170 644 645 cell_1rw
* cell instance $19892 m0 *1 36.66,174.72
X$19892 169 642 170 644 645 cell_1rw
* cell instance $19893 r0 *1 36.66,174.72
X$19893 169 643 170 644 645 cell_1rw
* cell instance $19894 m0 *1 37.365,90.09
X$19894 171 581 172 644 645 cell_1rw
* cell instance $19895 r0 *1 37.365,87.36
X$19895 171 322 172 644 645 cell_1rw
* cell instance $19896 r0 *1 37.365,90.09
X$19896 171 580 172 644 645 cell_1rw
* cell instance $19897 m0 *1 37.365,92.82
X$19897 171 583 172 644 645 cell_1rw
* cell instance $19898 r0 *1 37.365,92.82
X$19898 171 582 172 644 645 cell_1rw
* cell instance $19899 m0 *1 37.365,95.55
X$19899 171 584 172 644 645 cell_1rw
* cell instance $19900 r0 *1 37.365,95.55
X$19900 171 585 172 644 645 cell_1rw
* cell instance $19901 m0 *1 37.365,98.28
X$19901 171 586 172 644 645 cell_1rw
* cell instance $19902 m0 *1 37.365,101.01
X$19902 171 588 172 644 645 cell_1rw
* cell instance $19903 r0 *1 37.365,98.28
X$19903 171 587 172 644 645 cell_1rw
* cell instance $19904 r0 *1 37.365,101.01
X$19904 171 589 172 644 645 cell_1rw
* cell instance $19905 m0 *1 37.365,103.74
X$19905 171 590 172 644 645 cell_1rw
* cell instance $19906 r0 *1 37.365,103.74
X$19906 171 591 172 644 645 cell_1rw
* cell instance $19907 m0 *1 37.365,106.47
X$19907 171 593 172 644 645 cell_1rw
* cell instance $19908 r0 *1 37.365,106.47
X$19908 171 592 172 644 645 cell_1rw
* cell instance $19909 m0 *1 37.365,109.2
X$19909 171 594 172 644 645 cell_1rw
* cell instance $19910 r0 *1 37.365,109.2
X$19910 171 595 172 644 645 cell_1rw
* cell instance $19911 m0 *1 37.365,111.93
X$19911 171 597 172 644 645 cell_1rw
* cell instance $19912 r0 *1 37.365,111.93
X$19912 171 596 172 644 645 cell_1rw
* cell instance $19913 m0 *1 37.365,114.66
X$19913 171 598 172 644 645 cell_1rw
* cell instance $19914 r0 *1 37.365,114.66
X$19914 171 599 172 644 645 cell_1rw
* cell instance $19915 m0 *1 37.365,117.39
X$19915 171 600 172 644 645 cell_1rw
* cell instance $19916 r0 *1 37.365,117.39
X$19916 171 601 172 644 645 cell_1rw
* cell instance $19917 m0 *1 37.365,120.12
X$19917 171 602 172 644 645 cell_1rw
* cell instance $19918 m0 *1 37.365,122.85
X$19918 171 604 172 644 645 cell_1rw
* cell instance $19919 r0 *1 37.365,120.12
X$19919 171 603 172 644 645 cell_1rw
* cell instance $19920 m0 *1 37.365,125.58
X$19920 171 606 172 644 645 cell_1rw
* cell instance $19921 r0 *1 37.365,122.85
X$19921 171 605 172 644 645 cell_1rw
* cell instance $19922 r0 *1 37.365,125.58
X$19922 171 607 172 644 645 cell_1rw
* cell instance $19923 m0 *1 37.365,128.31
X$19923 171 609 172 644 645 cell_1rw
* cell instance $19924 r0 *1 37.365,128.31
X$19924 171 608 172 644 645 cell_1rw
* cell instance $19925 m0 *1 37.365,131.04
X$19925 171 610 172 644 645 cell_1rw
* cell instance $19926 m0 *1 37.365,133.77
X$19926 171 612 172 644 645 cell_1rw
* cell instance $19927 r0 *1 37.365,131.04
X$19927 171 611 172 644 645 cell_1rw
* cell instance $19928 r0 *1 37.365,133.77
X$19928 171 613 172 644 645 cell_1rw
* cell instance $19929 m0 *1 37.365,136.5
X$19929 171 615 172 644 645 cell_1rw
* cell instance $19930 r0 *1 37.365,136.5
X$19930 171 614 172 644 645 cell_1rw
* cell instance $19931 m0 *1 37.365,139.23
X$19931 171 617 172 644 645 cell_1rw
* cell instance $19932 r0 *1 37.365,139.23
X$19932 171 616 172 644 645 cell_1rw
* cell instance $19933 m0 *1 37.365,141.96
X$19933 171 618 172 644 645 cell_1rw
* cell instance $19934 r0 *1 37.365,141.96
X$19934 171 619 172 644 645 cell_1rw
* cell instance $19935 m0 *1 37.365,144.69
X$19935 171 620 172 644 645 cell_1rw
* cell instance $19936 r0 *1 37.365,144.69
X$19936 171 621 172 644 645 cell_1rw
* cell instance $19937 m0 *1 37.365,147.42
X$19937 171 622 172 644 645 cell_1rw
* cell instance $19938 r0 *1 37.365,147.42
X$19938 171 623 172 644 645 cell_1rw
* cell instance $19939 m0 *1 37.365,150.15
X$19939 171 624 172 644 645 cell_1rw
* cell instance $19940 m0 *1 37.365,152.88
X$19940 171 626 172 644 645 cell_1rw
* cell instance $19941 r0 *1 37.365,150.15
X$19941 171 625 172 644 645 cell_1rw
* cell instance $19942 r0 *1 37.365,152.88
X$19942 171 627 172 644 645 cell_1rw
* cell instance $19943 m0 *1 37.365,155.61
X$19943 171 628 172 644 645 cell_1rw
* cell instance $19944 r0 *1 37.365,155.61
X$19944 171 629 172 644 645 cell_1rw
* cell instance $19945 m0 *1 37.365,158.34
X$19945 171 630 172 644 645 cell_1rw
* cell instance $19946 r0 *1 37.365,158.34
X$19946 171 631 172 644 645 cell_1rw
* cell instance $19947 m0 *1 37.365,161.07
X$19947 171 632 172 644 645 cell_1rw
* cell instance $19948 r0 *1 37.365,161.07
X$19948 171 633 172 644 645 cell_1rw
* cell instance $19949 m0 *1 37.365,163.8
X$19949 171 634 172 644 645 cell_1rw
* cell instance $19950 r0 *1 37.365,163.8
X$19950 171 635 172 644 645 cell_1rw
* cell instance $19951 m0 *1 37.365,166.53
X$19951 171 637 172 644 645 cell_1rw
* cell instance $19952 r0 *1 37.365,166.53
X$19952 171 636 172 644 645 cell_1rw
* cell instance $19953 m0 *1 37.365,169.26
X$19953 171 639 172 644 645 cell_1rw
* cell instance $19954 r0 *1 37.365,169.26
X$19954 171 638 172 644 645 cell_1rw
* cell instance $19955 m0 *1 37.365,171.99
X$19955 171 640 172 644 645 cell_1rw
* cell instance $19956 r0 *1 37.365,171.99
X$19956 171 641 172 644 645 cell_1rw
* cell instance $19957 m0 *1 37.365,174.72
X$19957 171 642 172 644 645 cell_1rw
* cell instance $19958 r0 *1 37.365,174.72
X$19958 171 643 172 644 645 cell_1rw
* cell instance $19959 r0 *1 38.07,87.36
X$19959 173 322 174 644 645 cell_1rw
* cell instance $19960 m0 *1 38.07,90.09
X$19960 173 581 174 644 645 cell_1rw
* cell instance $19961 r0 *1 38.07,90.09
X$19961 173 580 174 644 645 cell_1rw
* cell instance $19962 m0 *1 38.07,92.82
X$19962 173 583 174 644 645 cell_1rw
* cell instance $19963 r0 *1 38.07,92.82
X$19963 173 582 174 644 645 cell_1rw
* cell instance $19964 m0 *1 38.07,95.55
X$19964 173 584 174 644 645 cell_1rw
* cell instance $19965 r0 *1 38.07,95.55
X$19965 173 585 174 644 645 cell_1rw
* cell instance $19966 m0 *1 38.07,98.28
X$19966 173 586 174 644 645 cell_1rw
* cell instance $19967 r0 *1 38.07,98.28
X$19967 173 587 174 644 645 cell_1rw
* cell instance $19968 m0 *1 38.07,101.01
X$19968 173 588 174 644 645 cell_1rw
* cell instance $19969 r0 *1 38.07,101.01
X$19969 173 589 174 644 645 cell_1rw
* cell instance $19970 m0 *1 38.07,103.74
X$19970 173 590 174 644 645 cell_1rw
* cell instance $19971 r0 *1 38.07,103.74
X$19971 173 591 174 644 645 cell_1rw
* cell instance $19972 m0 *1 38.07,106.47
X$19972 173 593 174 644 645 cell_1rw
* cell instance $19973 r0 *1 38.07,106.47
X$19973 173 592 174 644 645 cell_1rw
* cell instance $19974 m0 *1 38.07,109.2
X$19974 173 594 174 644 645 cell_1rw
* cell instance $19975 r0 *1 38.07,109.2
X$19975 173 595 174 644 645 cell_1rw
* cell instance $19976 m0 *1 38.07,111.93
X$19976 173 597 174 644 645 cell_1rw
* cell instance $19977 r0 *1 38.07,111.93
X$19977 173 596 174 644 645 cell_1rw
* cell instance $19978 m0 *1 38.07,114.66
X$19978 173 598 174 644 645 cell_1rw
* cell instance $19979 r0 *1 38.07,114.66
X$19979 173 599 174 644 645 cell_1rw
* cell instance $19980 m0 *1 38.07,117.39
X$19980 173 600 174 644 645 cell_1rw
* cell instance $19981 r0 *1 38.07,117.39
X$19981 173 601 174 644 645 cell_1rw
* cell instance $19982 m0 *1 38.07,120.12
X$19982 173 602 174 644 645 cell_1rw
* cell instance $19983 r0 *1 38.07,120.12
X$19983 173 603 174 644 645 cell_1rw
* cell instance $19984 m0 *1 38.07,122.85
X$19984 173 604 174 644 645 cell_1rw
* cell instance $19985 r0 *1 38.07,122.85
X$19985 173 605 174 644 645 cell_1rw
* cell instance $19986 m0 *1 38.07,125.58
X$19986 173 606 174 644 645 cell_1rw
* cell instance $19987 r0 *1 38.07,125.58
X$19987 173 607 174 644 645 cell_1rw
* cell instance $19988 m0 *1 38.07,128.31
X$19988 173 609 174 644 645 cell_1rw
* cell instance $19989 r0 *1 38.07,128.31
X$19989 173 608 174 644 645 cell_1rw
* cell instance $19990 m0 *1 38.07,131.04
X$19990 173 610 174 644 645 cell_1rw
* cell instance $19991 r0 *1 38.07,131.04
X$19991 173 611 174 644 645 cell_1rw
* cell instance $19992 m0 *1 38.07,133.77
X$19992 173 612 174 644 645 cell_1rw
* cell instance $19993 r0 *1 38.07,133.77
X$19993 173 613 174 644 645 cell_1rw
* cell instance $19994 m0 *1 38.07,136.5
X$19994 173 615 174 644 645 cell_1rw
* cell instance $19995 r0 *1 38.07,136.5
X$19995 173 614 174 644 645 cell_1rw
* cell instance $19996 m0 *1 38.07,139.23
X$19996 173 617 174 644 645 cell_1rw
* cell instance $19997 r0 *1 38.07,139.23
X$19997 173 616 174 644 645 cell_1rw
* cell instance $19998 m0 *1 38.07,141.96
X$19998 173 618 174 644 645 cell_1rw
* cell instance $19999 r0 *1 38.07,141.96
X$19999 173 619 174 644 645 cell_1rw
* cell instance $20000 m0 *1 38.07,144.69
X$20000 173 620 174 644 645 cell_1rw
* cell instance $20001 r0 *1 38.07,144.69
X$20001 173 621 174 644 645 cell_1rw
* cell instance $20002 m0 *1 38.07,147.42
X$20002 173 622 174 644 645 cell_1rw
* cell instance $20003 m0 *1 38.07,150.15
X$20003 173 624 174 644 645 cell_1rw
* cell instance $20004 r0 *1 38.07,147.42
X$20004 173 623 174 644 645 cell_1rw
* cell instance $20005 r0 *1 38.07,150.15
X$20005 173 625 174 644 645 cell_1rw
* cell instance $20006 m0 *1 38.07,152.88
X$20006 173 626 174 644 645 cell_1rw
* cell instance $20007 r0 *1 38.07,152.88
X$20007 173 627 174 644 645 cell_1rw
* cell instance $20008 m0 *1 38.07,155.61
X$20008 173 628 174 644 645 cell_1rw
* cell instance $20009 r0 *1 38.07,155.61
X$20009 173 629 174 644 645 cell_1rw
* cell instance $20010 m0 *1 38.07,158.34
X$20010 173 630 174 644 645 cell_1rw
* cell instance $20011 r0 *1 38.07,158.34
X$20011 173 631 174 644 645 cell_1rw
* cell instance $20012 m0 *1 38.07,161.07
X$20012 173 632 174 644 645 cell_1rw
* cell instance $20013 r0 *1 38.07,161.07
X$20013 173 633 174 644 645 cell_1rw
* cell instance $20014 m0 *1 38.07,163.8
X$20014 173 634 174 644 645 cell_1rw
* cell instance $20015 r0 *1 38.07,163.8
X$20015 173 635 174 644 645 cell_1rw
* cell instance $20016 m0 *1 38.07,166.53
X$20016 173 637 174 644 645 cell_1rw
* cell instance $20017 m0 *1 38.07,169.26
X$20017 173 639 174 644 645 cell_1rw
* cell instance $20018 r0 *1 38.07,166.53
X$20018 173 636 174 644 645 cell_1rw
* cell instance $20019 r0 *1 38.07,169.26
X$20019 173 638 174 644 645 cell_1rw
* cell instance $20020 m0 *1 38.07,171.99
X$20020 173 640 174 644 645 cell_1rw
* cell instance $20021 r0 *1 38.07,171.99
X$20021 173 641 174 644 645 cell_1rw
* cell instance $20022 m0 *1 38.07,174.72
X$20022 173 642 174 644 645 cell_1rw
* cell instance $20023 r0 *1 38.07,174.72
X$20023 173 643 174 644 645 cell_1rw
* cell instance $20024 r0 *1 38.775,87.36
X$20024 175 322 176 644 645 cell_1rw
* cell instance $20025 m0 *1 38.775,90.09
X$20025 175 581 176 644 645 cell_1rw
* cell instance $20026 r0 *1 38.775,90.09
X$20026 175 580 176 644 645 cell_1rw
* cell instance $20027 m0 *1 38.775,92.82
X$20027 175 583 176 644 645 cell_1rw
* cell instance $20028 m0 *1 38.775,95.55
X$20028 175 584 176 644 645 cell_1rw
* cell instance $20029 r0 *1 38.775,92.82
X$20029 175 582 176 644 645 cell_1rw
* cell instance $20030 r0 *1 38.775,95.55
X$20030 175 585 176 644 645 cell_1rw
* cell instance $20031 m0 *1 38.775,98.28
X$20031 175 586 176 644 645 cell_1rw
* cell instance $20032 m0 *1 38.775,101.01
X$20032 175 588 176 644 645 cell_1rw
* cell instance $20033 r0 *1 38.775,98.28
X$20033 175 587 176 644 645 cell_1rw
* cell instance $20034 m0 *1 38.775,103.74
X$20034 175 590 176 644 645 cell_1rw
* cell instance $20035 r0 *1 38.775,101.01
X$20035 175 589 176 644 645 cell_1rw
* cell instance $20036 r0 *1 38.775,103.74
X$20036 175 591 176 644 645 cell_1rw
* cell instance $20037 m0 *1 38.775,106.47
X$20037 175 593 176 644 645 cell_1rw
* cell instance $20038 m0 *1 38.775,109.2
X$20038 175 594 176 644 645 cell_1rw
* cell instance $20039 r0 *1 38.775,106.47
X$20039 175 592 176 644 645 cell_1rw
* cell instance $20040 r0 *1 38.775,109.2
X$20040 175 595 176 644 645 cell_1rw
* cell instance $20041 m0 *1 38.775,111.93
X$20041 175 597 176 644 645 cell_1rw
* cell instance $20042 m0 *1 38.775,114.66
X$20042 175 598 176 644 645 cell_1rw
* cell instance $20043 r0 *1 38.775,111.93
X$20043 175 596 176 644 645 cell_1rw
* cell instance $20044 r0 *1 38.775,114.66
X$20044 175 599 176 644 645 cell_1rw
* cell instance $20045 m0 *1 38.775,117.39
X$20045 175 600 176 644 645 cell_1rw
* cell instance $20046 r0 *1 38.775,117.39
X$20046 175 601 176 644 645 cell_1rw
* cell instance $20047 m0 *1 38.775,120.12
X$20047 175 602 176 644 645 cell_1rw
* cell instance $20048 m0 *1 38.775,122.85
X$20048 175 604 176 644 645 cell_1rw
* cell instance $20049 r0 *1 38.775,120.12
X$20049 175 603 176 644 645 cell_1rw
* cell instance $20050 r0 *1 38.775,122.85
X$20050 175 605 176 644 645 cell_1rw
* cell instance $20051 m0 *1 38.775,125.58
X$20051 175 606 176 644 645 cell_1rw
* cell instance $20052 r0 *1 38.775,125.58
X$20052 175 607 176 644 645 cell_1rw
* cell instance $20053 m0 *1 38.775,128.31
X$20053 175 609 176 644 645 cell_1rw
* cell instance $20054 r0 *1 38.775,128.31
X$20054 175 608 176 644 645 cell_1rw
* cell instance $20055 m0 *1 38.775,131.04
X$20055 175 610 176 644 645 cell_1rw
* cell instance $20056 r0 *1 38.775,131.04
X$20056 175 611 176 644 645 cell_1rw
* cell instance $20057 m0 *1 38.775,133.77
X$20057 175 612 176 644 645 cell_1rw
* cell instance $20058 r0 *1 38.775,133.77
X$20058 175 613 176 644 645 cell_1rw
* cell instance $20059 m0 *1 38.775,136.5
X$20059 175 615 176 644 645 cell_1rw
* cell instance $20060 r0 *1 38.775,136.5
X$20060 175 614 176 644 645 cell_1rw
* cell instance $20061 m0 *1 38.775,139.23
X$20061 175 617 176 644 645 cell_1rw
* cell instance $20062 r0 *1 38.775,139.23
X$20062 175 616 176 644 645 cell_1rw
* cell instance $20063 m0 *1 38.775,141.96
X$20063 175 618 176 644 645 cell_1rw
* cell instance $20064 r0 *1 38.775,141.96
X$20064 175 619 176 644 645 cell_1rw
* cell instance $20065 m0 *1 38.775,144.69
X$20065 175 620 176 644 645 cell_1rw
* cell instance $20066 r0 *1 38.775,144.69
X$20066 175 621 176 644 645 cell_1rw
* cell instance $20067 m0 *1 38.775,147.42
X$20067 175 622 176 644 645 cell_1rw
* cell instance $20068 r0 *1 38.775,147.42
X$20068 175 623 176 644 645 cell_1rw
* cell instance $20069 m0 *1 38.775,150.15
X$20069 175 624 176 644 645 cell_1rw
* cell instance $20070 m0 *1 38.775,152.88
X$20070 175 626 176 644 645 cell_1rw
* cell instance $20071 r0 *1 38.775,150.15
X$20071 175 625 176 644 645 cell_1rw
* cell instance $20072 r0 *1 38.775,152.88
X$20072 175 627 176 644 645 cell_1rw
* cell instance $20073 m0 *1 38.775,155.61
X$20073 175 628 176 644 645 cell_1rw
* cell instance $20074 r0 *1 38.775,155.61
X$20074 175 629 176 644 645 cell_1rw
* cell instance $20075 m0 *1 38.775,158.34
X$20075 175 630 176 644 645 cell_1rw
* cell instance $20076 r0 *1 38.775,158.34
X$20076 175 631 176 644 645 cell_1rw
* cell instance $20077 m0 *1 38.775,161.07
X$20077 175 632 176 644 645 cell_1rw
* cell instance $20078 m0 *1 38.775,163.8
X$20078 175 634 176 644 645 cell_1rw
* cell instance $20079 r0 *1 38.775,161.07
X$20079 175 633 176 644 645 cell_1rw
* cell instance $20080 r0 *1 38.775,163.8
X$20080 175 635 176 644 645 cell_1rw
* cell instance $20081 m0 *1 38.775,166.53
X$20081 175 637 176 644 645 cell_1rw
* cell instance $20082 r0 *1 38.775,166.53
X$20082 175 636 176 644 645 cell_1rw
* cell instance $20083 m0 *1 38.775,169.26
X$20083 175 639 176 644 645 cell_1rw
* cell instance $20084 r0 *1 38.775,169.26
X$20084 175 638 176 644 645 cell_1rw
* cell instance $20085 m0 *1 38.775,171.99
X$20085 175 640 176 644 645 cell_1rw
* cell instance $20086 r0 *1 38.775,171.99
X$20086 175 641 176 644 645 cell_1rw
* cell instance $20087 m0 *1 38.775,174.72
X$20087 175 642 176 644 645 cell_1rw
* cell instance $20088 r0 *1 38.775,174.72
X$20088 175 643 176 644 645 cell_1rw
* cell instance $20089 r0 *1 39.48,87.36
X$20089 177 322 178 644 645 cell_1rw
* cell instance $20090 m0 *1 39.48,90.09
X$20090 177 581 178 644 645 cell_1rw
* cell instance $20091 m0 *1 39.48,92.82
X$20091 177 583 178 644 645 cell_1rw
* cell instance $20092 r0 *1 39.48,90.09
X$20092 177 580 178 644 645 cell_1rw
* cell instance $20093 m0 *1 39.48,95.55
X$20093 177 584 178 644 645 cell_1rw
* cell instance $20094 r0 *1 39.48,92.82
X$20094 177 582 178 644 645 cell_1rw
* cell instance $20095 r0 *1 39.48,95.55
X$20095 177 585 178 644 645 cell_1rw
* cell instance $20096 m0 *1 39.48,98.28
X$20096 177 586 178 644 645 cell_1rw
* cell instance $20097 r0 *1 39.48,98.28
X$20097 177 587 178 644 645 cell_1rw
* cell instance $20098 m0 *1 39.48,101.01
X$20098 177 588 178 644 645 cell_1rw
* cell instance $20099 m0 *1 39.48,103.74
X$20099 177 590 178 644 645 cell_1rw
* cell instance $20100 r0 *1 39.48,101.01
X$20100 177 589 178 644 645 cell_1rw
* cell instance $20101 m0 *1 39.48,106.47
X$20101 177 593 178 644 645 cell_1rw
* cell instance $20102 r0 *1 39.48,103.74
X$20102 177 591 178 644 645 cell_1rw
* cell instance $20103 r0 *1 39.48,106.47
X$20103 177 592 178 644 645 cell_1rw
* cell instance $20104 m0 *1 39.48,109.2
X$20104 177 594 178 644 645 cell_1rw
* cell instance $20105 r0 *1 39.48,109.2
X$20105 177 595 178 644 645 cell_1rw
* cell instance $20106 m0 *1 39.48,111.93
X$20106 177 597 178 644 645 cell_1rw
* cell instance $20107 r0 *1 39.48,111.93
X$20107 177 596 178 644 645 cell_1rw
* cell instance $20108 m0 *1 39.48,114.66
X$20108 177 598 178 644 645 cell_1rw
* cell instance $20109 r0 *1 39.48,114.66
X$20109 177 599 178 644 645 cell_1rw
* cell instance $20110 m0 *1 39.48,117.39
X$20110 177 600 178 644 645 cell_1rw
* cell instance $20111 r0 *1 39.48,117.39
X$20111 177 601 178 644 645 cell_1rw
* cell instance $20112 m0 *1 39.48,120.12
X$20112 177 602 178 644 645 cell_1rw
* cell instance $20113 r0 *1 39.48,120.12
X$20113 177 603 178 644 645 cell_1rw
* cell instance $20114 m0 *1 39.48,122.85
X$20114 177 604 178 644 645 cell_1rw
* cell instance $20115 m0 *1 39.48,125.58
X$20115 177 606 178 644 645 cell_1rw
* cell instance $20116 r0 *1 39.48,122.85
X$20116 177 605 178 644 645 cell_1rw
* cell instance $20117 r0 *1 39.48,125.58
X$20117 177 607 178 644 645 cell_1rw
* cell instance $20118 m0 *1 39.48,128.31
X$20118 177 609 178 644 645 cell_1rw
* cell instance $20119 m0 *1 39.48,131.04
X$20119 177 610 178 644 645 cell_1rw
* cell instance $20120 r0 *1 39.48,128.31
X$20120 177 608 178 644 645 cell_1rw
* cell instance $20121 m0 *1 39.48,133.77
X$20121 177 612 178 644 645 cell_1rw
* cell instance $20122 r0 *1 39.48,131.04
X$20122 177 611 178 644 645 cell_1rw
* cell instance $20123 r0 *1 39.48,133.77
X$20123 177 613 178 644 645 cell_1rw
* cell instance $20124 m0 *1 39.48,136.5
X$20124 177 615 178 644 645 cell_1rw
* cell instance $20125 r0 *1 39.48,136.5
X$20125 177 614 178 644 645 cell_1rw
* cell instance $20126 m0 *1 39.48,139.23
X$20126 177 617 178 644 645 cell_1rw
* cell instance $20127 r0 *1 39.48,139.23
X$20127 177 616 178 644 645 cell_1rw
* cell instance $20128 m0 *1 39.48,141.96
X$20128 177 618 178 644 645 cell_1rw
* cell instance $20129 r0 *1 39.48,141.96
X$20129 177 619 178 644 645 cell_1rw
* cell instance $20130 m0 *1 39.48,144.69
X$20130 177 620 178 644 645 cell_1rw
* cell instance $20131 m0 *1 39.48,147.42
X$20131 177 622 178 644 645 cell_1rw
* cell instance $20132 r0 *1 39.48,144.69
X$20132 177 621 178 644 645 cell_1rw
* cell instance $20133 m0 *1 39.48,150.15
X$20133 177 624 178 644 645 cell_1rw
* cell instance $20134 r0 *1 39.48,147.42
X$20134 177 623 178 644 645 cell_1rw
* cell instance $20135 m0 *1 39.48,152.88
X$20135 177 626 178 644 645 cell_1rw
* cell instance $20136 r0 *1 39.48,150.15
X$20136 177 625 178 644 645 cell_1rw
* cell instance $20137 r0 *1 39.48,152.88
X$20137 177 627 178 644 645 cell_1rw
* cell instance $20138 m0 *1 39.48,155.61
X$20138 177 628 178 644 645 cell_1rw
* cell instance $20139 r0 *1 39.48,155.61
X$20139 177 629 178 644 645 cell_1rw
* cell instance $20140 m0 *1 39.48,158.34
X$20140 177 630 178 644 645 cell_1rw
* cell instance $20141 r0 *1 39.48,158.34
X$20141 177 631 178 644 645 cell_1rw
* cell instance $20142 m0 *1 39.48,161.07
X$20142 177 632 178 644 645 cell_1rw
* cell instance $20143 r0 *1 39.48,161.07
X$20143 177 633 178 644 645 cell_1rw
* cell instance $20144 m0 *1 39.48,163.8
X$20144 177 634 178 644 645 cell_1rw
* cell instance $20145 r0 *1 39.48,163.8
X$20145 177 635 178 644 645 cell_1rw
* cell instance $20146 m0 *1 39.48,166.53
X$20146 177 637 178 644 645 cell_1rw
* cell instance $20147 r0 *1 39.48,166.53
X$20147 177 636 178 644 645 cell_1rw
* cell instance $20148 m0 *1 39.48,169.26
X$20148 177 639 178 644 645 cell_1rw
* cell instance $20149 r0 *1 39.48,169.26
X$20149 177 638 178 644 645 cell_1rw
* cell instance $20150 m0 *1 39.48,171.99
X$20150 177 640 178 644 645 cell_1rw
* cell instance $20151 m0 *1 39.48,174.72
X$20151 177 642 178 644 645 cell_1rw
* cell instance $20152 r0 *1 39.48,171.99
X$20152 177 641 178 644 645 cell_1rw
* cell instance $20153 r0 *1 39.48,174.72
X$20153 177 643 178 644 645 cell_1rw
* cell instance $20154 r0 *1 40.185,87.36
X$20154 179 322 180 644 645 cell_1rw
* cell instance $20155 m0 *1 40.185,90.09
X$20155 179 581 180 644 645 cell_1rw
* cell instance $20156 r0 *1 40.185,90.09
X$20156 179 580 180 644 645 cell_1rw
* cell instance $20157 m0 *1 40.185,92.82
X$20157 179 583 180 644 645 cell_1rw
* cell instance $20158 r0 *1 40.185,92.82
X$20158 179 582 180 644 645 cell_1rw
* cell instance $20159 m0 *1 40.185,95.55
X$20159 179 584 180 644 645 cell_1rw
* cell instance $20160 r0 *1 40.185,95.55
X$20160 179 585 180 644 645 cell_1rw
* cell instance $20161 m0 *1 40.185,98.28
X$20161 179 586 180 644 645 cell_1rw
* cell instance $20162 r0 *1 40.185,98.28
X$20162 179 587 180 644 645 cell_1rw
* cell instance $20163 m0 *1 40.185,101.01
X$20163 179 588 180 644 645 cell_1rw
* cell instance $20164 m0 *1 40.185,103.74
X$20164 179 590 180 644 645 cell_1rw
* cell instance $20165 r0 *1 40.185,101.01
X$20165 179 589 180 644 645 cell_1rw
* cell instance $20166 r0 *1 40.185,103.74
X$20166 179 591 180 644 645 cell_1rw
* cell instance $20167 m0 *1 40.185,106.47
X$20167 179 593 180 644 645 cell_1rw
* cell instance $20168 r0 *1 40.185,106.47
X$20168 179 592 180 644 645 cell_1rw
* cell instance $20169 m0 *1 40.185,109.2
X$20169 179 594 180 644 645 cell_1rw
* cell instance $20170 r0 *1 40.185,109.2
X$20170 179 595 180 644 645 cell_1rw
* cell instance $20171 m0 *1 40.185,111.93
X$20171 179 597 180 644 645 cell_1rw
* cell instance $20172 r0 *1 40.185,111.93
X$20172 179 596 180 644 645 cell_1rw
* cell instance $20173 m0 *1 40.185,114.66
X$20173 179 598 180 644 645 cell_1rw
* cell instance $20174 r0 *1 40.185,114.66
X$20174 179 599 180 644 645 cell_1rw
* cell instance $20175 m0 *1 40.185,117.39
X$20175 179 600 180 644 645 cell_1rw
* cell instance $20176 m0 *1 40.185,120.12
X$20176 179 602 180 644 645 cell_1rw
* cell instance $20177 r0 *1 40.185,117.39
X$20177 179 601 180 644 645 cell_1rw
* cell instance $20178 r0 *1 40.185,120.12
X$20178 179 603 180 644 645 cell_1rw
* cell instance $20179 m0 *1 40.185,122.85
X$20179 179 604 180 644 645 cell_1rw
* cell instance $20180 r0 *1 40.185,122.85
X$20180 179 605 180 644 645 cell_1rw
* cell instance $20181 m0 *1 40.185,125.58
X$20181 179 606 180 644 645 cell_1rw
* cell instance $20182 r0 *1 40.185,125.58
X$20182 179 607 180 644 645 cell_1rw
* cell instance $20183 m0 *1 40.185,128.31
X$20183 179 609 180 644 645 cell_1rw
* cell instance $20184 r0 *1 40.185,128.31
X$20184 179 608 180 644 645 cell_1rw
* cell instance $20185 m0 *1 40.185,131.04
X$20185 179 610 180 644 645 cell_1rw
* cell instance $20186 r0 *1 40.185,131.04
X$20186 179 611 180 644 645 cell_1rw
* cell instance $20187 m0 *1 40.185,133.77
X$20187 179 612 180 644 645 cell_1rw
* cell instance $20188 m0 *1 40.185,136.5
X$20188 179 615 180 644 645 cell_1rw
* cell instance $20189 r0 *1 40.185,133.77
X$20189 179 613 180 644 645 cell_1rw
* cell instance $20190 r0 *1 40.185,136.5
X$20190 179 614 180 644 645 cell_1rw
* cell instance $20191 m0 *1 40.185,139.23
X$20191 179 617 180 644 645 cell_1rw
* cell instance $20192 r0 *1 40.185,139.23
X$20192 179 616 180 644 645 cell_1rw
* cell instance $20193 m0 *1 40.185,141.96
X$20193 179 618 180 644 645 cell_1rw
* cell instance $20194 r0 *1 40.185,141.96
X$20194 179 619 180 644 645 cell_1rw
* cell instance $20195 m0 *1 40.185,144.69
X$20195 179 620 180 644 645 cell_1rw
* cell instance $20196 r0 *1 40.185,144.69
X$20196 179 621 180 644 645 cell_1rw
* cell instance $20197 m0 *1 40.185,147.42
X$20197 179 622 180 644 645 cell_1rw
* cell instance $20198 r0 *1 40.185,147.42
X$20198 179 623 180 644 645 cell_1rw
* cell instance $20199 m0 *1 40.185,150.15
X$20199 179 624 180 644 645 cell_1rw
* cell instance $20200 m0 *1 40.185,152.88
X$20200 179 626 180 644 645 cell_1rw
* cell instance $20201 r0 *1 40.185,150.15
X$20201 179 625 180 644 645 cell_1rw
* cell instance $20202 m0 *1 40.185,155.61
X$20202 179 628 180 644 645 cell_1rw
* cell instance $20203 r0 *1 40.185,152.88
X$20203 179 627 180 644 645 cell_1rw
* cell instance $20204 m0 *1 40.185,158.34
X$20204 179 630 180 644 645 cell_1rw
* cell instance $20205 r0 *1 40.185,155.61
X$20205 179 629 180 644 645 cell_1rw
* cell instance $20206 m0 *1 40.185,161.07
X$20206 179 632 180 644 645 cell_1rw
* cell instance $20207 r0 *1 40.185,158.34
X$20207 179 631 180 644 645 cell_1rw
* cell instance $20208 r0 *1 40.185,161.07
X$20208 179 633 180 644 645 cell_1rw
* cell instance $20209 m0 *1 40.185,163.8
X$20209 179 634 180 644 645 cell_1rw
* cell instance $20210 r0 *1 40.185,163.8
X$20210 179 635 180 644 645 cell_1rw
* cell instance $20211 m0 *1 40.185,166.53
X$20211 179 637 180 644 645 cell_1rw
* cell instance $20212 r0 *1 40.185,166.53
X$20212 179 636 180 644 645 cell_1rw
* cell instance $20213 m0 *1 40.185,169.26
X$20213 179 639 180 644 645 cell_1rw
* cell instance $20214 r0 *1 40.185,169.26
X$20214 179 638 180 644 645 cell_1rw
* cell instance $20215 m0 *1 40.185,171.99
X$20215 179 640 180 644 645 cell_1rw
* cell instance $20216 r0 *1 40.185,171.99
X$20216 179 641 180 644 645 cell_1rw
* cell instance $20217 m0 *1 40.185,174.72
X$20217 179 642 180 644 645 cell_1rw
* cell instance $20218 r0 *1 40.185,174.72
X$20218 179 643 180 644 645 cell_1rw
* cell instance $20219 r0 *1 40.89,87.36
X$20219 181 322 182 644 645 cell_1rw
* cell instance $20220 m0 *1 40.89,90.09
X$20220 181 581 182 644 645 cell_1rw
* cell instance $20221 r0 *1 40.89,90.09
X$20221 181 580 182 644 645 cell_1rw
* cell instance $20222 m0 *1 40.89,92.82
X$20222 181 583 182 644 645 cell_1rw
* cell instance $20223 r0 *1 40.89,92.82
X$20223 181 582 182 644 645 cell_1rw
* cell instance $20224 m0 *1 40.89,95.55
X$20224 181 584 182 644 645 cell_1rw
* cell instance $20225 r0 *1 40.89,95.55
X$20225 181 585 182 644 645 cell_1rw
* cell instance $20226 m0 *1 40.89,98.28
X$20226 181 586 182 644 645 cell_1rw
* cell instance $20227 r0 *1 40.89,98.28
X$20227 181 587 182 644 645 cell_1rw
* cell instance $20228 m0 *1 40.89,101.01
X$20228 181 588 182 644 645 cell_1rw
* cell instance $20229 r0 *1 40.89,101.01
X$20229 181 589 182 644 645 cell_1rw
* cell instance $20230 m0 *1 40.89,103.74
X$20230 181 590 182 644 645 cell_1rw
* cell instance $20231 r0 *1 40.89,103.74
X$20231 181 591 182 644 645 cell_1rw
* cell instance $20232 m0 *1 40.89,106.47
X$20232 181 593 182 644 645 cell_1rw
* cell instance $20233 r0 *1 40.89,106.47
X$20233 181 592 182 644 645 cell_1rw
* cell instance $20234 m0 *1 40.89,109.2
X$20234 181 594 182 644 645 cell_1rw
* cell instance $20235 r0 *1 40.89,109.2
X$20235 181 595 182 644 645 cell_1rw
* cell instance $20236 m0 *1 40.89,111.93
X$20236 181 597 182 644 645 cell_1rw
* cell instance $20237 r0 *1 40.89,111.93
X$20237 181 596 182 644 645 cell_1rw
* cell instance $20238 m0 *1 40.89,114.66
X$20238 181 598 182 644 645 cell_1rw
* cell instance $20239 r0 *1 40.89,114.66
X$20239 181 599 182 644 645 cell_1rw
* cell instance $20240 m0 *1 40.89,117.39
X$20240 181 600 182 644 645 cell_1rw
* cell instance $20241 r0 *1 40.89,117.39
X$20241 181 601 182 644 645 cell_1rw
* cell instance $20242 m0 *1 40.89,120.12
X$20242 181 602 182 644 645 cell_1rw
* cell instance $20243 m0 *1 40.89,122.85
X$20243 181 604 182 644 645 cell_1rw
* cell instance $20244 r0 *1 40.89,120.12
X$20244 181 603 182 644 645 cell_1rw
* cell instance $20245 r0 *1 40.89,122.85
X$20245 181 605 182 644 645 cell_1rw
* cell instance $20246 m0 *1 40.89,125.58
X$20246 181 606 182 644 645 cell_1rw
* cell instance $20247 r0 *1 40.89,125.58
X$20247 181 607 182 644 645 cell_1rw
* cell instance $20248 m0 *1 40.89,128.31
X$20248 181 609 182 644 645 cell_1rw
* cell instance $20249 m0 *1 40.89,131.04
X$20249 181 610 182 644 645 cell_1rw
* cell instance $20250 r0 *1 40.89,128.31
X$20250 181 608 182 644 645 cell_1rw
* cell instance $20251 r0 *1 40.89,131.04
X$20251 181 611 182 644 645 cell_1rw
* cell instance $20252 m0 *1 40.89,133.77
X$20252 181 612 182 644 645 cell_1rw
* cell instance $20253 r0 *1 40.89,133.77
X$20253 181 613 182 644 645 cell_1rw
* cell instance $20254 m0 *1 40.89,136.5
X$20254 181 615 182 644 645 cell_1rw
* cell instance $20255 r0 *1 40.89,136.5
X$20255 181 614 182 644 645 cell_1rw
* cell instance $20256 m0 *1 40.89,139.23
X$20256 181 617 182 644 645 cell_1rw
* cell instance $20257 r0 *1 40.89,139.23
X$20257 181 616 182 644 645 cell_1rw
* cell instance $20258 m0 *1 40.89,141.96
X$20258 181 618 182 644 645 cell_1rw
* cell instance $20259 r0 *1 40.89,141.96
X$20259 181 619 182 644 645 cell_1rw
* cell instance $20260 m0 *1 40.89,144.69
X$20260 181 620 182 644 645 cell_1rw
* cell instance $20261 r0 *1 40.89,144.69
X$20261 181 621 182 644 645 cell_1rw
* cell instance $20262 m0 *1 40.89,147.42
X$20262 181 622 182 644 645 cell_1rw
* cell instance $20263 m0 *1 40.89,150.15
X$20263 181 624 182 644 645 cell_1rw
* cell instance $20264 r0 *1 40.89,147.42
X$20264 181 623 182 644 645 cell_1rw
* cell instance $20265 r0 *1 40.89,150.15
X$20265 181 625 182 644 645 cell_1rw
* cell instance $20266 m0 *1 40.89,152.88
X$20266 181 626 182 644 645 cell_1rw
* cell instance $20267 r0 *1 40.89,152.88
X$20267 181 627 182 644 645 cell_1rw
* cell instance $20268 m0 *1 40.89,155.61
X$20268 181 628 182 644 645 cell_1rw
* cell instance $20269 m0 *1 40.89,158.34
X$20269 181 630 182 644 645 cell_1rw
* cell instance $20270 r0 *1 40.89,155.61
X$20270 181 629 182 644 645 cell_1rw
* cell instance $20271 m0 *1 40.89,161.07
X$20271 181 632 182 644 645 cell_1rw
* cell instance $20272 r0 *1 40.89,158.34
X$20272 181 631 182 644 645 cell_1rw
* cell instance $20273 r0 *1 40.89,161.07
X$20273 181 633 182 644 645 cell_1rw
* cell instance $20274 m0 *1 40.89,163.8
X$20274 181 634 182 644 645 cell_1rw
* cell instance $20275 m0 *1 40.89,166.53
X$20275 181 637 182 644 645 cell_1rw
* cell instance $20276 r0 *1 40.89,163.8
X$20276 181 635 182 644 645 cell_1rw
* cell instance $20277 r0 *1 40.89,166.53
X$20277 181 636 182 644 645 cell_1rw
* cell instance $20278 m0 *1 40.89,169.26
X$20278 181 639 182 644 645 cell_1rw
* cell instance $20279 r0 *1 40.89,169.26
X$20279 181 638 182 644 645 cell_1rw
* cell instance $20280 m0 *1 40.89,171.99
X$20280 181 640 182 644 645 cell_1rw
* cell instance $20281 m0 *1 40.89,174.72
X$20281 181 642 182 644 645 cell_1rw
* cell instance $20282 r0 *1 40.89,171.99
X$20282 181 641 182 644 645 cell_1rw
* cell instance $20283 r0 *1 40.89,174.72
X$20283 181 643 182 644 645 cell_1rw
* cell instance $20284 m0 *1 41.595,90.09
X$20284 183 581 184 644 645 cell_1rw
* cell instance $20285 r0 *1 41.595,87.36
X$20285 183 322 184 644 645 cell_1rw
* cell instance $20286 m0 *1 41.595,92.82
X$20286 183 583 184 644 645 cell_1rw
* cell instance $20287 r0 *1 41.595,90.09
X$20287 183 580 184 644 645 cell_1rw
* cell instance $20288 r0 *1 41.595,92.82
X$20288 183 582 184 644 645 cell_1rw
* cell instance $20289 m0 *1 41.595,95.55
X$20289 183 584 184 644 645 cell_1rw
* cell instance $20290 r0 *1 41.595,95.55
X$20290 183 585 184 644 645 cell_1rw
* cell instance $20291 m0 *1 41.595,98.28
X$20291 183 586 184 644 645 cell_1rw
* cell instance $20292 r0 *1 41.595,98.28
X$20292 183 587 184 644 645 cell_1rw
* cell instance $20293 m0 *1 41.595,101.01
X$20293 183 588 184 644 645 cell_1rw
* cell instance $20294 r0 *1 41.595,101.01
X$20294 183 589 184 644 645 cell_1rw
* cell instance $20295 m0 *1 41.595,103.74
X$20295 183 590 184 644 645 cell_1rw
* cell instance $20296 r0 *1 41.595,103.74
X$20296 183 591 184 644 645 cell_1rw
* cell instance $20297 m0 *1 41.595,106.47
X$20297 183 593 184 644 645 cell_1rw
* cell instance $20298 r0 *1 41.595,106.47
X$20298 183 592 184 644 645 cell_1rw
* cell instance $20299 m0 *1 41.595,109.2
X$20299 183 594 184 644 645 cell_1rw
* cell instance $20300 r0 *1 41.595,109.2
X$20300 183 595 184 644 645 cell_1rw
* cell instance $20301 m0 *1 41.595,111.93
X$20301 183 597 184 644 645 cell_1rw
* cell instance $20302 r0 *1 41.595,111.93
X$20302 183 596 184 644 645 cell_1rw
* cell instance $20303 m0 *1 41.595,114.66
X$20303 183 598 184 644 645 cell_1rw
* cell instance $20304 r0 *1 41.595,114.66
X$20304 183 599 184 644 645 cell_1rw
* cell instance $20305 m0 *1 41.595,117.39
X$20305 183 600 184 644 645 cell_1rw
* cell instance $20306 m0 *1 41.595,120.12
X$20306 183 602 184 644 645 cell_1rw
* cell instance $20307 r0 *1 41.595,117.39
X$20307 183 601 184 644 645 cell_1rw
* cell instance $20308 r0 *1 41.595,120.12
X$20308 183 603 184 644 645 cell_1rw
* cell instance $20309 m0 *1 41.595,122.85
X$20309 183 604 184 644 645 cell_1rw
* cell instance $20310 r0 *1 41.595,122.85
X$20310 183 605 184 644 645 cell_1rw
* cell instance $20311 m0 *1 41.595,125.58
X$20311 183 606 184 644 645 cell_1rw
* cell instance $20312 r0 *1 41.595,125.58
X$20312 183 607 184 644 645 cell_1rw
* cell instance $20313 m0 *1 41.595,128.31
X$20313 183 609 184 644 645 cell_1rw
* cell instance $20314 r0 *1 41.595,128.31
X$20314 183 608 184 644 645 cell_1rw
* cell instance $20315 m0 *1 41.595,131.04
X$20315 183 610 184 644 645 cell_1rw
* cell instance $20316 m0 *1 41.595,133.77
X$20316 183 612 184 644 645 cell_1rw
* cell instance $20317 r0 *1 41.595,131.04
X$20317 183 611 184 644 645 cell_1rw
* cell instance $20318 r0 *1 41.595,133.77
X$20318 183 613 184 644 645 cell_1rw
* cell instance $20319 m0 *1 41.595,136.5
X$20319 183 615 184 644 645 cell_1rw
* cell instance $20320 r0 *1 41.595,136.5
X$20320 183 614 184 644 645 cell_1rw
* cell instance $20321 m0 *1 41.595,139.23
X$20321 183 617 184 644 645 cell_1rw
* cell instance $20322 r0 *1 41.595,139.23
X$20322 183 616 184 644 645 cell_1rw
* cell instance $20323 m0 *1 41.595,141.96
X$20323 183 618 184 644 645 cell_1rw
* cell instance $20324 r0 *1 41.595,141.96
X$20324 183 619 184 644 645 cell_1rw
* cell instance $20325 m0 *1 41.595,144.69
X$20325 183 620 184 644 645 cell_1rw
* cell instance $20326 r0 *1 41.595,144.69
X$20326 183 621 184 644 645 cell_1rw
* cell instance $20327 m0 *1 41.595,147.42
X$20327 183 622 184 644 645 cell_1rw
* cell instance $20328 r0 *1 41.595,147.42
X$20328 183 623 184 644 645 cell_1rw
* cell instance $20329 m0 *1 41.595,150.15
X$20329 183 624 184 644 645 cell_1rw
* cell instance $20330 r0 *1 41.595,150.15
X$20330 183 625 184 644 645 cell_1rw
* cell instance $20331 m0 *1 41.595,152.88
X$20331 183 626 184 644 645 cell_1rw
* cell instance $20332 r0 *1 41.595,152.88
X$20332 183 627 184 644 645 cell_1rw
* cell instance $20333 m0 *1 41.595,155.61
X$20333 183 628 184 644 645 cell_1rw
* cell instance $20334 r0 *1 41.595,155.61
X$20334 183 629 184 644 645 cell_1rw
* cell instance $20335 m0 *1 41.595,158.34
X$20335 183 630 184 644 645 cell_1rw
* cell instance $20336 r0 *1 41.595,158.34
X$20336 183 631 184 644 645 cell_1rw
* cell instance $20337 m0 *1 41.595,161.07
X$20337 183 632 184 644 645 cell_1rw
* cell instance $20338 r0 *1 41.595,161.07
X$20338 183 633 184 644 645 cell_1rw
* cell instance $20339 m0 *1 41.595,163.8
X$20339 183 634 184 644 645 cell_1rw
* cell instance $20340 r0 *1 41.595,163.8
X$20340 183 635 184 644 645 cell_1rw
* cell instance $20341 m0 *1 41.595,166.53
X$20341 183 637 184 644 645 cell_1rw
* cell instance $20342 m0 *1 41.595,169.26
X$20342 183 639 184 644 645 cell_1rw
* cell instance $20343 r0 *1 41.595,166.53
X$20343 183 636 184 644 645 cell_1rw
* cell instance $20344 r0 *1 41.595,169.26
X$20344 183 638 184 644 645 cell_1rw
* cell instance $20345 m0 *1 41.595,171.99
X$20345 183 640 184 644 645 cell_1rw
* cell instance $20346 r0 *1 41.595,171.99
X$20346 183 641 184 644 645 cell_1rw
* cell instance $20347 m0 *1 41.595,174.72
X$20347 183 642 184 644 645 cell_1rw
* cell instance $20348 r0 *1 41.595,174.72
X$20348 183 643 184 644 645 cell_1rw
* cell instance $20349 r0 *1 42.3,87.36
X$20349 185 322 186 644 645 cell_1rw
* cell instance $20350 m0 *1 42.3,90.09
X$20350 185 581 186 644 645 cell_1rw
* cell instance $20351 r0 *1 42.3,90.09
X$20351 185 580 186 644 645 cell_1rw
* cell instance $20352 m0 *1 42.3,92.82
X$20352 185 583 186 644 645 cell_1rw
* cell instance $20353 r0 *1 42.3,92.82
X$20353 185 582 186 644 645 cell_1rw
* cell instance $20354 m0 *1 42.3,95.55
X$20354 185 584 186 644 645 cell_1rw
* cell instance $20355 r0 *1 42.3,95.55
X$20355 185 585 186 644 645 cell_1rw
* cell instance $20356 m0 *1 42.3,98.28
X$20356 185 586 186 644 645 cell_1rw
* cell instance $20357 r0 *1 42.3,98.28
X$20357 185 587 186 644 645 cell_1rw
* cell instance $20358 m0 *1 42.3,101.01
X$20358 185 588 186 644 645 cell_1rw
* cell instance $20359 r0 *1 42.3,101.01
X$20359 185 589 186 644 645 cell_1rw
* cell instance $20360 m0 *1 42.3,103.74
X$20360 185 590 186 644 645 cell_1rw
* cell instance $20361 r0 *1 42.3,103.74
X$20361 185 591 186 644 645 cell_1rw
* cell instance $20362 m0 *1 42.3,106.47
X$20362 185 593 186 644 645 cell_1rw
* cell instance $20363 r0 *1 42.3,106.47
X$20363 185 592 186 644 645 cell_1rw
* cell instance $20364 m0 *1 42.3,109.2
X$20364 185 594 186 644 645 cell_1rw
* cell instance $20365 r0 *1 42.3,109.2
X$20365 185 595 186 644 645 cell_1rw
* cell instance $20366 m0 *1 42.3,111.93
X$20366 185 597 186 644 645 cell_1rw
* cell instance $20367 r0 *1 42.3,111.93
X$20367 185 596 186 644 645 cell_1rw
* cell instance $20368 m0 *1 42.3,114.66
X$20368 185 598 186 644 645 cell_1rw
* cell instance $20369 r0 *1 42.3,114.66
X$20369 185 599 186 644 645 cell_1rw
* cell instance $20370 m0 *1 42.3,117.39
X$20370 185 600 186 644 645 cell_1rw
* cell instance $20371 m0 *1 42.3,120.12
X$20371 185 602 186 644 645 cell_1rw
* cell instance $20372 r0 *1 42.3,117.39
X$20372 185 601 186 644 645 cell_1rw
* cell instance $20373 r0 *1 42.3,120.12
X$20373 185 603 186 644 645 cell_1rw
* cell instance $20374 m0 *1 42.3,122.85
X$20374 185 604 186 644 645 cell_1rw
* cell instance $20375 r0 *1 42.3,122.85
X$20375 185 605 186 644 645 cell_1rw
* cell instance $20376 m0 *1 42.3,125.58
X$20376 185 606 186 644 645 cell_1rw
* cell instance $20377 r0 *1 42.3,125.58
X$20377 185 607 186 644 645 cell_1rw
* cell instance $20378 m0 *1 42.3,128.31
X$20378 185 609 186 644 645 cell_1rw
* cell instance $20379 r0 *1 42.3,128.31
X$20379 185 608 186 644 645 cell_1rw
* cell instance $20380 m0 *1 42.3,131.04
X$20380 185 610 186 644 645 cell_1rw
* cell instance $20381 r0 *1 42.3,131.04
X$20381 185 611 186 644 645 cell_1rw
* cell instance $20382 m0 *1 42.3,133.77
X$20382 185 612 186 644 645 cell_1rw
* cell instance $20383 r0 *1 42.3,133.77
X$20383 185 613 186 644 645 cell_1rw
* cell instance $20384 m0 *1 42.3,136.5
X$20384 185 615 186 644 645 cell_1rw
* cell instance $20385 r0 *1 42.3,136.5
X$20385 185 614 186 644 645 cell_1rw
* cell instance $20386 m0 *1 42.3,139.23
X$20386 185 617 186 644 645 cell_1rw
* cell instance $20387 r0 *1 42.3,139.23
X$20387 185 616 186 644 645 cell_1rw
* cell instance $20388 m0 *1 42.3,141.96
X$20388 185 618 186 644 645 cell_1rw
* cell instance $20389 r0 *1 42.3,141.96
X$20389 185 619 186 644 645 cell_1rw
* cell instance $20390 m0 *1 42.3,144.69
X$20390 185 620 186 644 645 cell_1rw
* cell instance $20391 r0 *1 42.3,144.69
X$20391 185 621 186 644 645 cell_1rw
* cell instance $20392 m0 *1 42.3,147.42
X$20392 185 622 186 644 645 cell_1rw
* cell instance $20393 r0 *1 42.3,147.42
X$20393 185 623 186 644 645 cell_1rw
* cell instance $20394 m0 *1 42.3,150.15
X$20394 185 624 186 644 645 cell_1rw
* cell instance $20395 r0 *1 42.3,150.15
X$20395 185 625 186 644 645 cell_1rw
* cell instance $20396 m0 *1 42.3,152.88
X$20396 185 626 186 644 645 cell_1rw
* cell instance $20397 m0 *1 42.3,155.61
X$20397 185 628 186 644 645 cell_1rw
* cell instance $20398 r0 *1 42.3,152.88
X$20398 185 627 186 644 645 cell_1rw
* cell instance $20399 r0 *1 42.3,155.61
X$20399 185 629 186 644 645 cell_1rw
* cell instance $20400 m0 *1 42.3,158.34
X$20400 185 630 186 644 645 cell_1rw
* cell instance $20401 r0 *1 42.3,158.34
X$20401 185 631 186 644 645 cell_1rw
* cell instance $20402 m0 *1 42.3,161.07
X$20402 185 632 186 644 645 cell_1rw
* cell instance $20403 r0 *1 42.3,161.07
X$20403 185 633 186 644 645 cell_1rw
* cell instance $20404 m0 *1 42.3,163.8
X$20404 185 634 186 644 645 cell_1rw
* cell instance $20405 r0 *1 42.3,163.8
X$20405 185 635 186 644 645 cell_1rw
* cell instance $20406 m0 *1 42.3,166.53
X$20406 185 637 186 644 645 cell_1rw
* cell instance $20407 r0 *1 42.3,166.53
X$20407 185 636 186 644 645 cell_1rw
* cell instance $20408 m0 *1 42.3,169.26
X$20408 185 639 186 644 645 cell_1rw
* cell instance $20409 r0 *1 42.3,169.26
X$20409 185 638 186 644 645 cell_1rw
* cell instance $20410 m0 *1 42.3,171.99
X$20410 185 640 186 644 645 cell_1rw
* cell instance $20411 r0 *1 42.3,171.99
X$20411 185 641 186 644 645 cell_1rw
* cell instance $20412 m0 *1 42.3,174.72
X$20412 185 642 186 644 645 cell_1rw
* cell instance $20413 r0 *1 42.3,174.72
X$20413 185 643 186 644 645 cell_1rw
* cell instance $20414 r0 *1 43.005,87.36
X$20414 187 322 188 644 645 cell_1rw
* cell instance $20415 m0 *1 43.005,90.09
X$20415 187 581 188 644 645 cell_1rw
* cell instance $20416 r0 *1 43.005,90.09
X$20416 187 580 188 644 645 cell_1rw
* cell instance $20417 m0 *1 43.005,92.82
X$20417 187 583 188 644 645 cell_1rw
* cell instance $20418 r0 *1 43.005,92.82
X$20418 187 582 188 644 645 cell_1rw
* cell instance $20419 m0 *1 43.005,95.55
X$20419 187 584 188 644 645 cell_1rw
* cell instance $20420 r0 *1 43.005,95.55
X$20420 187 585 188 644 645 cell_1rw
* cell instance $20421 m0 *1 43.005,98.28
X$20421 187 586 188 644 645 cell_1rw
* cell instance $20422 r0 *1 43.005,98.28
X$20422 187 587 188 644 645 cell_1rw
* cell instance $20423 m0 *1 43.005,101.01
X$20423 187 588 188 644 645 cell_1rw
* cell instance $20424 r0 *1 43.005,101.01
X$20424 187 589 188 644 645 cell_1rw
* cell instance $20425 m0 *1 43.005,103.74
X$20425 187 590 188 644 645 cell_1rw
* cell instance $20426 r0 *1 43.005,103.74
X$20426 187 591 188 644 645 cell_1rw
* cell instance $20427 m0 *1 43.005,106.47
X$20427 187 593 188 644 645 cell_1rw
* cell instance $20428 r0 *1 43.005,106.47
X$20428 187 592 188 644 645 cell_1rw
* cell instance $20429 m0 *1 43.005,109.2
X$20429 187 594 188 644 645 cell_1rw
* cell instance $20430 r0 *1 43.005,109.2
X$20430 187 595 188 644 645 cell_1rw
* cell instance $20431 m0 *1 43.005,111.93
X$20431 187 597 188 644 645 cell_1rw
* cell instance $20432 r0 *1 43.005,111.93
X$20432 187 596 188 644 645 cell_1rw
* cell instance $20433 m0 *1 43.005,114.66
X$20433 187 598 188 644 645 cell_1rw
* cell instance $20434 m0 *1 43.005,117.39
X$20434 187 600 188 644 645 cell_1rw
* cell instance $20435 r0 *1 43.005,114.66
X$20435 187 599 188 644 645 cell_1rw
* cell instance $20436 m0 *1 43.005,120.12
X$20436 187 602 188 644 645 cell_1rw
* cell instance $20437 r0 *1 43.005,117.39
X$20437 187 601 188 644 645 cell_1rw
* cell instance $20438 r0 *1 43.005,120.12
X$20438 187 603 188 644 645 cell_1rw
* cell instance $20439 m0 *1 43.005,122.85
X$20439 187 604 188 644 645 cell_1rw
* cell instance $20440 m0 *1 43.005,125.58
X$20440 187 606 188 644 645 cell_1rw
* cell instance $20441 r0 *1 43.005,122.85
X$20441 187 605 188 644 645 cell_1rw
* cell instance $20442 m0 *1 43.005,128.31
X$20442 187 609 188 644 645 cell_1rw
* cell instance $20443 r0 *1 43.005,125.58
X$20443 187 607 188 644 645 cell_1rw
* cell instance $20444 r0 *1 43.005,128.31
X$20444 187 608 188 644 645 cell_1rw
* cell instance $20445 m0 *1 43.005,131.04
X$20445 187 610 188 644 645 cell_1rw
* cell instance $20446 r0 *1 43.005,131.04
X$20446 187 611 188 644 645 cell_1rw
* cell instance $20447 m0 *1 43.005,133.77
X$20447 187 612 188 644 645 cell_1rw
* cell instance $20448 m0 *1 43.005,136.5
X$20448 187 615 188 644 645 cell_1rw
* cell instance $20449 r0 *1 43.005,133.77
X$20449 187 613 188 644 645 cell_1rw
* cell instance $20450 r0 *1 43.005,136.5
X$20450 187 614 188 644 645 cell_1rw
* cell instance $20451 m0 *1 43.005,139.23
X$20451 187 617 188 644 645 cell_1rw
* cell instance $20452 m0 *1 43.005,141.96
X$20452 187 618 188 644 645 cell_1rw
* cell instance $20453 r0 *1 43.005,139.23
X$20453 187 616 188 644 645 cell_1rw
* cell instance $20454 r0 *1 43.005,141.96
X$20454 187 619 188 644 645 cell_1rw
* cell instance $20455 m0 *1 43.005,144.69
X$20455 187 620 188 644 645 cell_1rw
* cell instance $20456 r0 *1 43.005,144.69
X$20456 187 621 188 644 645 cell_1rw
* cell instance $20457 m0 *1 43.005,147.42
X$20457 187 622 188 644 645 cell_1rw
* cell instance $20458 r0 *1 43.005,147.42
X$20458 187 623 188 644 645 cell_1rw
* cell instance $20459 m0 *1 43.005,150.15
X$20459 187 624 188 644 645 cell_1rw
* cell instance $20460 r0 *1 43.005,150.15
X$20460 187 625 188 644 645 cell_1rw
* cell instance $20461 m0 *1 43.005,152.88
X$20461 187 626 188 644 645 cell_1rw
* cell instance $20462 r0 *1 43.005,152.88
X$20462 187 627 188 644 645 cell_1rw
* cell instance $20463 m0 *1 43.005,155.61
X$20463 187 628 188 644 645 cell_1rw
* cell instance $20464 r0 *1 43.005,155.61
X$20464 187 629 188 644 645 cell_1rw
* cell instance $20465 m0 *1 43.005,158.34
X$20465 187 630 188 644 645 cell_1rw
* cell instance $20466 r0 *1 43.005,158.34
X$20466 187 631 188 644 645 cell_1rw
* cell instance $20467 m0 *1 43.005,161.07
X$20467 187 632 188 644 645 cell_1rw
* cell instance $20468 r0 *1 43.005,161.07
X$20468 187 633 188 644 645 cell_1rw
* cell instance $20469 m0 *1 43.005,163.8
X$20469 187 634 188 644 645 cell_1rw
* cell instance $20470 r0 *1 43.005,163.8
X$20470 187 635 188 644 645 cell_1rw
* cell instance $20471 m0 *1 43.005,166.53
X$20471 187 637 188 644 645 cell_1rw
* cell instance $20472 m0 *1 43.005,169.26
X$20472 187 639 188 644 645 cell_1rw
* cell instance $20473 r0 *1 43.005,166.53
X$20473 187 636 188 644 645 cell_1rw
* cell instance $20474 m0 *1 43.005,171.99
X$20474 187 640 188 644 645 cell_1rw
* cell instance $20475 r0 *1 43.005,169.26
X$20475 187 638 188 644 645 cell_1rw
* cell instance $20476 r0 *1 43.005,171.99
X$20476 187 641 188 644 645 cell_1rw
* cell instance $20477 m0 *1 43.005,174.72
X$20477 187 642 188 644 645 cell_1rw
* cell instance $20478 r0 *1 43.005,174.72
X$20478 187 643 188 644 645 cell_1rw
* cell instance $20479 r0 *1 43.71,87.36
X$20479 189 322 190 644 645 cell_1rw
* cell instance $20480 m0 *1 43.71,90.09
X$20480 189 581 190 644 645 cell_1rw
* cell instance $20481 r0 *1 43.71,90.09
X$20481 189 580 190 644 645 cell_1rw
* cell instance $20482 m0 *1 43.71,92.82
X$20482 189 583 190 644 645 cell_1rw
* cell instance $20483 r0 *1 43.71,92.82
X$20483 189 582 190 644 645 cell_1rw
* cell instance $20484 m0 *1 43.71,95.55
X$20484 189 584 190 644 645 cell_1rw
* cell instance $20485 m0 *1 43.71,98.28
X$20485 189 586 190 644 645 cell_1rw
* cell instance $20486 r0 *1 43.71,95.55
X$20486 189 585 190 644 645 cell_1rw
* cell instance $20487 r0 *1 43.71,98.28
X$20487 189 587 190 644 645 cell_1rw
* cell instance $20488 m0 *1 43.71,101.01
X$20488 189 588 190 644 645 cell_1rw
* cell instance $20489 m0 *1 43.71,103.74
X$20489 189 590 190 644 645 cell_1rw
* cell instance $20490 r0 *1 43.71,101.01
X$20490 189 589 190 644 645 cell_1rw
* cell instance $20491 m0 *1 43.71,106.47
X$20491 189 593 190 644 645 cell_1rw
* cell instance $20492 r0 *1 43.71,103.74
X$20492 189 591 190 644 645 cell_1rw
* cell instance $20493 r0 *1 43.71,106.47
X$20493 189 592 190 644 645 cell_1rw
* cell instance $20494 m0 *1 43.71,109.2
X$20494 189 594 190 644 645 cell_1rw
* cell instance $20495 r0 *1 43.71,109.2
X$20495 189 595 190 644 645 cell_1rw
* cell instance $20496 m0 *1 43.71,111.93
X$20496 189 597 190 644 645 cell_1rw
* cell instance $20497 m0 *1 43.71,114.66
X$20497 189 598 190 644 645 cell_1rw
* cell instance $20498 r0 *1 43.71,111.93
X$20498 189 596 190 644 645 cell_1rw
* cell instance $20499 r0 *1 43.71,114.66
X$20499 189 599 190 644 645 cell_1rw
* cell instance $20500 m0 *1 43.71,117.39
X$20500 189 600 190 644 645 cell_1rw
* cell instance $20501 r0 *1 43.71,117.39
X$20501 189 601 190 644 645 cell_1rw
* cell instance $20502 m0 *1 43.71,120.12
X$20502 189 602 190 644 645 cell_1rw
* cell instance $20503 m0 *1 43.71,122.85
X$20503 189 604 190 644 645 cell_1rw
* cell instance $20504 r0 *1 43.71,120.12
X$20504 189 603 190 644 645 cell_1rw
* cell instance $20505 r0 *1 43.71,122.85
X$20505 189 605 190 644 645 cell_1rw
* cell instance $20506 m0 *1 43.71,125.58
X$20506 189 606 190 644 645 cell_1rw
* cell instance $20507 r0 *1 43.71,125.58
X$20507 189 607 190 644 645 cell_1rw
* cell instance $20508 m0 *1 43.71,128.31
X$20508 189 609 190 644 645 cell_1rw
* cell instance $20509 m0 *1 43.71,131.04
X$20509 189 610 190 644 645 cell_1rw
* cell instance $20510 r0 *1 43.71,128.31
X$20510 189 608 190 644 645 cell_1rw
* cell instance $20511 m0 *1 43.71,133.77
X$20511 189 612 190 644 645 cell_1rw
* cell instance $20512 r0 *1 43.71,131.04
X$20512 189 611 190 644 645 cell_1rw
* cell instance $20513 r0 *1 43.71,133.77
X$20513 189 613 190 644 645 cell_1rw
* cell instance $20514 m0 *1 43.71,136.5
X$20514 189 615 190 644 645 cell_1rw
* cell instance $20515 r0 *1 43.71,136.5
X$20515 189 614 190 644 645 cell_1rw
* cell instance $20516 m0 *1 43.71,139.23
X$20516 189 617 190 644 645 cell_1rw
* cell instance $20517 r0 *1 43.71,139.23
X$20517 189 616 190 644 645 cell_1rw
* cell instance $20518 m0 *1 43.71,141.96
X$20518 189 618 190 644 645 cell_1rw
* cell instance $20519 r0 *1 43.71,141.96
X$20519 189 619 190 644 645 cell_1rw
* cell instance $20520 m0 *1 43.71,144.69
X$20520 189 620 190 644 645 cell_1rw
* cell instance $20521 r0 *1 43.71,144.69
X$20521 189 621 190 644 645 cell_1rw
* cell instance $20522 m0 *1 43.71,147.42
X$20522 189 622 190 644 645 cell_1rw
* cell instance $20523 r0 *1 43.71,147.42
X$20523 189 623 190 644 645 cell_1rw
* cell instance $20524 m0 *1 43.71,150.15
X$20524 189 624 190 644 645 cell_1rw
* cell instance $20525 m0 *1 43.71,152.88
X$20525 189 626 190 644 645 cell_1rw
* cell instance $20526 r0 *1 43.71,150.15
X$20526 189 625 190 644 645 cell_1rw
* cell instance $20527 r0 *1 43.71,152.88
X$20527 189 627 190 644 645 cell_1rw
* cell instance $20528 m0 *1 43.71,155.61
X$20528 189 628 190 644 645 cell_1rw
* cell instance $20529 r0 *1 43.71,155.61
X$20529 189 629 190 644 645 cell_1rw
* cell instance $20530 m0 *1 43.71,158.34
X$20530 189 630 190 644 645 cell_1rw
* cell instance $20531 m0 *1 43.71,161.07
X$20531 189 632 190 644 645 cell_1rw
* cell instance $20532 r0 *1 43.71,158.34
X$20532 189 631 190 644 645 cell_1rw
* cell instance $20533 r0 *1 43.71,161.07
X$20533 189 633 190 644 645 cell_1rw
* cell instance $20534 m0 *1 43.71,163.8
X$20534 189 634 190 644 645 cell_1rw
* cell instance $20535 r0 *1 43.71,163.8
X$20535 189 635 190 644 645 cell_1rw
* cell instance $20536 m0 *1 43.71,166.53
X$20536 189 637 190 644 645 cell_1rw
* cell instance $20537 r0 *1 43.71,166.53
X$20537 189 636 190 644 645 cell_1rw
* cell instance $20538 m0 *1 43.71,169.26
X$20538 189 639 190 644 645 cell_1rw
* cell instance $20539 r0 *1 43.71,169.26
X$20539 189 638 190 644 645 cell_1rw
* cell instance $20540 m0 *1 43.71,171.99
X$20540 189 640 190 644 645 cell_1rw
* cell instance $20541 r0 *1 43.71,171.99
X$20541 189 641 190 644 645 cell_1rw
* cell instance $20542 m0 *1 43.71,174.72
X$20542 189 642 190 644 645 cell_1rw
* cell instance $20543 r0 *1 43.71,174.72
X$20543 189 643 190 644 645 cell_1rw
* cell instance $20544 r0 *1 44.415,87.36
X$20544 191 322 192 644 645 cell_1rw
* cell instance $20545 m0 *1 44.415,90.09
X$20545 191 581 192 644 645 cell_1rw
* cell instance $20546 m0 *1 44.415,92.82
X$20546 191 583 192 644 645 cell_1rw
* cell instance $20547 r0 *1 44.415,90.09
X$20547 191 580 192 644 645 cell_1rw
* cell instance $20548 r0 *1 44.415,92.82
X$20548 191 582 192 644 645 cell_1rw
* cell instance $20549 m0 *1 44.415,95.55
X$20549 191 584 192 644 645 cell_1rw
* cell instance $20550 r0 *1 44.415,95.55
X$20550 191 585 192 644 645 cell_1rw
* cell instance $20551 m0 *1 44.415,98.28
X$20551 191 586 192 644 645 cell_1rw
* cell instance $20552 r0 *1 44.415,98.28
X$20552 191 587 192 644 645 cell_1rw
* cell instance $20553 m0 *1 44.415,101.01
X$20553 191 588 192 644 645 cell_1rw
* cell instance $20554 r0 *1 44.415,101.01
X$20554 191 589 192 644 645 cell_1rw
* cell instance $20555 m0 *1 44.415,103.74
X$20555 191 590 192 644 645 cell_1rw
* cell instance $20556 r0 *1 44.415,103.74
X$20556 191 591 192 644 645 cell_1rw
* cell instance $20557 m0 *1 44.415,106.47
X$20557 191 593 192 644 645 cell_1rw
* cell instance $20558 r0 *1 44.415,106.47
X$20558 191 592 192 644 645 cell_1rw
* cell instance $20559 m0 *1 44.415,109.2
X$20559 191 594 192 644 645 cell_1rw
* cell instance $20560 m0 *1 44.415,111.93
X$20560 191 597 192 644 645 cell_1rw
* cell instance $20561 r0 *1 44.415,109.2
X$20561 191 595 192 644 645 cell_1rw
* cell instance $20562 r0 *1 44.415,111.93
X$20562 191 596 192 644 645 cell_1rw
* cell instance $20563 m0 *1 44.415,114.66
X$20563 191 598 192 644 645 cell_1rw
* cell instance $20564 r0 *1 44.415,114.66
X$20564 191 599 192 644 645 cell_1rw
* cell instance $20565 m0 *1 44.415,117.39
X$20565 191 600 192 644 645 cell_1rw
* cell instance $20566 m0 *1 44.415,120.12
X$20566 191 602 192 644 645 cell_1rw
* cell instance $20567 r0 *1 44.415,117.39
X$20567 191 601 192 644 645 cell_1rw
* cell instance $20568 m0 *1 44.415,122.85
X$20568 191 604 192 644 645 cell_1rw
* cell instance $20569 r0 *1 44.415,120.12
X$20569 191 603 192 644 645 cell_1rw
* cell instance $20570 r0 *1 44.415,122.85
X$20570 191 605 192 644 645 cell_1rw
* cell instance $20571 m0 *1 44.415,125.58
X$20571 191 606 192 644 645 cell_1rw
* cell instance $20572 m0 *1 44.415,128.31
X$20572 191 609 192 644 645 cell_1rw
* cell instance $20573 r0 *1 44.415,125.58
X$20573 191 607 192 644 645 cell_1rw
* cell instance $20574 r0 *1 44.415,128.31
X$20574 191 608 192 644 645 cell_1rw
* cell instance $20575 m0 *1 44.415,131.04
X$20575 191 610 192 644 645 cell_1rw
* cell instance $20576 m0 *1 44.415,133.77
X$20576 191 612 192 644 645 cell_1rw
* cell instance $20577 r0 *1 44.415,131.04
X$20577 191 611 192 644 645 cell_1rw
* cell instance $20578 r0 *1 44.415,133.77
X$20578 191 613 192 644 645 cell_1rw
* cell instance $20579 m0 *1 44.415,136.5
X$20579 191 615 192 644 645 cell_1rw
* cell instance $20580 r0 *1 44.415,136.5
X$20580 191 614 192 644 645 cell_1rw
* cell instance $20581 m0 *1 44.415,139.23
X$20581 191 617 192 644 645 cell_1rw
* cell instance $20582 r0 *1 44.415,139.23
X$20582 191 616 192 644 645 cell_1rw
* cell instance $20583 m0 *1 44.415,141.96
X$20583 191 618 192 644 645 cell_1rw
* cell instance $20584 r0 *1 44.415,141.96
X$20584 191 619 192 644 645 cell_1rw
* cell instance $20585 m0 *1 44.415,144.69
X$20585 191 620 192 644 645 cell_1rw
* cell instance $20586 r0 *1 44.415,144.69
X$20586 191 621 192 644 645 cell_1rw
* cell instance $20587 m0 *1 44.415,147.42
X$20587 191 622 192 644 645 cell_1rw
* cell instance $20588 m0 *1 44.415,150.15
X$20588 191 624 192 644 645 cell_1rw
* cell instance $20589 r0 *1 44.415,147.42
X$20589 191 623 192 644 645 cell_1rw
* cell instance $20590 r0 *1 44.415,150.15
X$20590 191 625 192 644 645 cell_1rw
* cell instance $20591 m0 *1 44.415,152.88
X$20591 191 626 192 644 645 cell_1rw
* cell instance $20592 r0 *1 44.415,152.88
X$20592 191 627 192 644 645 cell_1rw
* cell instance $20593 m0 *1 44.415,155.61
X$20593 191 628 192 644 645 cell_1rw
* cell instance $20594 r0 *1 44.415,155.61
X$20594 191 629 192 644 645 cell_1rw
* cell instance $20595 m0 *1 44.415,158.34
X$20595 191 630 192 644 645 cell_1rw
* cell instance $20596 m0 *1 44.415,161.07
X$20596 191 632 192 644 645 cell_1rw
* cell instance $20597 r0 *1 44.415,158.34
X$20597 191 631 192 644 645 cell_1rw
* cell instance $20598 r0 *1 44.415,161.07
X$20598 191 633 192 644 645 cell_1rw
* cell instance $20599 m0 *1 44.415,163.8
X$20599 191 634 192 644 645 cell_1rw
* cell instance $20600 r0 *1 44.415,163.8
X$20600 191 635 192 644 645 cell_1rw
* cell instance $20601 m0 *1 44.415,166.53
X$20601 191 637 192 644 645 cell_1rw
* cell instance $20602 r0 *1 44.415,166.53
X$20602 191 636 192 644 645 cell_1rw
* cell instance $20603 m0 *1 44.415,169.26
X$20603 191 639 192 644 645 cell_1rw
* cell instance $20604 r0 *1 44.415,169.26
X$20604 191 638 192 644 645 cell_1rw
* cell instance $20605 m0 *1 44.415,171.99
X$20605 191 640 192 644 645 cell_1rw
* cell instance $20606 r0 *1 44.415,171.99
X$20606 191 641 192 644 645 cell_1rw
* cell instance $20607 m0 *1 44.415,174.72
X$20607 191 642 192 644 645 cell_1rw
* cell instance $20608 r0 *1 44.415,174.72
X$20608 191 643 192 644 645 cell_1rw
* cell instance $20609 r0 *1 45.12,87.36
X$20609 193 322 194 644 645 cell_1rw
* cell instance $20610 m0 *1 45.12,90.09
X$20610 193 581 194 644 645 cell_1rw
* cell instance $20611 r0 *1 45.12,90.09
X$20611 193 580 194 644 645 cell_1rw
* cell instance $20612 m0 *1 45.12,92.82
X$20612 193 583 194 644 645 cell_1rw
* cell instance $20613 r0 *1 45.12,92.82
X$20613 193 582 194 644 645 cell_1rw
* cell instance $20614 m0 *1 45.12,95.55
X$20614 193 584 194 644 645 cell_1rw
* cell instance $20615 r0 *1 45.12,95.55
X$20615 193 585 194 644 645 cell_1rw
* cell instance $20616 m0 *1 45.12,98.28
X$20616 193 586 194 644 645 cell_1rw
* cell instance $20617 r0 *1 45.12,98.28
X$20617 193 587 194 644 645 cell_1rw
* cell instance $20618 m0 *1 45.12,101.01
X$20618 193 588 194 644 645 cell_1rw
* cell instance $20619 r0 *1 45.12,101.01
X$20619 193 589 194 644 645 cell_1rw
* cell instance $20620 m0 *1 45.12,103.74
X$20620 193 590 194 644 645 cell_1rw
* cell instance $20621 r0 *1 45.12,103.74
X$20621 193 591 194 644 645 cell_1rw
* cell instance $20622 m0 *1 45.12,106.47
X$20622 193 593 194 644 645 cell_1rw
* cell instance $20623 r0 *1 45.12,106.47
X$20623 193 592 194 644 645 cell_1rw
* cell instance $20624 m0 *1 45.12,109.2
X$20624 193 594 194 644 645 cell_1rw
* cell instance $20625 r0 *1 45.12,109.2
X$20625 193 595 194 644 645 cell_1rw
* cell instance $20626 m0 *1 45.12,111.93
X$20626 193 597 194 644 645 cell_1rw
* cell instance $20627 r0 *1 45.12,111.93
X$20627 193 596 194 644 645 cell_1rw
* cell instance $20628 m0 *1 45.12,114.66
X$20628 193 598 194 644 645 cell_1rw
* cell instance $20629 r0 *1 45.12,114.66
X$20629 193 599 194 644 645 cell_1rw
* cell instance $20630 m0 *1 45.12,117.39
X$20630 193 600 194 644 645 cell_1rw
* cell instance $20631 r0 *1 45.12,117.39
X$20631 193 601 194 644 645 cell_1rw
* cell instance $20632 m0 *1 45.12,120.12
X$20632 193 602 194 644 645 cell_1rw
* cell instance $20633 r0 *1 45.12,120.12
X$20633 193 603 194 644 645 cell_1rw
* cell instance $20634 m0 *1 45.12,122.85
X$20634 193 604 194 644 645 cell_1rw
* cell instance $20635 r0 *1 45.12,122.85
X$20635 193 605 194 644 645 cell_1rw
* cell instance $20636 m0 *1 45.12,125.58
X$20636 193 606 194 644 645 cell_1rw
* cell instance $20637 r0 *1 45.12,125.58
X$20637 193 607 194 644 645 cell_1rw
* cell instance $20638 m0 *1 45.12,128.31
X$20638 193 609 194 644 645 cell_1rw
* cell instance $20639 m0 *1 45.12,131.04
X$20639 193 610 194 644 645 cell_1rw
* cell instance $20640 r0 *1 45.12,128.31
X$20640 193 608 194 644 645 cell_1rw
* cell instance $20641 m0 *1 45.12,133.77
X$20641 193 612 194 644 645 cell_1rw
* cell instance $20642 r0 *1 45.12,131.04
X$20642 193 611 194 644 645 cell_1rw
* cell instance $20643 r0 *1 45.12,133.77
X$20643 193 613 194 644 645 cell_1rw
* cell instance $20644 m0 *1 45.12,136.5
X$20644 193 615 194 644 645 cell_1rw
* cell instance $20645 r0 *1 45.12,136.5
X$20645 193 614 194 644 645 cell_1rw
* cell instance $20646 m0 *1 45.12,139.23
X$20646 193 617 194 644 645 cell_1rw
* cell instance $20647 r0 *1 45.12,139.23
X$20647 193 616 194 644 645 cell_1rw
* cell instance $20648 m0 *1 45.12,141.96
X$20648 193 618 194 644 645 cell_1rw
* cell instance $20649 m0 *1 45.12,144.69
X$20649 193 620 194 644 645 cell_1rw
* cell instance $20650 r0 *1 45.12,141.96
X$20650 193 619 194 644 645 cell_1rw
* cell instance $20651 r0 *1 45.12,144.69
X$20651 193 621 194 644 645 cell_1rw
* cell instance $20652 m0 *1 45.12,147.42
X$20652 193 622 194 644 645 cell_1rw
* cell instance $20653 r0 *1 45.12,147.42
X$20653 193 623 194 644 645 cell_1rw
* cell instance $20654 m0 *1 45.12,150.15
X$20654 193 624 194 644 645 cell_1rw
* cell instance $20655 r0 *1 45.12,150.15
X$20655 193 625 194 644 645 cell_1rw
* cell instance $20656 m0 *1 45.12,152.88
X$20656 193 626 194 644 645 cell_1rw
* cell instance $20657 m0 *1 45.12,155.61
X$20657 193 628 194 644 645 cell_1rw
* cell instance $20658 r0 *1 45.12,152.88
X$20658 193 627 194 644 645 cell_1rw
* cell instance $20659 r0 *1 45.12,155.61
X$20659 193 629 194 644 645 cell_1rw
* cell instance $20660 m0 *1 45.12,158.34
X$20660 193 630 194 644 645 cell_1rw
* cell instance $20661 r0 *1 45.12,158.34
X$20661 193 631 194 644 645 cell_1rw
* cell instance $20662 m0 *1 45.12,161.07
X$20662 193 632 194 644 645 cell_1rw
* cell instance $20663 r0 *1 45.12,161.07
X$20663 193 633 194 644 645 cell_1rw
* cell instance $20664 m0 *1 45.12,163.8
X$20664 193 634 194 644 645 cell_1rw
* cell instance $20665 r0 *1 45.12,163.8
X$20665 193 635 194 644 645 cell_1rw
* cell instance $20666 m0 *1 45.12,166.53
X$20666 193 637 194 644 645 cell_1rw
* cell instance $20667 r0 *1 45.12,166.53
X$20667 193 636 194 644 645 cell_1rw
* cell instance $20668 m0 *1 45.12,169.26
X$20668 193 639 194 644 645 cell_1rw
* cell instance $20669 m0 *1 45.12,171.99
X$20669 193 640 194 644 645 cell_1rw
* cell instance $20670 r0 *1 45.12,169.26
X$20670 193 638 194 644 645 cell_1rw
* cell instance $20671 r0 *1 45.12,171.99
X$20671 193 641 194 644 645 cell_1rw
* cell instance $20672 m0 *1 45.12,174.72
X$20672 193 642 194 644 645 cell_1rw
* cell instance $20673 r0 *1 45.12,174.72
X$20673 193 643 194 644 645 cell_1rw
* cell instance $20674 m0 *1 45.825,90.09
X$20674 195 581 196 644 645 cell_1rw
* cell instance $20675 r0 *1 45.825,87.36
X$20675 195 322 196 644 645 cell_1rw
* cell instance $20676 r0 *1 45.825,90.09
X$20676 195 580 196 644 645 cell_1rw
* cell instance $20677 m0 *1 45.825,92.82
X$20677 195 583 196 644 645 cell_1rw
* cell instance $20678 r0 *1 45.825,92.82
X$20678 195 582 196 644 645 cell_1rw
* cell instance $20679 m0 *1 45.825,95.55
X$20679 195 584 196 644 645 cell_1rw
* cell instance $20680 m0 *1 45.825,98.28
X$20680 195 586 196 644 645 cell_1rw
* cell instance $20681 r0 *1 45.825,95.55
X$20681 195 585 196 644 645 cell_1rw
* cell instance $20682 r0 *1 45.825,98.28
X$20682 195 587 196 644 645 cell_1rw
* cell instance $20683 m0 *1 45.825,101.01
X$20683 195 588 196 644 645 cell_1rw
* cell instance $20684 r0 *1 45.825,101.01
X$20684 195 589 196 644 645 cell_1rw
* cell instance $20685 m0 *1 45.825,103.74
X$20685 195 590 196 644 645 cell_1rw
* cell instance $20686 r0 *1 45.825,103.74
X$20686 195 591 196 644 645 cell_1rw
* cell instance $20687 m0 *1 45.825,106.47
X$20687 195 593 196 644 645 cell_1rw
* cell instance $20688 r0 *1 45.825,106.47
X$20688 195 592 196 644 645 cell_1rw
* cell instance $20689 m0 *1 45.825,109.2
X$20689 195 594 196 644 645 cell_1rw
* cell instance $20690 r0 *1 45.825,109.2
X$20690 195 595 196 644 645 cell_1rw
* cell instance $20691 m0 *1 45.825,111.93
X$20691 195 597 196 644 645 cell_1rw
* cell instance $20692 r0 *1 45.825,111.93
X$20692 195 596 196 644 645 cell_1rw
* cell instance $20693 m0 *1 45.825,114.66
X$20693 195 598 196 644 645 cell_1rw
* cell instance $20694 r0 *1 45.825,114.66
X$20694 195 599 196 644 645 cell_1rw
* cell instance $20695 m0 *1 45.825,117.39
X$20695 195 600 196 644 645 cell_1rw
* cell instance $20696 m0 *1 45.825,120.12
X$20696 195 602 196 644 645 cell_1rw
* cell instance $20697 r0 *1 45.825,117.39
X$20697 195 601 196 644 645 cell_1rw
* cell instance $20698 m0 *1 45.825,122.85
X$20698 195 604 196 644 645 cell_1rw
* cell instance $20699 r0 *1 45.825,120.12
X$20699 195 603 196 644 645 cell_1rw
* cell instance $20700 m0 *1 45.825,125.58
X$20700 195 606 196 644 645 cell_1rw
* cell instance $20701 r0 *1 45.825,122.85
X$20701 195 605 196 644 645 cell_1rw
* cell instance $20702 m0 *1 45.825,128.31
X$20702 195 609 196 644 645 cell_1rw
* cell instance $20703 r0 *1 45.825,125.58
X$20703 195 607 196 644 645 cell_1rw
* cell instance $20704 r0 *1 45.825,128.31
X$20704 195 608 196 644 645 cell_1rw
* cell instance $20705 m0 *1 45.825,131.04
X$20705 195 610 196 644 645 cell_1rw
* cell instance $20706 m0 *1 45.825,133.77
X$20706 195 612 196 644 645 cell_1rw
* cell instance $20707 r0 *1 45.825,131.04
X$20707 195 611 196 644 645 cell_1rw
* cell instance $20708 r0 *1 45.825,133.77
X$20708 195 613 196 644 645 cell_1rw
* cell instance $20709 m0 *1 45.825,136.5
X$20709 195 615 196 644 645 cell_1rw
* cell instance $20710 r0 *1 45.825,136.5
X$20710 195 614 196 644 645 cell_1rw
* cell instance $20711 m0 *1 45.825,139.23
X$20711 195 617 196 644 645 cell_1rw
* cell instance $20712 r0 *1 45.825,139.23
X$20712 195 616 196 644 645 cell_1rw
* cell instance $20713 m0 *1 45.825,141.96
X$20713 195 618 196 644 645 cell_1rw
* cell instance $20714 r0 *1 45.825,141.96
X$20714 195 619 196 644 645 cell_1rw
* cell instance $20715 m0 *1 45.825,144.69
X$20715 195 620 196 644 645 cell_1rw
* cell instance $20716 r0 *1 45.825,144.69
X$20716 195 621 196 644 645 cell_1rw
* cell instance $20717 m0 *1 45.825,147.42
X$20717 195 622 196 644 645 cell_1rw
* cell instance $20718 r0 *1 45.825,147.42
X$20718 195 623 196 644 645 cell_1rw
* cell instance $20719 m0 *1 45.825,150.15
X$20719 195 624 196 644 645 cell_1rw
* cell instance $20720 r0 *1 45.825,150.15
X$20720 195 625 196 644 645 cell_1rw
* cell instance $20721 m0 *1 45.825,152.88
X$20721 195 626 196 644 645 cell_1rw
* cell instance $20722 r0 *1 45.825,152.88
X$20722 195 627 196 644 645 cell_1rw
* cell instance $20723 m0 *1 45.825,155.61
X$20723 195 628 196 644 645 cell_1rw
* cell instance $20724 r0 *1 45.825,155.61
X$20724 195 629 196 644 645 cell_1rw
* cell instance $20725 m0 *1 45.825,158.34
X$20725 195 630 196 644 645 cell_1rw
* cell instance $20726 r0 *1 45.825,158.34
X$20726 195 631 196 644 645 cell_1rw
* cell instance $20727 m0 *1 45.825,161.07
X$20727 195 632 196 644 645 cell_1rw
* cell instance $20728 r0 *1 45.825,161.07
X$20728 195 633 196 644 645 cell_1rw
* cell instance $20729 m0 *1 45.825,163.8
X$20729 195 634 196 644 645 cell_1rw
* cell instance $20730 r0 *1 45.825,163.8
X$20730 195 635 196 644 645 cell_1rw
* cell instance $20731 m0 *1 45.825,166.53
X$20731 195 637 196 644 645 cell_1rw
* cell instance $20732 r0 *1 45.825,166.53
X$20732 195 636 196 644 645 cell_1rw
* cell instance $20733 m0 *1 45.825,169.26
X$20733 195 639 196 644 645 cell_1rw
* cell instance $20734 m0 *1 45.825,171.99
X$20734 195 640 196 644 645 cell_1rw
* cell instance $20735 r0 *1 45.825,169.26
X$20735 195 638 196 644 645 cell_1rw
* cell instance $20736 m0 *1 45.825,174.72
X$20736 195 642 196 644 645 cell_1rw
* cell instance $20737 r0 *1 45.825,171.99
X$20737 195 641 196 644 645 cell_1rw
* cell instance $20738 r0 *1 45.825,174.72
X$20738 195 643 196 644 645 cell_1rw
* cell instance $20739 r0 *1 46.53,87.36
X$20739 197 322 198 644 645 cell_1rw
* cell instance $20740 m0 *1 46.53,90.09
X$20740 197 581 198 644 645 cell_1rw
* cell instance $20741 m0 *1 46.53,92.82
X$20741 197 583 198 644 645 cell_1rw
* cell instance $20742 r0 *1 46.53,90.09
X$20742 197 580 198 644 645 cell_1rw
* cell instance $20743 r0 *1 46.53,92.82
X$20743 197 582 198 644 645 cell_1rw
* cell instance $20744 m0 *1 46.53,95.55
X$20744 197 584 198 644 645 cell_1rw
* cell instance $20745 r0 *1 46.53,95.55
X$20745 197 585 198 644 645 cell_1rw
* cell instance $20746 m0 *1 46.53,98.28
X$20746 197 586 198 644 645 cell_1rw
* cell instance $20747 r0 *1 46.53,98.28
X$20747 197 587 198 644 645 cell_1rw
* cell instance $20748 m0 *1 46.53,101.01
X$20748 197 588 198 644 645 cell_1rw
* cell instance $20749 r0 *1 46.53,101.01
X$20749 197 589 198 644 645 cell_1rw
* cell instance $20750 m0 *1 46.53,103.74
X$20750 197 590 198 644 645 cell_1rw
* cell instance $20751 r0 *1 46.53,103.74
X$20751 197 591 198 644 645 cell_1rw
* cell instance $20752 m0 *1 46.53,106.47
X$20752 197 593 198 644 645 cell_1rw
* cell instance $20753 r0 *1 46.53,106.47
X$20753 197 592 198 644 645 cell_1rw
* cell instance $20754 m0 *1 46.53,109.2
X$20754 197 594 198 644 645 cell_1rw
* cell instance $20755 r0 *1 46.53,109.2
X$20755 197 595 198 644 645 cell_1rw
* cell instance $20756 m0 *1 46.53,111.93
X$20756 197 597 198 644 645 cell_1rw
* cell instance $20757 r0 *1 46.53,111.93
X$20757 197 596 198 644 645 cell_1rw
* cell instance $20758 m0 *1 46.53,114.66
X$20758 197 598 198 644 645 cell_1rw
* cell instance $20759 m0 *1 46.53,117.39
X$20759 197 600 198 644 645 cell_1rw
* cell instance $20760 r0 *1 46.53,114.66
X$20760 197 599 198 644 645 cell_1rw
* cell instance $20761 r0 *1 46.53,117.39
X$20761 197 601 198 644 645 cell_1rw
* cell instance $20762 m0 *1 46.53,120.12
X$20762 197 602 198 644 645 cell_1rw
* cell instance $20763 r0 *1 46.53,120.12
X$20763 197 603 198 644 645 cell_1rw
* cell instance $20764 m0 *1 46.53,122.85
X$20764 197 604 198 644 645 cell_1rw
* cell instance $20765 m0 *1 46.53,125.58
X$20765 197 606 198 644 645 cell_1rw
* cell instance $20766 r0 *1 46.53,122.85
X$20766 197 605 198 644 645 cell_1rw
* cell instance $20767 r0 *1 46.53,125.58
X$20767 197 607 198 644 645 cell_1rw
* cell instance $20768 m0 *1 46.53,128.31
X$20768 197 609 198 644 645 cell_1rw
* cell instance $20769 r0 *1 46.53,128.31
X$20769 197 608 198 644 645 cell_1rw
* cell instance $20770 m0 *1 46.53,131.04
X$20770 197 610 198 644 645 cell_1rw
* cell instance $20771 r0 *1 46.53,131.04
X$20771 197 611 198 644 645 cell_1rw
* cell instance $20772 m0 *1 46.53,133.77
X$20772 197 612 198 644 645 cell_1rw
* cell instance $20773 r0 *1 46.53,133.77
X$20773 197 613 198 644 645 cell_1rw
* cell instance $20774 m0 *1 46.53,136.5
X$20774 197 615 198 644 645 cell_1rw
* cell instance $20775 r0 *1 46.53,136.5
X$20775 197 614 198 644 645 cell_1rw
* cell instance $20776 m0 *1 46.53,139.23
X$20776 197 617 198 644 645 cell_1rw
* cell instance $20777 m0 *1 46.53,141.96
X$20777 197 618 198 644 645 cell_1rw
* cell instance $20778 r0 *1 46.53,139.23
X$20778 197 616 198 644 645 cell_1rw
* cell instance $20779 r0 *1 46.53,141.96
X$20779 197 619 198 644 645 cell_1rw
* cell instance $20780 m0 *1 46.53,144.69
X$20780 197 620 198 644 645 cell_1rw
* cell instance $20781 r0 *1 46.53,144.69
X$20781 197 621 198 644 645 cell_1rw
* cell instance $20782 m0 *1 46.53,147.42
X$20782 197 622 198 644 645 cell_1rw
* cell instance $20783 r0 *1 46.53,147.42
X$20783 197 623 198 644 645 cell_1rw
* cell instance $20784 m0 *1 46.53,150.15
X$20784 197 624 198 644 645 cell_1rw
* cell instance $20785 r0 *1 46.53,150.15
X$20785 197 625 198 644 645 cell_1rw
* cell instance $20786 m0 *1 46.53,152.88
X$20786 197 626 198 644 645 cell_1rw
* cell instance $20787 r0 *1 46.53,152.88
X$20787 197 627 198 644 645 cell_1rw
* cell instance $20788 m0 *1 46.53,155.61
X$20788 197 628 198 644 645 cell_1rw
* cell instance $20789 r0 *1 46.53,155.61
X$20789 197 629 198 644 645 cell_1rw
* cell instance $20790 m0 *1 46.53,158.34
X$20790 197 630 198 644 645 cell_1rw
* cell instance $20791 m0 *1 46.53,161.07
X$20791 197 632 198 644 645 cell_1rw
* cell instance $20792 r0 *1 46.53,158.34
X$20792 197 631 198 644 645 cell_1rw
* cell instance $20793 r0 *1 46.53,161.07
X$20793 197 633 198 644 645 cell_1rw
* cell instance $20794 m0 *1 46.53,163.8
X$20794 197 634 198 644 645 cell_1rw
* cell instance $20795 r0 *1 46.53,163.8
X$20795 197 635 198 644 645 cell_1rw
* cell instance $20796 m0 *1 46.53,166.53
X$20796 197 637 198 644 645 cell_1rw
* cell instance $20797 r0 *1 46.53,166.53
X$20797 197 636 198 644 645 cell_1rw
* cell instance $20798 m0 *1 46.53,169.26
X$20798 197 639 198 644 645 cell_1rw
* cell instance $20799 m0 *1 46.53,171.99
X$20799 197 640 198 644 645 cell_1rw
* cell instance $20800 r0 *1 46.53,169.26
X$20800 197 638 198 644 645 cell_1rw
* cell instance $20801 r0 *1 46.53,171.99
X$20801 197 641 198 644 645 cell_1rw
* cell instance $20802 m0 *1 46.53,174.72
X$20802 197 642 198 644 645 cell_1rw
* cell instance $20803 r0 *1 46.53,174.72
X$20803 197 643 198 644 645 cell_1rw
* cell instance $20804 r0 *1 47.235,87.36
X$20804 199 322 200 644 645 cell_1rw
* cell instance $20805 m0 *1 47.235,90.09
X$20805 199 581 200 644 645 cell_1rw
* cell instance $20806 r0 *1 47.235,90.09
X$20806 199 580 200 644 645 cell_1rw
* cell instance $20807 m0 *1 47.235,92.82
X$20807 199 583 200 644 645 cell_1rw
* cell instance $20808 r0 *1 47.235,92.82
X$20808 199 582 200 644 645 cell_1rw
* cell instance $20809 m0 *1 47.235,95.55
X$20809 199 584 200 644 645 cell_1rw
* cell instance $20810 m0 *1 47.235,98.28
X$20810 199 586 200 644 645 cell_1rw
* cell instance $20811 r0 *1 47.235,95.55
X$20811 199 585 200 644 645 cell_1rw
* cell instance $20812 r0 *1 47.235,98.28
X$20812 199 587 200 644 645 cell_1rw
* cell instance $20813 m0 *1 47.235,101.01
X$20813 199 588 200 644 645 cell_1rw
* cell instance $20814 r0 *1 47.235,101.01
X$20814 199 589 200 644 645 cell_1rw
* cell instance $20815 m0 *1 47.235,103.74
X$20815 199 590 200 644 645 cell_1rw
* cell instance $20816 r0 *1 47.235,103.74
X$20816 199 591 200 644 645 cell_1rw
* cell instance $20817 m0 *1 47.235,106.47
X$20817 199 593 200 644 645 cell_1rw
* cell instance $20818 m0 *1 47.235,109.2
X$20818 199 594 200 644 645 cell_1rw
* cell instance $20819 r0 *1 47.235,106.47
X$20819 199 592 200 644 645 cell_1rw
* cell instance $20820 r0 *1 47.235,109.2
X$20820 199 595 200 644 645 cell_1rw
* cell instance $20821 m0 *1 47.235,111.93
X$20821 199 597 200 644 645 cell_1rw
* cell instance $20822 m0 *1 47.235,114.66
X$20822 199 598 200 644 645 cell_1rw
* cell instance $20823 r0 *1 47.235,111.93
X$20823 199 596 200 644 645 cell_1rw
* cell instance $20824 r0 *1 47.235,114.66
X$20824 199 599 200 644 645 cell_1rw
* cell instance $20825 m0 *1 47.235,117.39
X$20825 199 600 200 644 645 cell_1rw
* cell instance $20826 m0 *1 47.235,120.12
X$20826 199 602 200 644 645 cell_1rw
* cell instance $20827 r0 *1 47.235,117.39
X$20827 199 601 200 644 645 cell_1rw
* cell instance $20828 r0 *1 47.235,120.12
X$20828 199 603 200 644 645 cell_1rw
* cell instance $20829 m0 *1 47.235,122.85
X$20829 199 604 200 644 645 cell_1rw
* cell instance $20830 r0 *1 47.235,122.85
X$20830 199 605 200 644 645 cell_1rw
* cell instance $20831 m0 *1 47.235,125.58
X$20831 199 606 200 644 645 cell_1rw
* cell instance $20832 r0 *1 47.235,125.58
X$20832 199 607 200 644 645 cell_1rw
* cell instance $20833 m0 *1 47.235,128.31
X$20833 199 609 200 644 645 cell_1rw
* cell instance $20834 r0 *1 47.235,128.31
X$20834 199 608 200 644 645 cell_1rw
* cell instance $20835 m0 *1 47.235,131.04
X$20835 199 610 200 644 645 cell_1rw
* cell instance $20836 m0 *1 47.235,133.77
X$20836 199 612 200 644 645 cell_1rw
* cell instance $20837 r0 *1 47.235,131.04
X$20837 199 611 200 644 645 cell_1rw
* cell instance $20838 r0 *1 47.235,133.77
X$20838 199 613 200 644 645 cell_1rw
* cell instance $20839 m0 *1 47.235,136.5
X$20839 199 615 200 644 645 cell_1rw
* cell instance $20840 r0 *1 47.235,136.5
X$20840 199 614 200 644 645 cell_1rw
* cell instance $20841 m0 *1 47.235,139.23
X$20841 199 617 200 644 645 cell_1rw
* cell instance $20842 r0 *1 47.235,139.23
X$20842 199 616 200 644 645 cell_1rw
* cell instance $20843 m0 *1 47.235,141.96
X$20843 199 618 200 644 645 cell_1rw
* cell instance $20844 r0 *1 47.235,141.96
X$20844 199 619 200 644 645 cell_1rw
* cell instance $20845 m0 *1 47.235,144.69
X$20845 199 620 200 644 645 cell_1rw
* cell instance $20846 r0 *1 47.235,144.69
X$20846 199 621 200 644 645 cell_1rw
* cell instance $20847 m0 *1 47.235,147.42
X$20847 199 622 200 644 645 cell_1rw
* cell instance $20848 r0 *1 47.235,147.42
X$20848 199 623 200 644 645 cell_1rw
* cell instance $20849 m0 *1 47.235,150.15
X$20849 199 624 200 644 645 cell_1rw
* cell instance $20850 r0 *1 47.235,150.15
X$20850 199 625 200 644 645 cell_1rw
* cell instance $20851 m0 *1 47.235,152.88
X$20851 199 626 200 644 645 cell_1rw
* cell instance $20852 r0 *1 47.235,152.88
X$20852 199 627 200 644 645 cell_1rw
* cell instance $20853 m0 *1 47.235,155.61
X$20853 199 628 200 644 645 cell_1rw
* cell instance $20854 r0 *1 47.235,155.61
X$20854 199 629 200 644 645 cell_1rw
* cell instance $20855 m0 *1 47.235,158.34
X$20855 199 630 200 644 645 cell_1rw
* cell instance $20856 m0 *1 47.235,161.07
X$20856 199 632 200 644 645 cell_1rw
* cell instance $20857 r0 *1 47.235,158.34
X$20857 199 631 200 644 645 cell_1rw
* cell instance $20858 r0 *1 47.235,161.07
X$20858 199 633 200 644 645 cell_1rw
* cell instance $20859 m0 *1 47.235,163.8
X$20859 199 634 200 644 645 cell_1rw
* cell instance $20860 m0 *1 47.235,166.53
X$20860 199 637 200 644 645 cell_1rw
* cell instance $20861 r0 *1 47.235,163.8
X$20861 199 635 200 644 645 cell_1rw
* cell instance $20862 m0 *1 47.235,169.26
X$20862 199 639 200 644 645 cell_1rw
* cell instance $20863 r0 *1 47.235,166.53
X$20863 199 636 200 644 645 cell_1rw
* cell instance $20864 r0 *1 47.235,169.26
X$20864 199 638 200 644 645 cell_1rw
* cell instance $20865 m0 *1 47.235,171.99
X$20865 199 640 200 644 645 cell_1rw
* cell instance $20866 m0 *1 47.235,174.72
X$20866 199 642 200 644 645 cell_1rw
* cell instance $20867 r0 *1 47.235,171.99
X$20867 199 641 200 644 645 cell_1rw
* cell instance $20868 r0 *1 47.235,174.72
X$20868 199 643 200 644 645 cell_1rw
* cell instance $20869 r0 *1 47.94,87.36
X$20869 201 322 202 644 645 cell_1rw
* cell instance $20870 m0 *1 47.94,90.09
X$20870 201 581 202 644 645 cell_1rw
* cell instance $20871 m0 *1 47.94,92.82
X$20871 201 583 202 644 645 cell_1rw
* cell instance $20872 r0 *1 47.94,90.09
X$20872 201 580 202 644 645 cell_1rw
* cell instance $20873 r0 *1 47.94,92.82
X$20873 201 582 202 644 645 cell_1rw
* cell instance $20874 m0 *1 47.94,95.55
X$20874 201 584 202 644 645 cell_1rw
* cell instance $20875 m0 *1 47.94,98.28
X$20875 201 586 202 644 645 cell_1rw
* cell instance $20876 r0 *1 47.94,95.55
X$20876 201 585 202 644 645 cell_1rw
* cell instance $20877 r0 *1 47.94,98.28
X$20877 201 587 202 644 645 cell_1rw
* cell instance $20878 m0 *1 47.94,101.01
X$20878 201 588 202 644 645 cell_1rw
* cell instance $20879 r0 *1 47.94,101.01
X$20879 201 589 202 644 645 cell_1rw
* cell instance $20880 m0 *1 47.94,103.74
X$20880 201 590 202 644 645 cell_1rw
* cell instance $20881 r0 *1 47.94,103.74
X$20881 201 591 202 644 645 cell_1rw
* cell instance $20882 m0 *1 47.94,106.47
X$20882 201 593 202 644 645 cell_1rw
* cell instance $20883 r0 *1 47.94,106.47
X$20883 201 592 202 644 645 cell_1rw
* cell instance $20884 m0 *1 47.94,109.2
X$20884 201 594 202 644 645 cell_1rw
* cell instance $20885 m0 *1 47.94,111.93
X$20885 201 597 202 644 645 cell_1rw
* cell instance $20886 r0 *1 47.94,109.2
X$20886 201 595 202 644 645 cell_1rw
* cell instance $20887 r0 *1 47.94,111.93
X$20887 201 596 202 644 645 cell_1rw
* cell instance $20888 m0 *1 47.94,114.66
X$20888 201 598 202 644 645 cell_1rw
* cell instance $20889 m0 *1 47.94,117.39
X$20889 201 600 202 644 645 cell_1rw
* cell instance $20890 r0 *1 47.94,114.66
X$20890 201 599 202 644 645 cell_1rw
* cell instance $20891 r0 *1 47.94,117.39
X$20891 201 601 202 644 645 cell_1rw
* cell instance $20892 m0 *1 47.94,120.12
X$20892 201 602 202 644 645 cell_1rw
* cell instance $20893 m0 *1 47.94,122.85
X$20893 201 604 202 644 645 cell_1rw
* cell instance $20894 r0 *1 47.94,120.12
X$20894 201 603 202 644 645 cell_1rw
* cell instance $20895 r0 *1 47.94,122.85
X$20895 201 605 202 644 645 cell_1rw
* cell instance $20896 m0 *1 47.94,125.58
X$20896 201 606 202 644 645 cell_1rw
* cell instance $20897 m0 *1 47.94,128.31
X$20897 201 609 202 644 645 cell_1rw
* cell instance $20898 r0 *1 47.94,125.58
X$20898 201 607 202 644 645 cell_1rw
* cell instance $20899 m0 *1 47.94,131.04
X$20899 201 610 202 644 645 cell_1rw
* cell instance $20900 r0 *1 47.94,128.31
X$20900 201 608 202 644 645 cell_1rw
* cell instance $20901 r0 *1 47.94,131.04
X$20901 201 611 202 644 645 cell_1rw
* cell instance $20902 m0 *1 47.94,133.77
X$20902 201 612 202 644 645 cell_1rw
* cell instance $20903 r0 *1 47.94,133.77
X$20903 201 613 202 644 645 cell_1rw
* cell instance $20904 m0 *1 47.94,136.5
X$20904 201 615 202 644 645 cell_1rw
* cell instance $20905 r0 *1 47.94,136.5
X$20905 201 614 202 644 645 cell_1rw
* cell instance $20906 m0 *1 47.94,139.23
X$20906 201 617 202 644 645 cell_1rw
* cell instance $20907 m0 *1 47.94,141.96
X$20907 201 618 202 644 645 cell_1rw
* cell instance $20908 r0 *1 47.94,139.23
X$20908 201 616 202 644 645 cell_1rw
* cell instance $20909 r0 *1 47.94,141.96
X$20909 201 619 202 644 645 cell_1rw
* cell instance $20910 m0 *1 47.94,144.69
X$20910 201 620 202 644 645 cell_1rw
* cell instance $20911 r0 *1 47.94,144.69
X$20911 201 621 202 644 645 cell_1rw
* cell instance $20912 m0 *1 47.94,147.42
X$20912 201 622 202 644 645 cell_1rw
* cell instance $20913 r0 *1 47.94,147.42
X$20913 201 623 202 644 645 cell_1rw
* cell instance $20914 m0 *1 47.94,150.15
X$20914 201 624 202 644 645 cell_1rw
* cell instance $20915 r0 *1 47.94,150.15
X$20915 201 625 202 644 645 cell_1rw
* cell instance $20916 m0 *1 47.94,152.88
X$20916 201 626 202 644 645 cell_1rw
* cell instance $20917 r0 *1 47.94,152.88
X$20917 201 627 202 644 645 cell_1rw
* cell instance $20918 m0 *1 47.94,155.61
X$20918 201 628 202 644 645 cell_1rw
* cell instance $20919 r0 *1 47.94,155.61
X$20919 201 629 202 644 645 cell_1rw
* cell instance $20920 m0 *1 47.94,158.34
X$20920 201 630 202 644 645 cell_1rw
* cell instance $20921 r0 *1 47.94,158.34
X$20921 201 631 202 644 645 cell_1rw
* cell instance $20922 m0 *1 47.94,161.07
X$20922 201 632 202 644 645 cell_1rw
* cell instance $20923 r0 *1 47.94,161.07
X$20923 201 633 202 644 645 cell_1rw
* cell instance $20924 m0 *1 47.94,163.8
X$20924 201 634 202 644 645 cell_1rw
* cell instance $20925 r0 *1 47.94,163.8
X$20925 201 635 202 644 645 cell_1rw
* cell instance $20926 m0 *1 47.94,166.53
X$20926 201 637 202 644 645 cell_1rw
* cell instance $20927 r0 *1 47.94,166.53
X$20927 201 636 202 644 645 cell_1rw
* cell instance $20928 m0 *1 47.94,169.26
X$20928 201 639 202 644 645 cell_1rw
* cell instance $20929 r0 *1 47.94,169.26
X$20929 201 638 202 644 645 cell_1rw
* cell instance $20930 m0 *1 47.94,171.99
X$20930 201 640 202 644 645 cell_1rw
* cell instance $20931 r0 *1 47.94,171.99
X$20931 201 641 202 644 645 cell_1rw
* cell instance $20932 m0 *1 47.94,174.72
X$20932 201 642 202 644 645 cell_1rw
* cell instance $20933 r0 *1 47.94,174.72
X$20933 201 643 202 644 645 cell_1rw
* cell instance $20934 r0 *1 48.645,87.36
X$20934 203 322 204 644 645 cell_1rw
* cell instance $20935 m0 *1 48.645,90.09
X$20935 203 581 204 644 645 cell_1rw
* cell instance $20936 m0 *1 48.645,92.82
X$20936 203 583 204 644 645 cell_1rw
* cell instance $20937 r0 *1 48.645,90.09
X$20937 203 580 204 644 645 cell_1rw
* cell instance $20938 m0 *1 48.645,95.55
X$20938 203 584 204 644 645 cell_1rw
* cell instance $20939 r0 *1 48.645,92.82
X$20939 203 582 204 644 645 cell_1rw
* cell instance $20940 m0 *1 48.645,98.28
X$20940 203 586 204 644 645 cell_1rw
* cell instance $20941 r0 *1 48.645,95.55
X$20941 203 585 204 644 645 cell_1rw
* cell instance $20942 r0 *1 48.645,98.28
X$20942 203 587 204 644 645 cell_1rw
* cell instance $20943 m0 *1 48.645,101.01
X$20943 203 588 204 644 645 cell_1rw
* cell instance $20944 m0 *1 48.645,103.74
X$20944 203 590 204 644 645 cell_1rw
* cell instance $20945 r0 *1 48.645,101.01
X$20945 203 589 204 644 645 cell_1rw
* cell instance $20946 r0 *1 48.645,103.74
X$20946 203 591 204 644 645 cell_1rw
* cell instance $20947 m0 *1 48.645,106.47
X$20947 203 593 204 644 645 cell_1rw
* cell instance $20948 r0 *1 48.645,106.47
X$20948 203 592 204 644 645 cell_1rw
* cell instance $20949 m0 *1 48.645,109.2
X$20949 203 594 204 644 645 cell_1rw
* cell instance $20950 r0 *1 48.645,109.2
X$20950 203 595 204 644 645 cell_1rw
* cell instance $20951 m0 *1 48.645,111.93
X$20951 203 597 204 644 645 cell_1rw
* cell instance $20952 r0 *1 48.645,111.93
X$20952 203 596 204 644 645 cell_1rw
* cell instance $20953 m0 *1 48.645,114.66
X$20953 203 598 204 644 645 cell_1rw
* cell instance $20954 r0 *1 48.645,114.66
X$20954 203 599 204 644 645 cell_1rw
* cell instance $20955 m0 *1 48.645,117.39
X$20955 203 600 204 644 645 cell_1rw
* cell instance $20956 r0 *1 48.645,117.39
X$20956 203 601 204 644 645 cell_1rw
* cell instance $20957 m0 *1 48.645,120.12
X$20957 203 602 204 644 645 cell_1rw
* cell instance $20958 m0 *1 48.645,122.85
X$20958 203 604 204 644 645 cell_1rw
* cell instance $20959 r0 *1 48.645,120.12
X$20959 203 603 204 644 645 cell_1rw
* cell instance $20960 r0 *1 48.645,122.85
X$20960 203 605 204 644 645 cell_1rw
* cell instance $20961 m0 *1 48.645,125.58
X$20961 203 606 204 644 645 cell_1rw
* cell instance $20962 r0 *1 48.645,125.58
X$20962 203 607 204 644 645 cell_1rw
* cell instance $20963 m0 *1 48.645,128.31
X$20963 203 609 204 644 645 cell_1rw
* cell instance $20964 r0 *1 48.645,128.31
X$20964 203 608 204 644 645 cell_1rw
* cell instance $20965 m0 *1 48.645,131.04
X$20965 203 610 204 644 645 cell_1rw
* cell instance $20966 r0 *1 48.645,131.04
X$20966 203 611 204 644 645 cell_1rw
* cell instance $20967 m0 *1 48.645,133.77
X$20967 203 612 204 644 645 cell_1rw
* cell instance $20968 r0 *1 48.645,133.77
X$20968 203 613 204 644 645 cell_1rw
* cell instance $20969 m0 *1 48.645,136.5
X$20969 203 615 204 644 645 cell_1rw
* cell instance $20970 r0 *1 48.645,136.5
X$20970 203 614 204 644 645 cell_1rw
* cell instance $20971 m0 *1 48.645,139.23
X$20971 203 617 204 644 645 cell_1rw
* cell instance $20972 r0 *1 48.645,139.23
X$20972 203 616 204 644 645 cell_1rw
* cell instance $20973 m0 *1 48.645,141.96
X$20973 203 618 204 644 645 cell_1rw
* cell instance $20974 m0 *1 48.645,144.69
X$20974 203 620 204 644 645 cell_1rw
* cell instance $20975 r0 *1 48.645,141.96
X$20975 203 619 204 644 645 cell_1rw
* cell instance $20976 m0 *1 48.645,147.42
X$20976 203 622 204 644 645 cell_1rw
* cell instance $20977 r0 *1 48.645,144.69
X$20977 203 621 204 644 645 cell_1rw
* cell instance $20978 r0 *1 48.645,147.42
X$20978 203 623 204 644 645 cell_1rw
* cell instance $20979 m0 *1 48.645,150.15
X$20979 203 624 204 644 645 cell_1rw
* cell instance $20980 r0 *1 48.645,150.15
X$20980 203 625 204 644 645 cell_1rw
* cell instance $20981 m0 *1 48.645,152.88
X$20981 203 626 204 644 645 cell_1rw
* cell instance $20982 r0 *1 48.645,152.88
X$20982 203 627 204 644 645 cell_1rw
* cell instance $20983 m0 *1 48.645,155.61
X$20983 203 628 204 644 645 cell_1rw
* cell instance $20984 r0 *1 48.645,155.61
X$20984 203 629 204 644 645 cell_1rw
* cell instance $20985 m0 *1 48.645,158.34
X$20985 203 630 204 644 645 cell_1rw
* cell instance $20986 r0 *1 48.645,158.34
X$20986 203 631 204 644 645 cell_1rw
* cell instance $20987 m0 *1 48.645,161.07
X$20987 203 632 204 644 645 cell_1rw
* cell instance $20988 r0 *1 48.645,161.07
X$20988 203 633 204 644 645 cell_1rw
* cell instance $20989 m0 *1 48.645,163.8
X$20989 203 634 204 644 645 cell_1rw
* cell instance $20990 r0 *1 48.645,163.8
X$20990 203 635 204 644 645 cell_1rw
* cell instance $20991 m0 *1 48.645,166.53
X$20991 203 637 204 644 645 cell_1rw
* cell instance $20992 r0 *1 48.645,166.53
X$20992 203 636 204 644 645 cell_1rw
* cell instance $20993 m0 *1 48.645,169.26
X$20993 203 639 204 644 645 cell_1rw
* cell instance $20994 r0 *1 48.645,169.26
X$20994 203 638 204 644 645 cell_1rw
* cell instance $20995 m0 *1 48.645,171.99
X$20995 203 640 204 644 645 cell_1rw
* cell instance $20996 r0 *1 48.645,171.99
X$20996 203 641 204 644 645 cell_1rw
* cell instance $20997 m0 *1 48.645,174.72
X$20997 203 642 204 644 645 cell_1rw
* cell instance $20998 r0 *1 48.645,174.72
X$20998 203 643 204 644 645 cell_1rw
* cell instance $20999 r0 *1 49.35,87.36
X$20999 205 322 206 644 645 cell_1rw
* cell instance $21000 m0 *1 49.35,90.09
X$21000 205 581 206 644 645 cell_1rw
* cell instance $21001 r0 *1 49.35,90.09
X$21001 205 580 206 644 645 cell_1rw
* cell instance $21002 m0 *1 49.35,92.82
X$21002 205 583 206 644 645 cell_1rw
* cell instance $21003 r0 *1 49.35,92.82
X$21003 205 582 206 644 645 cell_1rw
* cell instance $21004 m0 *1 49.35,95.55
X$21004 205 584 206 644 645 cell_1rw
* cell instance $21005 m0 *1 49.35,98.28
X$21005 205 586 206 644 645 cell_1rw
* cell instance $21006 r0 *1 49.35,95.55
X$21006 205 585 206 644 645 cell_1rw
* cell instance $21007 r0 *1 49.35,98.28
X$21007 205 587 206 644 645 cell_1rw
* cell instance $21008 m0 *1 49.35,101.01
X$21008 205 588 206 644 645 cell_1rw
* cell instance $21009 r0 *1 49.35,101.01
X$21009 205 589 206 644 645 cell_1rw
* cell instance $21010 m0 *1 49.35,103.74
X$21010 205 590 206 644 645 cell_1rw
* cell instance $21011 m0 *1 49.35,106.47
X$21011 205 593 206 644 645 cell_1rw
* cell instance $21012 r0 *1 49.35,103.74
X$21012 205 591 206 644 645 cell_1rw
* cell instance $21013 r0 *1 49.35,106.47
X$21013 205 592 206 644 645 cell_1rw
* cell instance $21014 m0 *1 49.35,109.2
X$21014 205 594 206 644 645 cell_1rw
* cell instance $21015 r0 *1 49.35,109.2
X$21015 205 595 206 644 645 cell_1rw
* cell instance $21016 m0 *1 49.35,111.93
X$21016 205 597 206 644 645 cell_1rw
* cell instance $21017 r0 *1 49.35,111.93
X$21017 205 596 206 644 645 cell_1rw
* cell instance $21018 m0 *1 49.35,114.66
X$21018 205 598 206 644 645 cell_1rw
* cell instance $21019 r0 *1 49.35,114.66
X$21019 205 599 206 644 645 cell_1rw
* cell instance $21020 m0 *1 49.35,117.39
X$21020 205 600 206 644 645 cell_1rw
* cell instance $21021 r0 *1 49.35,117.39
X$21021 205 601 206 644 645 cell_1rw
* cell instance $21022 m0 *1 49.35,120.12
X$21022 205 602 206 644 645 cell_1rw
* cell instance $21023 r0 *1 49.35,120.12
X$21023 205 603 206 644 645 cell_1rw
* cell instance $21024 m0 *1 49.35,122.85
X$21024 205 604 206 644 645 cell_1rw
* cell instance $21025 r0 *1 49.35,122.85
X$21025 205 605 206 644 645 cell_1rw
* cell instance $21026 m0 *1 49.35,125.58
X$21026 205 606 206 644 645 cell_1rw
* cell instance $21027 r0 *1 49.35,125.58
X$21027 205 607 206 644 645 cell_1rw
* cell instance $21028 m0 *1 49.35,128.31
X$21028 205 609 206 644 645 cell_1rw
* cell instance $21029 r0 *1 49.35,128.31
X$21029 205 608 206 644 645 cell_1rw
* cell instance $21030 m0 *1 49.35,131.04
X$21030 205 610 206 644 645 cell_1rw
* cell instance $21031 r0 *1 49.35,131.04
X$21031 205 611 206 644 645 cell_1rw
* cell instance $21032 m0 *1 49.35,133.77
X$21032 205 612 206 644 645 cell_1rw
* cell instance $21033 r0 *1 49.35,133.77
X$21033 205 613 206 644 645 cell_1rw
* cell instance $21034 m0 *1 49.35,136.5
X$21034 205 615 206 644 645 cell_1rw
* cell instance $21035 r0 *1 49.35,136.5
X$21035 205 614 206 644 645 cell_1rw
* cell instance $21036 m0 *1 49.35,139.23
X$21036 205 617 206 644 645 cell_1rw
* cell instance $21037 r0 *1 49.35,139.23
X$21037 205 616 206 644 645 cell_1rw
* cell instance $21038 m0 *1 49.35,141.96
X$21038 205 618 206 644 645 cell_1rw
* cell instance $21039 r0 *1 49.35,141.96
X$21039 205 619 206 644 645 cell_1rw
* cell instance $21040 m0 *1 49.35,144.69
X$21040 205 620 206 644 645 cell_1rw
* cell instance $21041 r0 *1 49.35,144.69
X$21041 205 621 206 644 645 cell_1rw
* cell instance $21042 m0 *1 49.35,147.42
X$21042 205 622 206 644 645 cell_1rw
* cell instance $21043 r0 *1 49.35,147.42
X$21043 205 623 206 644 645 cell_1rw
* cell instance $21044 m0 *1 49.35,150.15
X$21044 205 624 206 644 645 cell_1rw
* cell instance $21045 r0 *1 49.35,150.15
X$21045 205 625 206 644 645 cell_1rw
* cell instance $21046 m0 *1 49.35,152.88
X$21046 205 626 206 644 645 cell_1rw
* cell instance $21047 r0 *1 49.35,152.88
X$21047 205 627 206 644 645 cell_1rw
* cell instance $21048 m0 *1 49.35,155.61
X$21048 205 628 206 644 645 cell_1rw
* cell instance $21049 r0 *1 49.35,155.61
X$21049 205 629 206 644 645 cell_1rw
* cell instance $21050 m0 *1 49.35,158.34
X$21050 205 630 206 644 645 cell_1rw
* cell instance $21051 r0 *1 49.35,158.34
X$21051 205 631 206 644 645 cell_1rw
* cell instance $21052 m0 *1 49.35,161.07
X$21052 205 632 206 644 645 cell_1rw
* cell instance $21053 m0 *1 49.35,163.8
X$21053 205 634 206 644 645 cell_1rw
* cell instance $21054 r0 *1 49.35,161.07
X$21054 205 633 206 644 645 cell_1rw
* cell instance $21055 m0 *1 49.35,166.53
X$21055 205 637 206 644 645 cell_1rw
* cell instance $21056 r0 *1 49.35,163.8
X$21056 205 635 206 644 645 cell_1rw
* cell instance $21057 r0 *1 49.35,166.53
X$21057 205 636 206 644 645 cell_1rw
* cell instance $21058 m0 *1 49.35,169.26
X$21058 205 639 206 644 645 cell_1rw
* cell instance $21059 r0 *1 49.35,169.26
X$21059 205 638 206 644 645 cell_1rw
* cell instance $21060 m0 *1 49.35,171.99
X$21060 205 640 206 644 645 cell_1rw
* cell instance $21061 r0 *1 49.35,171.99
X$21061 205 641 206 644 645 cell_1rw
* cell instance $21062 m0 *1 49.35,174.72
X$21062 205 642 206 644 645 cell_1rw
* cell instance $21063 r0 *1 49.35,174.72
X$21063 205 643 206 644 645 cell_1rw
* cell instance $21064 r0 *1 50.055,87.36
X$21064 207 322 208 644 645 cell_1rw
* cell instance $21065 m0 *1 50.055,90.09
X$21065 207 581 208 644 645 cell_1rw
* cell instance $21066 r0 *1 50.055,90.09
X$21066 207 580 208 644 645 cell_1rw
* cell instance $21067 m0 *1 50.055,92.82
X$21067 207 583 208 644 645 cell_1rw
* cell instance $21068 r0 *1 50.055,92.82
X$21068 207 582 208 644 645 cell_1rw
* cell instance $21069 m0 *1 50.055,95.55
X$21069 207 584 208 644 645 cell_1rw
* cell instance $21070 r0 *1 50.055,95.55
X$21070 207 585 208 644 645 cell_1rw
* cell instance $21071 m0 *1 50.055,98.28
X$21071 207 586 208 644 645 cell_1rw
* cell instance $21072 r0 *1 50.055,98.28
X$21072 207 587 208 644 645 cell_1rw
* cell instance $21073 m0 *1 50.055,101.01
X$21073 207 588 208 644 645 cell_1rw
* cell instance $21074 r0 *1 50.055,101.01
X$21074 207 589 208 644 645 cell_1rw
* cell instance $21075 m0 *1 50.055,103.74
X$21075 207 590 208 644 645 cell_1rw
* cell instance $21076 r0 *1 50.055,103.74
X$21076 207 591 208 644 645 cell_1rw
* cell instance $21077 m0 *1 50.055,106.47
X$21077 207 593 208 644 645 cell_1rw
* cell instance $21078 r0 *1 50.055,106.47
X$21078 207 592 208 644 645 cell_1rw
* cell instance $21079 m0 *1 50.055,109.2
X$21079 207 594 208 644 645 cell_1rw
* cell instance $21080 r0 *1 50.055,109.2
X$21080 207 595 208 644 645 cell_1rw
* cell instance $21081 m0 *1 50.055,111.93
X$21081 207 597 208 644 645 cell_1rw
* cell instance $21082 r0 *1 50.055,111.93
X$21082 207 596 208 644 645 cell_1rw
* cell instance $21083 m0 *1 50.055,114.66
X$21083 207 598 208 644 645 cell_1rw
* cell instance $21084 r0 *1 50.055,114.66
X$21084 207 599 208 644 645 cell_1rw
* cell instance $21085 m0 *1 50.055,117.39
X$21085 207 600 208 644 645 cell_1rw
* cell instance $21086 r0 *1 50.055,117.39
X$21086 207 601 208 644 645 cell_1rw
* cell instance $21087 m0 *1 50.055,120.12
X$21087 207 602 208 644 645 cell_1rw
* cell instance $21088 r0 *1 50.055,120.12
X$21088 207 603 208 644 645 cell_1rw
* cell instance $21089 m0 *1 50.055,122.85
X$21089 207 604 208 644 645 cell_1rw
* cell instance $21090 r0 *1 50.055,122.85
X$21090 207 605 208 644 645 cell_1rw
* cell instance $21091 m0 *1 50.055,125.58
X$21091 207 606 208 644 645 cell_1rw
* cell instance $21092 r0 *1 50.055,125.58
X$21092 207 607 208 644 645 cell_1rw
* cell instance $21093 m0 *1 50.055,128.31
X$21093 207 609 208 644 645 cell_1rw
* cell instance $21094 m0 *1 50.055,131.04
X$21094 207 610 208 644 645 cell_1rw
* cell instance $21095 r0 *1 50.055,128.31
X$21095 207 608 208 644 645 cell_1rw
* cell instance $21096 r0 *1 50.055,131.04
X$21096 207 611 208 644 645 cell_1rw
* cell instance $21097 m0 *1 50.055,133.77
X$21097 207 612 208 644 645 cell_1rw
* cell instance $21098 r0 *1 50.055,133.77
X$21098 207 613 208 644 645 cell_1rw
* cell instance $21099 m0 *1 50.055,136.5
X$21099 207 615 208 644 645 cell_1rw
* cell instance $21100 r0 *1 50.055,136.5
X$21100 207 614 208 644 645 cell_1rw
* cell instance $21101 m0 *1 50.055,139.23
X$21101 207 617 208 644 645 cell_1rw
* cell instance $21102 m0 *1 50.055,141.96
X$21102 207 618 208 644 645 cell_1rw
* cell instance $21103 r0 *1 50.055,139.23
X$21103 207 616 208 644 645 cell_1rw
* cell instance $21104 r0 *1 50.055,141.96
X$21104 207 619 208 644 645 cell_1rw
* cell instance $21105 m0 *1 50.055,144.69
X$21105 207 620 208 644 645 cell_1rw
* cell instance $21106 r0 *1 50.055,144.69
X$21106 207 621 208 644 645 cell_1rw
* cell instance $21107 m0 *1 50.055,147.42
X$21107 207 622 208 644 645 cell_1rw
* cell instance $21108 m0 *1 50.055,150.15
X$21108 207 624 208 644 645 cell_1rw
* cell instance $21109 r0 *1 50.055,147.42
X$21109 207 623 208 644 645 cell_1rw
* cell instance $21110 r0 *1 50.055,150.15
X$21110 207 625 208 644 645 cell_1rw
* cell instance $21111 m0 *1 50.055,152.88
X$21111 207 626 208 644 645 cell_1rw
* cell instance $21112 r0 *1 50.055,152.88
X$21112 207 627 208 644 645 cell_1rw
* cell instance $21113 m0 *1 50.055,155.61
X$21113 207 628 208 644 645 cell_1rw
* cell instance $21114 r0 *1 50.055,155.61
X$21114 207 629 208 644 645 cell_1rw
* cell instance $21115 m0 *1 50.055,158.34
X$21115 207 630 208 644 645 cell_1rw
* cell instance $21116 r0 *1 50.055,158.34
X$21116 207 631 208 644 645 cell_1rw
* cell instance $21117 m0 *1 50.055,161.07
X$21117 207 632 208 644 645 cell_1rw
* cell instance $21118 r0 *1 50.055,161.07
X$21118 207 633 208 644 645 cell_1rw
* cell instance $21119 m0 *1 50.055,163.8
X$21119 207 634 208 644 645 cell_1rw
* cell instance $21120 r0 *1 50.055,163.8
X$21120 207 635 208 644 645 cell_1rw
* cell instance $21121 m0 *1 50.055,166.53
X$21121 207 637 208 644 645 cell_1rw
* cell instance $21122 m0 *1 50.055,169.26
X$21122 207 639 208 644 645 cell_1rw
* cell instance $21123 r0 *1 50.055,166.53
X$21123 207 636 208 644 645 cell_1rw
* cell instance $21124 r0 *1 50.055,169.26
X$21124 207 638 208 644 645 cell_1rw
* cell instance $21125 m0 *1 50.055,171.99
X$21125 207 640 208 644 645 cell_1rw
* cell instance $21126 r0 *1 50.055,171.99
X$21126 207 641 208 644 645 cell_1rw
* cell instance $21127 m0 *1 50.055,174.72
X$21127 207 642 208 644 645 cell_1rw
* cell instance $21128 r0 *1 50.055,174.72
X$21128 207 643 208 644 645 cell_1rw
* cell instance $21129 r0 *1 50.76,87.36
X$21129 209 322 210 644 645 cell_1rw
* cell instance $21130 m0 *1 50.76,90.09
X$21130 209 581 210 644 645 cell_1rw
* cell instance $21131 r0 *1 50.76,90.09
X$21131 209 580 210 644 645 cell_1rw
* cell instance $21132 m0 *1 50.76,92.82
X$21132 209 583 210 644 645 cell_1rw
* cell instance $21133 r0 *1 50.76,92.82
X$21133 209 582 210 644 645 cell_1rw
* cell instance $21134 m0 *1 50.76,95.55
X$21134 209 584 210 644 645 cell_1rw
* cell instance $21135 r0 *1 50.76,95.55
X$21135 209 585 210 644 645 cell_1rw
* cell instance $21136 m0 *1 50.76,98.28
X$21136 209 586 210 644 645 cell_1rw
* cell instance $21137 r0 *1 50.76,98.28
X$21137 209 587 210 644 645 cell_1rw
* cell instance $21138 m0 *1 50.76,101.01
X$21138 209 588 210 644 645 cell_1rw
* cell instance $21139 r0 *1 50.76,101.01
X$21139 209 589 210 644 645 cell_1rw
* cell instance $21140 m0 *1 50.76,103.74
X$21140 209 590 210 644 645 cell_1rw
* cell instance $21141 r0 *1 50.76,103.74
X$21141 209 591 210 644 645 cell_1rw
* cell instance $21142 m0 *1 50.76,106.47
X$21142 209 593 210 644 645 cell_1rw
* cell instance $21143 m0 *1 50.76,109.2
X$21143 209 594 210 644 645 cell_1rw
* cell instance $21144 r0 *1 50.76,106.47
X$21144 209 592 210 644 645 cell_1rw
* cell instance $21145 r0 *1 50.76,109.2
X$21145 209 595 210 644 645 cell_1rw
* cell instance $21146 m0 *1 50.76,111.93
X$21146 209 597 210 644 645 cell_1rw
* cell instance $21147 r0 *1 50.76,111.93
X$21147 209 596 210 644 645 cell_1rw
* cell instance $21148 m0 *1 50.76,114.66
X$21148 209 598 210 644 645 cell_1rw
* cell instance $21149 r0 *1 50.76,114.66
X$21149 209 599 210 644 645 cell_1rw
* cell instance $21150 m0 *1 50.76,117.39
X$21150 209 600 210 644 645 cell_1rw
* cell instance $21151 r0 *1 50.76,117.39
X$21151 209 601 210 644 645 cell_1rw
* cell instance $21152 m0 *1 50.76,120.12
X$21152 209 602 210 644 645 cell_1rw
* cell instance $21153 r0 *1 50.76,120.12
X$21153 209 603 210 644 645 cell_1rw
* cell instance $21154 m0 *1 50.76,122.85
X$21154 209 604 210 644 645 cell_1rw
* cell instance $21155 r0 *1 50.76,122.85
X$21155 209 605 210 644 645 cell_1rw
* cell instance $21156 m0 *1 50.76,125.58
X$21156 209 606 210 644 645 cell_1rw
* cell instance $21157 r0 *1 50.76,125.58
X$21157 209 607 210 644 645 cell_1rw
* cell instance $21158 m0 *1 50.76,128.31
X$21158 209 609 210 644 645 cell_1rw
* cell instance $21159 r0 *1 50.76,128.31
X$21159 209 608 210 644 645 cell_1rw
* cell instance $21160 m0 *1 50.76,131.04
X$21160 209 610 210 644 645 cell_1rw
* cell instance $21161 r0 *1 50.76,131.04
X$21161 209 611 210 644 645 cell_1rw
* cell instance $21162 m0 *1 50.76,133.77
X$21162 209 612 210 644 645 cell_1rw
* cell instance $21163 r0 *1 50.76,133.77
X$21163 209 613 210 644 645 cell_1rw
* cell instance $21164 m0 *1 50.76,136.5
X$21164 209 615 210 644 645 cell_1rw
* cell instance $21165 r0 *1 50.76,136.5
X$21165 209 614 210 644 645 cell_1rw
* cell instance $21166 m0 *1 50.76,139.23
X$21166 209 617 210 644 645 cell_1rw
* cell instance $21167 m0 *1 50.76,141.96
X$21167 209 618 210 644 645 cell_1rw
* cell instance $21168 r0 *1 50.76,139.23
X$21168 209 616 210 644 645 cell_1rw
* cell instance $21169 r0 *1 50.76,141.96
X$21169 209 619 210 644 645 cell_1rw
* cell instance $21170 m0 *1 50.76,144.69
X$21170 209 620 210 644 645 cell_1rw
* cell instance $21171 r0 *1 50.76,144.69
X$21171 209 621 210 644 645 cell_1rw
* cell instance $21172 m0 *1 50.76,147.42
X$21172 209 622 210 644 645 cell_1rw
* cell instance $21173 r0 *1 50.76,147.42
X$21173 209 623 210 644 645 cell_1rw
* cell instance $21174 m0 *1 50.76,150.15
X$21174 209 624 210 644 645 cell_1rw
* cell instance $21175 r0 *1 50.76,150.15
X$21175 209 625 210 644 645 cell_1rw
* cell instance $21176 m0 *1 50.76,152.88
X$21176 209 626 210 644 645 cell_1rw
* cell instance $21177 r0 *1 50.76,152.88
X$21177 209 627 210 644 645 cell_1rw
* cell instance $21178 m0 *1 50.76,155.61
X$21178 209 628 210 644 645 cell_1rw
* cell instance $21179 m0 *1 50.76,158.34
X$21179 209 630 210 644 645 cell_1rw
* cell instance $21180 r0 *1 50.76,155.61
X$21180 209 629 210 644 645 cell_1rw
* cell instance $21181 r0 *1 50.76,158.34
X$21181 209 631 210 644 645 cell_1rw
* cell instance $21182 m0 *1 50.76,161.07
X$21182 209 632 210 644 645 cell_1rw
* cell instance $21183 r0 *1 50.76,161.07
X$21183 209 633 210 644 645 cell_1rw
* cell instance $21184 m0 *1 50.76,163.8
X$21184 209 634 210 644 645 cell_1rw
* cell instance $21185 r0 *1 50.76,163.8
X$21185 209 635 210 644 645 cell_1rw
* cell instance $21186 m0 *1 50.76,166.53
X$21186 209 637 210 644 645 cell_1rw
* cell instance $21187 r0 *1 50.76,166.53
X$21187 209 636 210 644 645 cell_1rw
* cell instance $21188 m0 *1 50.76,169.26
X$21188 209 639 210 644 645 cell_1rw
* cell instance $21189 r0 *1 50.76,169.26
X$21189 209 638 210 644 645 cell_1rw
* cell instance $21190 m0 *1 50.76,171.99
X$21190 209 640 210 644 645 cell_1rw
* cell instance $21191 r0 *1 50.76,171.99
X$21191 209 641 210 644 645 cell_1rw
* cell instance $21192 m0 *1 50.76,174.72
X$21192 209 642 210 644 645 cell_1rw
* cell instance $21193 r0 *1 50.76,174.72
X$21193 209 643 210 644 645 cell_1rw
* cell instance $21194 r0 *1 51.465,87.36
X$21194 211 322 212 644 645 cell_1rw
* cell instance $21195 m0 *1 51.465,90.09
X$21195 211 581 212 644 645 cell_1rw
* cell instance $21196 r0 *1 51.465,90.09
X$21196 211 580 212 644 645 cell_1rw
* cell instance $21197 m0 *1 51.465,92.82
X$21197 211 583 212 644 645 cell_1rw
* cell instance $21198 r0 *1 51.465,92.82
X$21198 211 582 212 644 645 cell_1rw
* cell instance $21199 m0 *1 51.465,95.55
X$21199 211 584 212 644 645 cell_1rw
* cell instance $21200 r0 *1 51.465,95.55
X$21200 211 585 212 644 645 cell_1rw
* cell instance $21201 m0 *1 51.465,98.28
X$21201 211 586 212 644 645 cell_1rw
* cell instance $21202 m0 *1 51.465,101.01
X$21202 211 588 212 644 645 cell_1rw
* cell instance $21203 r0 *1 51.465,98.28
X$21203 211 587 212 644 645 cell_1rw
* cell instance $21204 r0 *1 51.465,101.01
X$21204 211 589 212 644 645 cell_1rw
* cell instance $21205 m0 *1 51.465,103.74
X$21205 211 590 212 644 645 cell_1rw
* cell instance $21206 r0 *1 51.465,103.74
X$21206 211 591 212 644 645 cell_1rw
* cell instance $21207 m0 *1 51.465,106.47
X$21207 211 593 212 644 645 cell_1rw
* cell instance $21208 r0 *1 51.465,106.47
X$21208 211 592 212 644 645 cell_1rw
* cell instance $21209 m0 *1 51.465,109.2
X$21209 211 594 212 644 645 cell_1rw
* cell instance $21210 r0 *1 51.465,109.2
X$21210 211 595 212 644 645 cell_1rw
* cell instance $21211 m0 *1 51.465,111.93
X$21211 211 597 212 644 645 cell_1rw
* cell instance $21212 m0 *1 51.465,114.66
X$21212 211 598 212 644 645 cell_1rw
* cell instance $21213 r0 *1 51.465,111.93
X$21213 211 596 212 644 645 cell_1rw
* cell instance $21214 r0 *1 51.465,114.66
X$21214 211 599 212 644 645 cell_1rw
* cell instance $21215 m0 *1 51.465,117.39
X$21215 211 600 212 644 645 cell_1rw
* cell instance $21216 r0 *1 51.465,117.39
X$21216 211 601 212 644 645 cell_1rw
* cell instance $21217 m0 *1 51.465,120.12
X$21217 211 602 212 644 645 cell_1rw
* cell instance $21218 r0 *1 51.465,120.12
X$21218 211 603 212 644 645 cell_1rw
* cell instance $21219 m0 *1 51.465,122.85
X$21219 211 604 212 644 645 cell_1rw
* cell instance $21220 r0 *1 51.465,122.85
X$21220 211 605 212 644 645 cell_1rw
* cell instance $21221 m0 *1 51.465,125.58
X$21221 211 606 212 644 645 cell_1rw
* cell instance $21222 r0 *1 51.465,125.58
X$21222 211 607 212 644 645 cell_1rw
* cell instance $21223 m0 *1 51.465,128.31
X$21223 211 609 212 644 645 cell_1rw
* cell instance $21224 r0 *1 51.465,128.31
X$21224 211 608 212 644 645 cell_1rw
* cell instance $21225 m0 *1 51.465,131.04
X$21225 211 610 212 644 645 cell_1rw
* cell instance $21226 m0 *1 51.465,133.77
X$21226 211 612 212 644 645 cell_1rw
* cell instance $21227 r0 *1 51.465,131.04
X$21227 211 611 212 644 645 cell_1rw
* cell instance $21228 r0 *1 51.465,133.77
X$21228 211 613 212 644 645 cell_1rw
* cell instance $21229 m0 *1 51.465,136.5
X$21229 211 615 212 644 645 cell_1rw
* cell instance $21230 m0 *1 51.465,139.23
X$21230 211 617 212 644 645 cell_1rw
* cell instance $21231 r0 *1 51.465,136.5
X$21231 211 614 212 644 645 cell_1rw
* cell instance $21232 r0 *1 51.465,139.23
X$21232 211 616 212 644 645 cell_1rw
* cell instance $21233 m0 *1 51.465,141.96
X$21233 211 618 212 644 645 cell_1rw
* cell instance $21234 m0 *1 51.465,144.69
X$21234 211 620 212 644 645 cell_1rw
* cell instance $21235 r0 *1 51.465,141.96
X$21235 211 619 212 644 645 cell_1rw
* cell instance $21236 r0 *1 51.465,144.69
X$21236 211 621 212 644 645 cell_1rw
* cell instance $21237 m0 *1 51.465,147.42
X$21237 211 622 212 644 645 cell_1rw
* cell instance $21238 r0 *1 51.465,147.42
X$21238 211 623 212 644 645 cell_1rw
* cell instance $21239 m0 *1 51.465,150.15
X$21239 211 624 212 644 645 cell_1rw
* cell instance $21240 r0 *1 51.465,150.15
X$21240 211 625 212 644 645 cell_1rw
* cell instance $21241 m0 *1 51.465,152.88
X$21241 211 626 212 644 645 cell_1rw
* cell instance $21242 r0 *1 51.465,152.88
X$21242 211 627 212 644 645 cell_1rw
* cell instance $21243 m0 *1 51.465,155.61
X$21243 211 628 212 644 645 cell_1rw
* cell instance $21244 r0 *1 51.465,155.61
X$21244 211 629 212 644 645 cell_1rw
* cell instance $21245 m0 *1 51.465,158.34
X$21245 211 630 212 644 645 cell_1rw
* cell instance $21246 r0 *1 51.465,158.34
X$21246 211 631 212 644 645 cell_1rw
* cell instance $21247 m0 *1 51.465,161.07
X$21247 211 632 212 644 645 cell_1rw
* cell instance $21248 r0 *1 51.465,161.07
X$21248 211 633 212 644 645 cell_1rw
* cell instance $21249 m0 *1 51.465,163.8
X$21249 211 634 212 644 645 cell_1rw
* cell instance $21250 m0 *1 51.465,166.53
X$21250 211 637 212 644 645 cell_1rw
* cell instance $21251 r0 *1 51.465,163.8
X$21251 211 635 212 644 645 cell_1rw
* cell instance $21252 r0 *1 51.465,166.53
X$21252 211 636 212 644 645 cell_1rw
* cell instance $21253 m0 *1 51.465,169.26
X$21253 211 639 212 644 645 cell_1rw
* cell instance $21254 r0 *1 51.465,169.26
X$21254 211 638 212 644 645 cell_1rw
* cell instance $21255 m0 *1 51.465,171.99
X$21255 211 640 212 644 645 cell_1rw
* cell instance $21256 r0 *1 51.465,171.99
X$21256 211 641 212 644 645 cell_1rw
* cell instance $21257 m0 *1 51.465,174.72
X$21257 211 642 212 644 645 cell_1rw
* cell instance $21258 r0 *1 51.465,174.72
X$21258 211 643 212 644 645 cell_1rw
* cell instance $21259 m0 *1 52.17,90.09
X$21259 213 581 214 644 645 cell_1rw
* cell instance $21260 r0 *1 52.17,87.36
X$21260 213 322 214 644 645 cell_1rw
* cell instance $21261 r0 *1 52.17,90.09
X$21261 213 580 214 644 645 cell_1rw
* cell instance $21262 m0 *1 52.17,92.82
X$21262 213 583 214 644 645 cell_1rw
* cell instance $21263 r0 *1 52.17,92.82
X$21263 213 582 214 644 645 cell_1rw
* cell instance $21264 m0 *1 52.17,95.55
X$21264 213 584 214 644 645 cell_1rw
* cell instance $21265 m0 *1 52.17,98.28
X$21265 213 586 214 644 645 cell_1rw
* cell instance $21266 r0 *1 52.17,95.55
X$21266 213 585 214 644 645 cell_1rw
* cell instance $21267 r0 *1 52.17,98.28
X$21267 213 587 214 644 645 cell_1rw
* cell instance $21268 m0 *1 52.17,101.01
X$21268 213 588 214 644 645 cell_1rw
* cell instance $21269 r0 *1 52.17,101.01
X$21269 213 589 214 644 645 cell_1rw
* cell instance $21270 m0 *1 52.17,103.74
X$21270 213 590 214 644 645 cell_1rw
* cell instance $21271 r0 *1 52.17,103.74
X$21271 213 591 214 644 645 cell_1rw
* cell instance $21272 m0 *1 52.17,106.47
X$21272 213 593 214 644 645 cell_1rw
* cell instance $21273 r0 *1 52.17,106.47
X$21273 213 592 214 644 645 cell_1rw
* cell instance $21274 m0 *1 52.17,109.2
X$21274 213 594 214 644 645 cell_1rw
* cell instance $21275 r0 *1 52.17,109.2
X$21275 213 595 214 644 645 cell_1rw
* cell instance $21276 m0 *1 52.17,111.93
X$21276 213 597 214 644 645 cell_1rw
* cell instance $21277 r0 *1 52.17,111.93
X$21277 213 596 214 644 645 cell_1rw
* cell instance $21278 m0 *1 52.17,114.66
X$21278 213 598 214 644 645 cell_1rw
* cell instance $21279 r0 *1 52.17,114.66
X$21279 213 599 214 644 645 cell_1rw
* cell instance $21280 m0 *1 52.17,117.39
X$21280 213 600 214 644 645 cell_1rw
* cell instance $21281 r0 *1 52.17,117.39
X$21281 213 601 214 644 645 cell_1rw
* cell instance $21282 m0 *1 52.17,120.12
X$21282 213 602 214 644 645 cell_1rw
* cell instance $21283 m0 *1 52.17,122.85
X$21283 213 604 214 644 645 cell_1rw
* cell instance $21284 r0 *1 52.17,120.12
X$21284 213 603 214 644 645 cell_1rw
* cell instance $21285 m0 *1 52.17,125.58
X$21285 213 606 214 644 645 cell_1rw
* cell instance $21286 r0 *1 52.17,122.85
X$21286 213 605 214 644 645 cell_1rw
* cell instance $21287 r0 *1 52.17,125.58
X$21287 213 607 214 644 645 cell_1rw
* cell instance $21288 m0 *1 52.17,128.31
X$21288 213 609 214 644 645 cell_1rw
* cell instance $21289 m0 *1 52.17,131.04
X$21289 213 610 214 644 645 cell_1rw
* cell instance $21290 r0 *1 52.17,128.31
X$21290 213 608 214 644 645 cell_1rw
* cell instance $21291 r0 *1 52.17,131.04
X$21291 213 611 214 644 645 cell_1rw
* cell instance $21292 m0 *1 52.17,133.77
X$21292 213 612 214 644 645 cell_1rw
* cell instance $21293 r0 *1 52.17,133.77
X$21293 213 613 214 644 645 cell_1rw
* cell instance $21294 m0 *1 52.17,136.5
X$21294 213 615 214 644 645 cell_1rw
* cell instance $21295 r0 *1 52.17,136.5
X$21295 213 614 214 644 645 cell_1rw
* cell instance $21296 m0 *1 52.17,139.23
X$21296 213 617 214 644 645 cell_1rw
* cell instance $21297 r0 *1 52.17,139.23
X$21297 213 616 214 644 645 cell_1rw
* cell instance $21298 m0 *1 52.17,141.96
X$21298 213 618 214 644 645 cell_1rw
* cell instance $21299 m0 *1 52.17,144.69
X$21299 213 620 214 644 645 cell_1rw
* cell instance $21300 r0 *1 52.17,141.96
X$21300 213 619 214 644 645 cell_1rw
* cell instance $21301 r0 *1 52.17,144.69
X$21301 213 621 214 644 645 cell_1rw
* cell instance $21302 m0 *1 52.17,147.42
X$21302 213 622 214 644 645 cell_1rw
* cell instance $21303 r0 *1 52.17,147.42
X$21303 213 623 214 644 645 cell_1rw
* cell instance $21304 m0 *1 52.17,150.15
X$21304 213 624 214 644 645 cell_1rw
* cell instance $21305 r0 *1 52.17,150.15
X$21305 213 625 214 644 645 cell_1rw
* cell instance $21306 m0 *1 52.17,152.88
X$21306 213 626 214 644 645 cell_1rw
* cell instance $21307 m0 *1 52.17,155.61
X$21307 213 628 214 644 645 cell_1rw
* cell instance $21308 r0 *1 52.17,152.88
X$21308 213 627 214 644 645 cell_1rw
* cell instance $21309 r0 *1 52.17,155.61
X$21309 213 629 214 644 645 cell_1rw
* cell instance $21310 m0 *1 52.17,158.34
X$21310 213 630 214 644 645 cell_1rw
* cell instance $21311 r0 *1 52.17,158.34
X$21311 213 631 214 644 645 cell_1rw
* cell instance $21312 m0 *1 52.17,161.07
X$21312 213 632 214 644 645 cell_1rw
* cell instance $21313 m0 *1 52.17,163.8
X$21313 213 634 214 644 645 cell_1rw
* cell instance $21314 r0 *1 52.17,161.07
X$21314 213 633 214 644 645 cell_1rw
* cell instance $21315 m0 *1 52.17,166.53
X$21315 213 637 214 644 645 cell_1rw
* cell instance $21316 r0 *1 52.17,163.8
X$21316 213 635 214 644 645 cell_1rw
* cell instance $21317 r0 *1 52.17,166.53
X$21317 213 636 214 644 645 cell_1rw
* cell instance $21318 m0 *1 52.17,169.26
X$21318 213 639 214 644 645 cell_1rw
* cell instance $21319 r0 *1 52.17,169.26
X$21319 213 638 214 644 645 cell_1rw
* cell instance $21320 m0 *1 52.17,171.99
X$21320 213 640 214 644 645 cell_1rw
* cell instance $21321 r0 *1 52.17,171.99
X$21321 213 641 214 644 645 cell_1rw
* cell instance $21322 m0 *1 52.17,174.72
X$21322 213 642 214 644 645 cell_1rw
* cell instance $21323 r0 *1 52.17,174.72
X$21323 213 643 214 644 645 cell_1rw
* cell instance $21324 m0 *1 52.875,90.09
X$21324 215 581 216 644 645 cell_1rw
* cell instance $21325 r0 *1 52.875,87.36
X$21325 215 322 216 644 645 cell_1rw
* cell instance $21326 r0 *1 52.875,90.09
X$21326 215 580 216 644 645 cell_1rw
* cell instance $21327 m0 *1 52.875,92.82
X$21327 215 583 216 644 645 cell_1rw
* cell instance $21328 r0 *1 52.875,92.82
X$21328 215 582 216 644 645 cell_1rw
* cell instance $21329 m0 *1 52.875,95.55
X$21329 215 584 216 644 645 cell_1rw
* cell instance $21330 r0 *1 52.875,95.55
X$21330 215 585 216 644 645 cell_1rw
* cell instance $21331 m0 *1 52.875,98.28
X$21331 215 586 216 644 645 cell_1rw
* cell instance $21332 r0 *1 52.875,98.28
X$21332 215 587 216 644 645 cell_1rw
* cell instance $21333 m0 *1 52.875,101.01
X$21333 215 588 216 644 645 cell_1rw
* cell instance $21334 m0 *1 52.875,103.74
X$21334 215 590 216 644 645 cell_1rw
* cell instance $21335 r0 *1 52.875,101.01
X$21335 215 589 216 644 645 cell_1rw
* cell instance $21336 r0 *1 52.875,103.74
X$21336 215 591 216 644 645 cell_1rw
* cell instance $21337 m0 *1 52.875,106.47
X$21337 215 593 216 644 645 cell_1rw
* cell instance $21338 r0 *1 52.875,106.47
X$21338 215 592 216 644 645 cell_1rw
* cell instance $21339 m0 *1 52.875,109.2
X$21339 215 594 216 644 645 cell_1rw
* cell instance $21340 m0 *1 52.875,111.93
X$21340 215 597 216 644 645 cell_1rw
* cell instance $21341 r0 *1 52.875,109.2
X$21341 215 595 216 644 645 cell_1rw
* cell instance $21342 r0 *1 52.875,111.93
X$21342 215 596 216 644 645 cell_1rw
* cell instance $21343 m0 *1 52.875,114.66
X$21343 215 598 216 644 645 cell_1rw
* cell instance $21344 r0 *1 52.875,114.66
X$21344 215 599 216 644 645 cell_1rw
* cell instance $21345 m0 *1 52.875,117.39
X$21345 215 600 216 644 645 cell_1rw
* cell instance $21346 r0 *1 52.875,117.39
X$21346 215 601 216 644 645 cell_1rw
* cell instance $21347 m0 *1 52.875,120.12
X$21347 215 602 216 644 645 cell_1rw
* cell instance $21348 r0 *1 52.875,120.12
X$21348 215 603 216 644 645 cell_1rw
* cell instance $21349 m0 *1 52.875,122.85
X$21349 215 604 216 644 645 cell_1rw
* cell instance $21350 r0 *1 52.875,122.85
X$21350 215 605 216 644 645 cell_1rw
* cell instance $21351 m0 *1 52.875,125.58
X$21351 215 606 216 644 645 cell_1rw
* cell instance $21352 r0 *1 52.875,125.58
X$21352 215 607 216 644 645 cell_1rw
* cell instance $21353 m0 *1 52.875,128.31
X$21353 215 609 216 644 645 cell_1rw
* cell instance $21354 r0 *1 52.875,128.31
X$21354 215 608 216 644 645 cell_1rw
* cell instance $21355 m0 *1 52.875,131.04
X$21355 215 610 216 644 645 cell_1rw
* cell instance $21356 r0 *1 52.875,131.04
X$21356 215 611 216 644 645 cell_1rw
* cell instance $21357 m0 *1 52.875,133.77
X$21357 215 612 216 644 645 cell_1rw
* cell instance $21358 r0 *1 52.875,133.77
X$21358 215 613 216 644 645 cell_1rw
* cell instance $21359 m0 *1 52.875,136.5
X$21359 215 615 216 644 645 cell_1rw
* cell instance $21360 r0 *1 52.875,136.5
X$21360 215 614 216 644 645 cell_1rw
* cell instance $21361 m0 *1 52.875,139.23
X$21361 215 617 216 644 645 cell_1rw
* cell instance $21362 r0 *1 52.875,139.23
X$21362 215 616 216 644 645 cell_1rw
* cell instance $21363 m0 *1 52.875,141.96
X$21363 215 618 216 644 645 cell_1rw
* cell instance $21364 r0 *1 52.875,141.96
X$21364 215 619 216 644 645 cell_1rw
* cell instance $21365 m0 *1 52.875,144.69
X$21365 215 620 216 644 645 cell_1rw
* cell instance $21366 r0 *1 52.875,144.69
X$21366 215 621 216 644 645 cell_1rw
* cell instance $21367 m0 *1 52.875,147.42
X$21367 215 622 216 644 645 cell_1rw
* cell instance $21368 r0 *1 52.875,147.42
X$21368 215 623 216 644 645 cell_1rw
* cell instance $21369 m0 *1 52.875,150.15
X$21369 215 624 216 644 645 cell_1rw
* cell instance $21370 r0 *1 52.875,150.15
X$21370 215 625 216 644 645 cell_1rw
* cell instance $21371 m0 *1 52.875,152.88
X$21371 215 626 216 644 645 cell_1rw
* cell instance $21372 r0 *1 52.875,152.88
X$21372 215 627 216 644 645 cell_1rw
* cell instance $21373 m0 *1 52.875,155.61
X$21373 215 628 216 644 645 cell_1rw
* cell instance $21374 m0 *1 52.875,158.34
X$21374 215 630 216 644 645 cell_1rw
* cell instance $21375 r0 *1 52.875,155.61
X$21375 215 629 216 644 645 cell_1rw
* cell instance $21376 r0 *1 52.875,158.34
X$21376 215 631 216 644 645 cell_1rw
* cell instance $21377 m0 *1 52.875,161.07
X$21377 215 632 216 644 645 cell_1rw
* cell instance $21378 r0 *1 52.875,161.07
X$21378 215 633 216 644 645 cell_1rw
* cell instance $21379 m0 *1 52.875,163.8
X$21379 215 634 216 644 645 cell_1rw
* cell instance $21380 r0 *1 52.875,163.8
X$21380 215 635 216 644 645 cell_1rw
* cell instance $21381 m0 *1 52.875,166.53
X$21381 215 637 216 644 645 cell_1rw
* cell instance $21382 r0 *1 52.875,166.53
X$21382 215 636 216 644 645 cell_1rw
* cell instance $21383 m0 *1 52.875,169.26
X$21383 215 639 216 644 645 cell_1rw
* cell instance $21384 r0 *1 52.875,169.26
X$21384 215 638 216 644 645 cell_1rw
* cell instance $21385 m0 *1 52.875,171.99
X$21385 215 640 216 644 645 cell_1rw
* cell instance $21386 m0 *1 52.875,174.72
X$21386 215 642 216 644 645 cell_1rw
* cell instance $21387 r0 *1 52.875,171.99
X$21387 215 641 216 644 645 cell_1rw
* cell instance $21388 r0 *1 52.875,174.72
X$21388 215 643 216 644 645 cell_1rw
* cell instance $21389 m0 *1 53.58,90.09
X$21389 217 581 218 644 645 cell_1rw
* cell instance $21390 r0 *1 53.58,87.36
X$21390 217 322 218 644 645 cell_1rw
* cell instance $21391 r0 *1 53.58,90.09
X$21391 217 580 218 644 645 cell_1rw
* cell instance $21392 m0 *1 53.58,92.82
X$21392 217 583 218 644 645 cell_1rw
* cell instance $21393 r0 *1 53.58,92.82
X$21393 217 582 218 644 645 cell_1rw
* cell instance $21394 m0 *1 53.58,95.55
X$21394 217 584 218 644 645 cell_1rw
* cell instance $21395 r0 *1 53.58,95.55
X$21395 217 585 218 644 645 cell_1rw
* cell instance $21396 m0 *1 53.58,98.28
X$21396 217 586 218 644 645 cell_1rw
* cell instance $21397 m0 *1 53.58,101.01
X$21397 217 588 218 644 645 cell_1rw
* cell instance $21398 r0 *1 53.58,98.28
X$21398 217 587 218 644 645 cell_1rw
* cell instance $21399 r0 *1 53.58,101.01
X$21399 217 589 218 644 645 cell_1rw
* cell instance $21400 m0 *1 53.58,103.74
X$21400 217 590 218 644 645 cell_1rw
* cell instance $21401 r0 *1 53.58,103.74
X$21401 217 591 218 644 645 cell_1rw
* cell instance $21402 m0 *1 53.58,106.47
X$21402 217 593 218 644 645 cell_1rw
* cell instance $21403 r0 *1 53.58,106.47
X$21403 217 592 218 644 645 cell_1rw
* cell instance $21404 m0 *1 53.58,109.2
X$21404 217 594 218 644 645 cell_1rw
* cell instance $21405 r0 *1 53.58,109.2
X$21405 217 595 218 644 645 cell_1rw
* cell instance $21406 m0 *1 53.58,111.93
X$21406 217 597 218 644 645 cell_1rw
* cell instance $21407 r0 *1 53.58,111.93
X$21407 217 596 218 644 645 cell_1rw
* cell instance $21408 m0 *1 53.58,114.66
X$21408 217 598 218 644 645 cell_1rw
* cell instance $21409 m0 *1 53.58,117.39
X$21409 217 600 218 644 645 cell_1rw
* cell instance $21410 r0 *1 53.58,114.66
X$21410 217 599 218 644 645 cell_1rw
* cell instance $21411 r0 *1 53.58,117.39
X$21411 217 601 218 644 645 cell_1rw
* cell instance $21412 m0 *1 53.58,120.12
X$21412 217 602 218 644 645 cell_1rw
* cell instance $21413 r0 *1 53.58,120.12
X$21413 217 603 218 644 645 cell_1rw
* cell instance $21414 m0 *1 53.58,122.85
X$21414 217 604 218 644 645 cell_1rw
* cell instance $21415 m0 *1 53.58,125.58
X$21415 217 606 218 644 645 cell_1rw
* cell instance $21416 r0 *1 53.58,122.85
X$21416 217 605 218 644 645 cell_1rw
* cell instance $21417 r0 *1 53.58,125.58
X$21417 217 607 218 644 645 cell_1rw
* cell instance $21418 m0 *1 53.58,128.31
X$21418 217 609 218 644 645 cell_1rw
* cell instance $21419 r0 *1 53.58,128.31
X$21419 217 608 218 644 645 cell_1rw
* cell instance $21420 m0 *1 53.58,131.04
X$21420 217 610 218 644 645 cell_1rw
* cell instance $21421 r0 *1 53.58,131.04
X$21421 217 611 218 644 645 cell_1rw
* cell instance $21422 m0 *1 53.58,133.77
X$21422 217 612 218 644 645 cell_1rw
* cell instance $21423 r0 *1 53.58,133.77
X$21423 217 613 218 644 645 cell_1rw
* cell instance $21424 m0 *1 53.58,136.5
X$21424 217 615 218 644 645 cell_1rw
* cell instance $21425 r0 *1 53.58,136.5
X$21425 217 614 218 644 645 cell_1rw
* cell instance $21426 m0 *1 53.58,139.23
X$21426 217 617 218 644 645 cell_1rw
* cell instance $21427 r0 *1 53.58,139.23
X$21427 217 616 218 644 645 cell_1rw
* cell instance $21428 m0 *1 53.58,141.96
X$21428 217 618 218 644 645 cell_1rw
* cell instance $21429 r0 *1 53.58,141.96
X$21429 217 619 218 644 645 cell_1rw
* cell instance $21430 m0 *1 53.58,144.69
X$21430 217 620 218 644 645 cell_1rw
* cell instance $21431 r0 *1 53.58,144.69
X$21431 217 621 218 644 645 cell_1rw
* cell instance $21432 m0 *1 53.58,147.42
X$21432 217 622 218 644 645 cell_1rw
* cell instance $21433 r0 *1 53.58,147.42
X$21433 217 623 218 644 645 cell_1rw
* cell instance $21434 m0 *1 53.58,150.15
X$21434 217 624 218 644 645 cell_1rw
* cell instance $21435 r0 *1 53.58,150.15
X$21435 217 625 218 644 645 cell_1rw
* cell instance $21436 m0 *1 53.58,152.88
X$21436 217 626 218 644 645 cell_1rw
* cell instance $21437 r0 *1 53.58,152.88
X$21437 217 627 218 644 645 cell_1rw
* cell instance $21438 m0 *1 53.58,155.61
X$21438 217 628 218 644 645 cell_1rw
* cell instance $21439 r0 *1 53.58,155.61
X$21439 217 629 218 644 645 cell_1rw
* cell instance $21440 m0 *1 53.58,158.34
X$21440 217 630 218 644 645 cell_1rw
* cell instance $21441 r0 *1 53.58,158.34
X$21441 217 631 218 644 645 cell_1rw
* cell instance $21442 m0 *1 53.58,161.07
X$21442 217 632 218 644 645 cell_1rw
* cell instance $21443 r0 *1 53.58,161.07
X$21443 217 633 218 644 645 cell_1rw
* cell instance $21444 m0 *1 53.58,163.8
X$21444 217 634 218 644 645 cell_1rw
* cell instance $21445 m0 *1 53.58,166.53
X$21445 217 637 218 644 645 cell_1rw
* cell instance $21446 r0 *1 53.58,163.8
X$21446 217 635 218 644 645 cell_1rw
* cell instance $21447 r0 *1 53.58,166.53
X$21447 217 636 218 644 645 cell_1rw
* cell instance $21448 m0 *1 53.58,169.26
X$21448 217 639 218 644 645 cell_1rw
* cell instance $21449 r0 *1 53.58,169.26
X$21449 217 638 218 644 645 cell_1rw
* cell instance $21450 m0 *1 53.58,171.99
X$21450 217 640 218 644 645 cell_1rw
* cell instance $21451 r0 *1 53.58,171.99
X$21451 217 641 218 644 645 cell_1rw
* cell instance $21452 m0 *1 53.58,174.72
X$21452 217 642 218 644 645 cell_1rw
* cell instance $21453 r0 *1 53.58,174.72
X$21453 217 643 218 644 645 cell_1rw
* cell instance $21454 m0 *1 54.285,90.09
X$21454 219 581 220 644 645 cell_1rw
* cell instance $21455 r0 *1 54.285,87.36
X$21455 219 322 220 644 645 cell_1rw
* cell instance $21456 r0 *1 54.285,90.09
X$21456 219 580 220 644 645 cell_1rw
* cell instance $21457 m0 *1 54.285,92.82
X$21457 219 583 220 644 645 cell_1rw
* cell instance $21458 r0 *1 54.285,92.82
X$21458 219 582 220 644 645 cell_1rw
* cell instance $21459 m0 *1 54.285,95.55
X$21459 219 584 220 644 645 cell_1rw
* cell instance $21460 r0 *1 54.285,95.55
X$21460 219 585 220 644 645 cell_1rw
* cell instance $21461 m0 *1 54.285,98.28
X$21461 219 586 220 644 645 cell_1rw
* cell instance $21462 r0 *1 54.285,98.28
X$21462 219 587 220 644 645 cell_1rw
* cell instance $21463 m0 *1 54.285,101.01
X$21463 219 588 220 644 645 cell_1rw
* cell instance $21464 r0 *1 54.285,101.01
X$21464 219 589 220 644 645 cell_1rw
* cell instance $21465 m0 *1 54.285,103.74
X$21465 219 590 220 644 645 cell_1rw
* cell instance $21466 r0 *1 54.285,103.74
X$21466 219 591 220 644 645 cell_1rw
* cell instance $21467 m0 *1 54.285,106.47
X$21467 219 593 220 644 645 cell_1rw
* cell instance $21468 r0 *1 54.285,106.47
X$21468 219 592 220 644 645 cell_1rw
* cell instance $21469 m0 *1 54.285,109.2
X$21469 219 594 220 644 645 cell_1rw
* cell instance $21470 r0 *1 54.285,109.2
X$21470 219 595 220 644 645 cell_1rw
* cell instance $21471 m0 *1 54.285,111.93
X$21471 219 597 220 644 645 cell_1rw
* cell instance $21472 m0 *1 54.285,114.66
X$21472 219 598 220 644 645 cell_1rw
* cell instance $21473 r0 *1 54.285,111.93
X$21473 219 596 220 644 645 cell_1rw
* cell instance $21474 r0 *1 54.285,114.66
X$21474 219 599 220 644 645 cell_1rw
* cell instance $21475 m0 *1 54.285,117.39
X$21475 219 600 220 644 645 cell_1rw
* cell instance $21476 r0 *1 54.285,117.39
X$21476 219 601 220 644 645 cell_1rw
* cell instance $21477 m0 *1 54.285,120.12
X$21477 219 602 220 644 645 cell_1rw
* cell instance $21478 r0 *1 54.285,120.12
X$21478 219 603 220 644 645 cell_1rw
* cell instance $21479 m0 *1 54.285,122.85
X$21479 219 604 220 644 645 cell_1rw
* cell instance $21480 r0 *1 54.285,122.85
X$21480 219 605 220 644 645 cell_1rw
* cell instance $21481 m0 *1 54.285,125.58
X$21481 219 606 220 644 645 cell_1rw
* cell instance $21482 r0 *1 54.285,125.58
X$21482 219 607 220 644 645 cell_1rw
* cell instance $21483 m0 *1 54.285,128.31
X$21483 219 609 220 644 645 cell_1rw
* cell instance $21484 r0 *1 54.285,128.31
X$21484 219 608 220 644 645 cell_1rw
* cell instance $21485 m0 *1 54.285,131.04
X$21485 219 610 220 644 645 cell_1rw
* cell instance $21486 r0 *1 54.285,131.04
X$21486 219 611 220 644 645 cell_1rw
* cell instance $21487 m0 *1 54.285,133.77
X$21487 219 612 220 644 645 cell_1rw
* cell instance $21488 r0 *1 54.285,133.77
X$21488 219 613 220 644 645 cell_1rw
* cell instance $21489 m0 *1 54.285,136.5
X$21489 219 615 220 644 645 cell_1rw
* cell instance $21490 r0 *1 54.285,136.5
X$21490 219 614 220 644 645 cell_1rw
* cell instance $21491 m0 *1 54.285,139.23
X$21491 219 617 220 644 645 cell_1rw
* cell instance $21492 r0 *1 54.285,139.23
X$21492 219 616 220 644 645 cell_1rw
* cell instance $21493 m0 *1 54.285,141.96
X$21493 219 618 220 644 645 cell_1rw
* cell instance $21494 r0 *1 54.285,141.96
X$21494 219 619 220 644 645 cell_1rw
* cell instance $21495 m0 *1 54.285,144.69
X$21495 219 620 220 644 645 cell_1rw
* cell instance $21496 r0 *1 54.285,144.69
X$21496 219 621 220 644 645 cell_1rw
* cell instance $21497 m0 *1 54.285,147.42
X$21497 219 622 220 644 645 cell_1rw
* cell instance $21498 r0 *1 54.285,147.42
X$21498 219 623 220 644 645 cell_1rw
* cell instance $21499 m0 *1 54.285,150.15
X$21499 219 624 220 644 645 cell_1rw
* cell instance $21500 r0 *1 54.285,150.15
X$21500 219 625 220 644 645 cell_1rw
* cell instance $21501 m0 *1 54.285,152.88
X$21501 219 626 220 644 645 cell_1rw
* cell instance $21502 r0 *1 54.285,152.88
X$21502 219 627 220 644 645 cell_1rw
* cell instance $21503 m0 *1 54.285,155.61
X$21503 219 628 220 644 645 cell_1rw
* cell instance $21504 m0 *1 54.285,158.34
X$21504 219 630 220 644 645 cell_1rw
* cell instance $21505 r0 *1 54.285,155.61
X$21505 219 629 220 644 645 cell_1rw
* cell instance $21506 m0 *1 54.285,161.07
X$21506 219 632 220 644 645 cell_1rw
* cell instance $21507 r0 *1 54.285,158.34
X$21507 219 631 220 644 645 cell_1rw
* cell instance $21508 m0 *1 54.285,163.8
X$21508 219 634 220 644 645 cell_1rw
* cell instance $21509 r0 *1 54.285,161.07
X$21509 219 633 220 644 645 cell_1rw
* cell instance $21510 r0 *1 54.285,163.8
X$21510 219 635 220 644 645 cell_1rw
* cell instance $21511 m0 *1 54.285,166.53
X$21511 219 637 220 644 645 cell_1rw
* cell instance $21512 r0 *1 54.285,166.53
X$21512 219 636 220 644 645 cell_1rw
* cell instance $21513 m0 *1 54.285,169.26
X$21513 219 639 220 644 645 cell_1rw
* cell instance $21514 r0 *1 54.285,169.26
X$21514 219 638 220 644 645 cell_1rw
* cell instance $21515 m0 *1 54.285,171.99
X$21515 219 640 220 644 645 cell_1rw
* cell instance $21516 m0 *1 54.285,174.72
X$21516 219 642 220 644 645 cell_1rw
* cell instance $21517 r0 *1 54.285,171.99
X$21517 219 641 220 644 645 cell_1rw
* cell instance $21518 r0 *1 54.285,174.72
X$21518 219 643 220 644 645 cell_1rw
* cell instance $21519 r0 *1 54.99,87.36
X$21519 221 322 222 644 645 cell_1rw
* cell instance $21520 m0 *1 54.99,90.09
X$21520 221 581 222 644 645 cell_1rw
* cell instance $21521 r0 *1 54.99,90.09
X$21521 221 580 222 644 645 cell_1rw
* cell instance $21522 m0 *1 54.99,92.82
X$21522 221 583 222 644 645 cell_1rw
* cell instance $21523 r0 *1 54.99,92.82
X$21523 221 582 222 644 645 cell_1rw
* cell instance $21524 m0 *1 54.99,95.55
X$21524 221 584 222 644 645 cell_1rw
* cell instance $21525 r0 *1 54.99,95.55
X$21525 221 585 222 644 645 cell_1rw
* cell instance $21526 m0 *1 54.99,98.28
X$21526 221 586 222 644 645 cell_1rw
* cell instance $21527 r0 *1 54.99,98.28
X$21527 221 587 222 644 645 cell_1rw
* cell instance $21528 m0 *1 54.99,101.01
X$21528 221 588 222 644 645 cell_1rw
* cell instance $21529 m0 *1 54.99,103.74
X$21529 221 590 222 644 645 cell_1rw
* cell instance $21530 r0 *1 54.99,101.01
X$21530 221 589 222 644 645 cell_1rw
* cell instance $21531 r0 *1 54.99,103.74
X$21531 221 591 222 644 645 cell_1rw
* cell instance $21532 m0 *1 54.99,106.47
X$21532 221 593 222 644 645 cell_1rw
* cell instance $21533 r0 *1 54.99,106.47
X$21533 221 592 222 644 645 cell_1rw
* cell instance $21534 m0 *1 54.99,109.2
X$21534 221 594 222 644 645 cell_1rw
* cell instance $21535 m0 *1 54.99,111.93
X$21535 221 597 222 644 645 cell_1rw
* cell instance $21536 r0 *1 54.99,109.2
X$21536 221 595 222 644 645 cell_1rw
* cell instance $21537 m0 *1 54.99,114.66
X$21537 221 598 222 644 645 cell_1rw
* cell instance $21538 r0 *1 54.99,111.93
X$21538 221 596 222 644 645 cell_1rw
* cell instance $21539 r0 *1 54.99,114.66
X$21539 221 599 222 644 645 cell_1rw
* cell instance $21540 m0 *1 54.99,117.39
X$21540 221 600 222 644 645 cell_1rw
* cell instance $21541 r0 *1 54.99,117.39
X$21541 221 601 222 644 645 cell_1rw
* cell instance $21542 m0 *1 54.99,120.12
X$21542 221 602 222 644 645 cell_1rw
* cell instance $21543 r0 *1 54.99,120.12
X$21543 221 603 222 644 645 cell_1rw
* cell instance $21544 m0 *1 54.99,122.85
X$21544 221 604 222 644 645 cell_1rw
* cell instance $21545 r0 *1 54.99,122.85
X$21545 221 605 222 644 645 cell_1rw
* cell instance $21546 m0 *1 54.99,125.58
X$21546 221 606 222 644 645 cell_1rw
* cell instance $21547 m0 *1 54.99,128.31
X$21547 221 609 222 644 645 cell_1rw
* cell instance $21548 r0 *1 54.99,125.58
X$21548 221 607 222 644 645 cell_1rw
* cell instance $21549 r0 *1 54.99,128.31
X$21549 221 608 222 644 645 cell_1rw
* cell instance $21550 m0 *1 54.99,131.04
X$21550 221 610 222 644 645 cell_1rw
* cell instance $21551 r0 *1 54.99,131.04
X$21551 221 611 222 644 645 cell_1rw
* cell instance $21552 m0 *1 54.99,133.77
X$21552 221 612 222 644 645 cell_1rw
* cell instance $21553 r0 *1 54.99,133.77
X$21553 221 613 222 644 645 cell_1rw
* cell instance $21554 m0 *1 54.99,136.5
X$21554 221 615 222 644 645 cell_1rw
* cell instance $21555 r0 *1 54.99,136.5
X$21555 221 614 222 644 645 cell_1rw
* cell instance $21556 m0 *1 54.99,139.23
X$21556 221 617 222 644 645 cell_1rw
* cell instance $21557 r0 *1 54.99,139.23
X$21557 221 616 222 644 645 cell_1rw
* cell instance $21558 m0 *1 54.99,141.96
X$21558 221 618 222 644 645 cell_1rw
* cell instance $21559 r0 *1 54.99,141.96
X$21559 221 619 222 644 645 cell_1rw
* cell instance $21560 m0 *1 54.99,144.69
X$21560 221 620 222 644 645 cell_1rw
* cell instance $21561 r0 *1 54.99,144.69
X$21561 221 621 222 644 645 cell_1rw
* cell instance $21562 m0 *1 54.99,147.42
X$21562 221 622 222 644 645 cell_1rw
* cell instance $21563 r0 *1 54.99,147.42
X$21563 221 623 222 644 645 cell_1rw
* cell instance $21564 m0 *1 54.99,150.15
X$21564 221 624 222 644 645 cell_1rw
* cell instance $21565 m0 *1 54.99,152.88
X$21565 221 626 222 644 645 cell_1rw
* cell instance $21566 r0 *1 54.99,150.15
X$21566 221 625 222 644 645 cell_1rw
* cell instance $21567 r0 *1 54.99,152.88
X$21567 221 627 222 644 645 cell_1rw
* cell instance $21568 m0 *1 54.99,155.61
X$21568 221 628 222 644 645 cell_1rw
* cell instance $21569 r0 *1 54.99,155.61
X$21569 221 629 222 644 645 cell_1rw
* cell instance $21570 m0 *1 54.99,158.34
X$21570 221 630 222 644 645 cell_1rw
* cell instance $21571 r0 *1 54.99,158.34
X$21571 221 631 222 644 645 cell_1rw
* cell instance $21572 m0 *1 54.99,161.07
X$21572 221 632 222 644 645 cell_1rw
* cell instance $21573 r0 *1 54.99,161.07
X$21573 221 633 222 644 645 cell_1rw
* cell instance $21574 m0 *1 54.99,163.8
X$21574 221 634 222 644 645 cell_1rw
* cell instance $21575 r0 *1 54.99,163.8
X$21575 221 635 222 644 645 cell_1rw
* cell instance $21576 m0 *1 54.99,166.53
X$21576 221 637 222 644 645 cell_1rw
* cell instance $21577 m0 *1 54.99,169.26
X$21577 221 639 222 644 645 cell_1rw
* cell instance $21578 r0 *1 54.99,166.53
X$21578 221 636 222 644 645 cell_1rw
* cell instance $21579 r0 *1 54.99,169.26
X$21579 221 638 222 644 645 cell_1rw
* cell instance $21580 m0 *1 54.99,171.99
X$21580 221 640 222 644 645 cell_1rw
* cell instance $21581 r0 *1 54.99,171.99
X$21581 221 641 222 644 645 cell_1rw
* cell instance $21582 m0 *1 54.99,174.72
X$21582 221 642 222 644 645 cell_1rw
* cell instance $21583 r0 *1 54.99,174.72
X$21583 221 643 222 644 645 cell_1rw
* cell instance $21584 r0 *1 55.695,87.36
X$21584 223 322 224 644 645 cell_1rw
* cell instance $21585 m0 *1 55.695,90.09
X$21585 223 581 224 644 645 cell_1rw
* cell instance $21586 r0 *1 55.695,90.09
X$21586 223 580 224 644 645 cell_1rw
* cell instance $21587 m0 *1 55.695,92.82
X$21587 223 583 224 644 645 cell_1rw
* cell instance $21588 m0 *1 55.695,95.55
X$21588 223 584 224 644 645 cell_1rw
* cell instance $21589 r0 *1 55.695,92.82
X$21589 223 582 224 644 645 cell_1rw
* cell instance $21590 r0 *1 55.695,95.55
X$21590 223 585 224 644 645 cell_1rw
* cell instance $21591 m0 *1 55.695,98.28
X$21591 223 586 224 644 645 cell_1rw
* cell instance $21592 r0 *1 55.695,98.28
X$21592 223 587 224 644 645 cell_1rw
* cell instance $21593 m0 *1 55.695,101.01
X$21593 223 588 224 644 645 cell_1rw
* cell instance $21594 r0 *1 55.695,101.01
X$21594 223 589 224 644 645 cell_1rw
* cell instance $21595 m0 *1 55.695,103.74
X$21595 223 590 224 644 645 cell_1rw
* cell instance $21596 r0 *1 55.695,103.74
X$21596 223 591 224 644 645 cell_1rw
* cell instance $21597 m0 *1 55.695,106.47
X$21597 223 593 224 644 645 cell_1rw
* cell instance $21598 r0 *1 55.695,106.47
X$21598 223 592 224 644 645 cell_1rw
* cell instance $21599 m0 *1 55.695,109.2
X$21599 223 594 224 644 645 cell_1rw
* cell instance $21600 r0 *1 55.695,109.2
X$21600 223 595 224 644 645 cell_1rw
* cell instance $21601 m0 *1 55.695,111.93
X$21601 223 597 224 644 645 cell_1rw
* cell instance $21602 r0 *1 55.695,111.93
X$21602 223 596 224 644 645 cell_1rw
* cell instance $21603 m0 *1 55.695,114.66
X$21603 223 598 224 644 645 cell_1rw
* cell instance $21604 r0 *1 55.695,114.66
X$21604 223 599 224 644 645 cell_1rw
* cell instance $21605 m0 *1 55.695,117.39
X$21605 223 600 224 644 645 cell_1rw
* cell instance $21606 r0 *1 55.695,117.39
X$21606 223 601 224 644 645 cell_1rw
* cell instance $21607 m0 *1 55.695,120.12
X$21607 223 602 224 644 645 cell_1rw
* cell instance $21608 r0 *1 55.695,120.12
X$21608 223 603 224 644 645 cell_1rw
* cell instance $21609 m0 *1 55.695,122.85
X$21609 223 604 224 644 645 cell_1rw
* cell instance $21610 m0 *1 55.695,125.58
X$21610 223 606 224 644 645 cell_1rw
* cell instance $21611 r0 *1 55.695,122.85
X$21611 223 605 224 644 645 cell_1rw
* cell instance $21612 r0 *1 55.695,125.58
X$21612 223 607 224 644 645 cell_1rw
* cell instance $21613 m0 *1 55.695,128.31
X$21613 223 609 224 644 645 cell_1rw
* cell instance $21614 r0 *1 55.695,128.31
X$21614 223 608 224 644 645 cell_1rw
* cell instance $21615 m0 *1 55.695,131.04
X$21615 223 610 224 644 645 cell_1rw
* cell instance $21616 r0 *1 55.695,131.04
X$21616 223 611 224 644 645 cell_1rw
* cell instance $21617 m0 *1 55.695,133.77
X$21617 223 612 224 644 645 cell_1rw
* cell instance $21618 r0 *1 55.695,133.77
X$21618 223 613 224 644 645 cell_1rw
* cell instance $21619 m0 *1 55.695,136.5
X$21619 223 615 224 644 645 cell_1rw
* cell instance $21620 r0 *1 55.695,136.5
X$21620 223 614 224 644 645 cell_1rw
* cell instance $21621 m0 *1 55.695,139.23
X$21621 223 617 224 644 645 cell_1rw
* cell instance $21622 r0 *1 55.695,139.23
X$21622 223 616 224 644 645 cell_1rw
* cell instance $21623 m0 *1 55.695,141.96
X$21623 223 618 224 644 645 cell_1rw
* cell instance $21624 r0 *1 55.695,141.96
X$21624 223 619 224 644 645 cell_1rw
* cell instance $21625 m0 *1 55.695,144.69
X$21625 223 620 224 644 645 cell_1rw
* cell instance $21626 m0 *1 55.695,147.42
X$21626 223 622 224 644 645 cell_1rw
* cell instance $21627 r0 *1 55.695,144.69
X$21627 223 621 224 644 645 cell_1rw
* cell instance $21628 r0 *1 55.695,147.42
X$21628 223 623 224 644 645 cell_1rw
* cell instance $21629 m0 *1 55.695,150.15
X$21629 223 624 224 644 645 cell_1rw
* cell instance $21630 r0 *1 55.695,150.15
X$21630 223 625 224 644 645 cell_1rw
* cell instance $21631 m0 *1 55.695,152.88
X$21631 223 626 224 644 645 cell_1rw
* cell instance $21632 r0 *1 55.695,152.88
X$21632 223 627 224 644 645 cell_1rw
* cell instance $21633 m0 *1 55.695,155.61
X$21633 223 628 224 644 645 cell_1rw
* cell instance $21634 r0 *1 55.695,155.61
X$21634 223 629 224 644 645 cell_1rw
* cell instance $21635 m0 *1 55.695,158.34
X$21635 223 630 224 644 645 cell_1rw
* cell instance $21636 r0 *1 55.695,158.34
X$21636 223 631 224 644 645 cell_1rw
* cell instance $21637 m0 *1 55.695,161.07
X$21637 223 632 224 644 645 cell_1rw
* cell instance $21638 m0 *1 55.695,163.8
X$21638 223 634 224 644 645 cell_1rw
* cell instance $21639 r0 *1 55.695,161.07
X$21639 223 633 224 644 645 cell_1rw
* cell instance $21640 r0 *1 55.695,163.8
X$21640 223 635 224 644 645 cell_1rw
* cell instance $21641 m0 *1 55.695,166.53
X$21641 223 637 224 644 645 cell_1rw
* cell instance $21642 r0 *1 55.695,166.53
X$21642 223 636 224 644 645 cell_1rw
* cell instance $21643 m0 *1 55.695,169.26
X$21643 223 639 224 644 645 cell_1rw
* cell instance $21644 r0 *1 55.695,169.26
X$21644 223 638 224 644 645 cell_1rw
* cell instance $21645 m0 *1 55.695,171.99
X$21645 223 640 224 644 645 cell_1rw
* cell instance $21646 r0 *1 55.695,171.99
X$21646 223 641 224 644 645 cell_1rw
* cell instance $21647 m0 *1 55.695,174.72
X$21647 223 642 224 644 645 cell_1rw
* cell instance $21648 r0 *1 55.695,174.72
X$21648 223 643 224 644 645 cell_1rw
* cell instance $21649 r0 *1 56.4,87.36
X$21649 225 322 226 644 645 cell_1rw
* cell instance $21650 m0 *1 56.4,90.09
X$21650 225 581 226 644 645 cell_1rw
* cell instance $21651 r0 *1 56.4,90.09
X$21651 225 580 226 644 645 cell_1rw
* cell instance $21652 m0 *1 56.4,92.82
X$21652 225 583 226 644 645 cell_1rw
* cell instance $21653 r0 *1 56.4,92.82
X$21653 225 582 226 644 645 cell_1rw
* cell instance $21654 m0 *1 56.4,95.55
X$21654 225 584 226 644 645 cell_1rw
* cell instance $21655 r0 *1 56.4,95.55
X$21655 225 585 226 644 645 cell_1rw
* cell instance $21656 m0 *1 56.4,98.28
X$21656 225 586 226 644 645 cell_1rw
* cell instance $21657 r0 *1 56.4,98.28
X$21657 225 587 226 644 645 cell_1rw
* cell instance $21658 m0 *1 56.4,101.01
X$21658 225 588 226 644 645 cell_1rw
* cell instance $21659 r0 *1 56.4,101.01
X$21659 225 589 226 644 645 cell_1rw
* cell instance $21660 m0 *1 56.4,103.74
X$21660 225 590 226 644 645 cell_1rw
* cell instance $21661 m0 *1 56.4,106.47
X$21661 225 593 226 644 645 cell_1rw
* cell instance $21662 r0 *1 56.4,103.74
X$21662 225 591 226 644 645 cell_1rw
* cell instance $21663 r0 *1 56.4,106.47
X$21663 225 592 226 644 645 cell_1rw
* cell instance $21664 m0 *1 56.4,109.2
X$21664 225 594 226 644 645 cell_1rw
* cell instance $21665 r0 *1 56.4,109.2
X$21665 225 595 226 644 645 cell_1rw
* cell instance $21666 m0 *1 56.4,111.93
X$21666 225 597 226 644 645 cell_1rw
* cell instance $21667 r0 *1 56.4,111.93
X$21667 225 596 226 644 645 cell_1rw
* cell instance $21668 m0 *1 56.4,114.66
X$21668 225 598 226 644 645 cell_1rw
* cell instance $21669 r0 *1 56.4,114.66
X$21669 225 599 226 644 645 cell_1rw
* cell instance $21670 m0 *1 56.4,117.39
X$21670 225 600 226 644 645 cell_1rw
* cell instance $21671 r0 *1 56.4,117.39
X$21671 225 601 226 644 645 cell_1rw
* cell instance $21672 m0 *1 56.4,120.12
X$21672 225 602 226 644 645 cell_1rw
* cell instance $21673 m0 *1 56.4,122.85
X$21673 225 604 226 644 645 cell_1rw
* cell instance $21674 r0 *1 56.4,120.12
X$21674 225 603 226 644 645 cell_1rw
* cell instance $21675 r0 *1 56.4,122.85
X$21675 225 605 226 644 645 cell_1rw
* cell instance $21676 m0 *1 56.4,125.58
X$21676 225 606 226 644 645 cell_1rw
* cell instance $21677 m0 *1 56.4,128.31
X$21677 225 609 226 644 645 cell_1rw
* cell instance $21678 r0 *1 56.4,125.58
X$21678 225 607 226 644 645 cell_1rw
* cell instance $21679 r0 *1 56.4,128.31
X$21679 225 608 226 644 645 cell_1rw
* cell instance $21680 m0 *1 56.4,131.04
X$21680 225 610 226 644 645 cell_1rw
* cell instance $21681 r0 *1 56.4,131.04
X$21681 225 611 226 644 645 cell_1rw
* cell instance $21682 m0 *1 56.4,133.77
X$21682 225 612 226 644 645 cell_1rw
* cell instance $21683 r0 *1 56.4,133.77
X$21683 225 613 226 644 645 cell_1rw
* cell instance $21684 m0 *1 56.4,136.5
X$21684 225 615 226 644 645 cell_1rw
* cell instance $21685 r0 *1 56.4,136.5
X$21685 225 614 226 644 645 cell_1rw
* cell instance $21686 m0 *1 56.4,139.23
X$21686 225 617 226 644 645 cell_1rw
* cell instance $21687 r0 *1 56.4,139.23
X$21687 225 616 226 644 645 cell_1rw
* cell instance $21688 m0 *1 56.4,141.96
X$21688 225 618 226 644 645 cell_1rw
* cell instance $21689 r0 *1 56.4,141.96
X$21689 225 619 226 644 645 cell_1rw
* cell instance $21690 m0 *1 56.4,144.69
X$21690 225 620 226 644 645 cell_1rw
* cell instance $21691 r0 *1 56.4,144.69
X$21691 225 621 226 644 645 cell_1rw
* cell instance $21692 m0 *1 56.4,147.42
X$21692 225 622 226 644 645 cell_1rw
* cell instance $21693 m0 *1 56.4,150.15
X$21693 225 624 226 644 645 cell_1rw
* cell instance $21694 r0 *1 56.4,147.42
X$21694 225 623 226 644 645 cell_1rw
* cell instance $21695 r0 *1 56.4,150.15
X$21695 225 625 226 644 645 cell_1rw
* cell instance $21696 m0 *1 56.4,152.88
X$21696 225 626 226 644 645 cell_1rw
* cell instance $21697 r0 *1 56.4,152.88
X$21697 225 627 226 644 645 cell_1rw
* cell instance $21698 m0 *1 56.4,155.61
X$21698 225 628 226 644 645 cell_1rw
* cell instance $21699 r0 *1 56.4,155.61
X$21699 225 629 226 644 645 cell_1rw
* cell instance $21700 m0 *1 56.4,158.34
X$21700 225 630 226 644 645 cell_1rw
* cell instance $21701 r0 *1 56.4,158.34
X$21701 225 631 226 644 645 cell_1rw
* cell instance $21702 m0 *1 56.4,161.07
X$21702 225 632 226 644 645 cell_1rw
* cell instance $21703 r0 *1 56.4,161.07
X$21703 225 633 226 644 645 cell_1rw
* cell instance $21704 m0 *1 56.4,163.8
X$21704 225 634 226 644 645 cell_1rw
* cell instance $21705 m0 *1 56.4,166.53
X$21705 225 637 226 644 645 cell_1rw
* cell instance $21706 r0 *1 56.4,163.8
X$21706 225 635 226 644 645 cell_1rw
* cell instance $21707 r0 *1 56.4,166.53
X$21707 225 636 226 644 645 cell_1rw
* cell instance $21708 m0 *1 56.4,169.26
X$21708 225 639 226 644 645 cell_1rw
* cell instance $21709 r0 *1 56.4,169.26
X$21709 225 638 226 644 645 cell_1rw
* cell instance $21710 m0 *1 56.4,171.99
X$21710 225 640 226 644 645 cell_1rw
* cell instance $21711 r0 *1 56.4,171.99
X$21711 225 641 226 644 645 cell_1rw
* cell instance $21712 m0 *1 56.4,174.72
X$21712 225 642 226 644 645 cell_1rw
* cell instance $21713 r0 *1 56.4,174.72
X$21713 225 643 226 644 645 cell_1rw
* cell instance $21714 r0 *1 57.105,87.36
X$21714 227 322 228 644 645 cell_1rw
* cell instance $21715 m0 *1 57.105,90.09
X$21715 227 581 228 644 645 cell_1rw
* cell instance $21716 r0 *1 57.105,90.09
X$21716 227 580 228 644 645 cell_1rw
* cell instance $21717 m0 *1 57.105,92.82
X$21717 227 583 228 644 645 cell_1rw
* cell instance $21718 r0 *1 57.105,92.82
X$21718 227 582 228 644 645 cell_1rw
* cell instance $21719 m0 *1 57.105,95.55
X$21719 227 584 228 644 645 cell_1rw
* cell instance $21720 r0 *1 57.105,95.55
X$21720 227 585 228 644 645 cell_1rw
* cell instance $21721 m0 *1 57.105,98.28
X$21721 227 586 228 644 645 cell_1rw
* cell instance $21722 r0 *1 57.105,98.28
X$21722 227 587 228 644 645 cell_1rw
* cell instance $21723 m0 *1 57.105,101.01
X$21723 227 588 228 644 645 cell_1rw
* cell instance $21724 r0 *1 57.105,101.01
X$21724 227 589 228 644 645 cell_1rw
* cell instance $21725 m0 *1 57.105,103.74
X$21725 227 590 228 644 645 cell_1rw
* cell instance $21726 m0 *1 57.105,106.47
X$21726 227 593 228 644 645 cell_1rw
* cell instance $21727 r0 *1 57.105,103.74
X$21727 227 591 228 644 645 cell_1rw
* cell instance $21728 r0 *1 57.105,106.47
X$21728 227 592 228 644 645 cell_1rw
* cell instance $21729 m0 *1 57.105,109.2
X$21729 227 594 228 644 645 cell_1rw
* cell instance $21730 r0 *1 57.105,109.2
X$21730 227 595 228 644 645 cell_1rw
* cell instance $21731 m0 *1 57.105,111.93
X$21731 227 597 228 644 645 cell_1rw
* cell instance $21732 r0 *1 57.105,111.93
X$21732 227 596 228 644 645 cell_1rw
* cell instance $21733 m0 *1 57.105,114.66
X$21733 227 598 228 644 645 cell_1rw
* cell instance $21734 r0 *1 57.105,114.66
X$21734 227 599 228 644 645 cell_1rw
* cell instance $21735 m0 *1 57.105,117.39
X$21735 227 600 228 644 645 cell_1rw
* cell instance $21736 r0 *1 57.105,117.39
X$21736 227 601 228 644 645 cell_1rw
* cell instance $21737 m0 *1 57.105,120.12
X$21737 227 602 228 644 645 cell_1rw
* cell instance $21738 r0 *1 57.105,120.12
X$21738 227 603 228 644 645 cell_1rw
* cell instance $21739 m0 *1 57.105,122.85
X$21739 227 604 228 644 645 cell_1rw
* cell instance $21740 r0 *1 57.105,122.85
X$21740 227 605 228 644 645 cell_1rw
* cell instance $21741 m0 *1 57.105,125.58
X$21741 227 606 228 644 645 cell_1rw
* cell instance $21742 r0 *1 57.105,125.58
X$21742 227 607 228 644 645 cell_1rw
* cell instance $21743 m0 *1 57.105,128.31
X$21743 227 609 228 644 645 cell_1rw
* cell instance $21744 r0 *1 57.105,128.31
X$21744 227 608 228 644 645 cell_1rw
* cell instance $21745 m0 *1 57.105,131.04
X$21745 227 610 228 644 645 cell_1rw
* cell instance $21746 r0 *1 57.105,131.04
X$21746 227 611 228 644 645 cell_1rw
* cell instance $21747 m0 *1 57.105,133.77
X$21747 227 612 228 644 645 cell_1rw
* cell instance $21748 r0 *1 57.105,133.77
X$21748 227 613 228 644 645 cell_1rw
* cell instance $21749 m0 *1 57.105,136.5
X$21749 227 615 228 644 645 cell_1rw
* cell instance $21750 r0 *1 57.105,136.5
X$21750 227 614 228 644 645 cell_1rw
* cell instance $21751 m0 *1 57.105,139.23
X$21751 227 617 228 644 645 cell_1rw
* cell instance $21752 r0 *1 57.105,139.23
X$21752 227 616 228 644 645 cell_1rw
* cell instance $21753 m0 *1 57.105,141.96
X$21753 227 618 228 644 645 cell_1rw
* cell instance $21754 r0 *1 57.105,141.96
X$21754 227 619 228 644 645 cell_1rw
* cell instance $21755 m0 *1 57.105,144.69
X$21755 227 620 228 644 645 cell_1rw
* cell instance $21756 m0 *1 57.105,147.42
X$21756 227 622 228 644 645 cell_1rw
* cell instance $21757 r0 *1 57.105,144.69
X$21757 227 621 228 644 645 cell_1rw
* cell instance $21758 r0 *1 57.105,147.42
X$21758 227 623 228 644 645 cell_1rw
* cell instance $21759 m0 *1 57.105,150.15
X$21759 227 624 228 644 645 cell_1rw
* cell instance $21760 r0 *1 57.105,150.15
X$21760 227 625 228 644 645 cell_1rw
* cell instance $21761 m0 *1 57.105,152.88
X$21761 227 626 228 644 645 cell_1rw
* cell instance $21762 m0 *1 57.105,155.61
X$21762 227 628 228 644 645 cell_1rw
* cell instance $21763 r0 *1 57.105,152.88
X$21763 227 627 228 644 645 cell_1rw
* cell instance $21764 r0 *1 57.105,155.61
X$21764 227 629 228 644 645 cell_1rw
* cell instance $21765 m0 *1 57.105,158.34
X$21765 227 630 228 644 645 cell_1rw
* cell instance $21766 r0 *1 57.105,158.34
X$21766 227 631 228 644 645 cell_1rw
* cell instance $21767 m0 *1 57.105,161.07
X$21767 227 632 228 644 645 cell_1rw
* cell instance $21768 r0 *1 57.105,161.07
X$21768 227 633 228 644 645 cell_1rw
* cell instance $21769 m0 *1 57.105,163.8
X$21769 227 634 228 644 645 cell_1rw
* cell instance $21770 m0 *1 57.105,166.53
X$21770 227 637 228 644 645 cell_1rw
* cell instance $21771 r0 *1 57.105,163.8
X$21771 227 635 228 644 645 cell_1rw
* cell instance $21772 r0 *1 57.105,166.53
X$21772 227 636 228 644 645 cell_1rw
* cell instance $21773 m0 *1 57.105,169.26
X$21773 227 639 228 644 645 cell_1rw
* cell instance $21774 r0 *1 57.105,169.26
X$21774 227 638 228 644 645 cell_1rw
* cell instance $21775 m0 *1 57.105,171.99
X$21775 227 640 228 644 645 cell_1rw
* cell instance $21776 r0 *1 57.105,171.99
X$21776 227 641 228 644 645 cell_1rw
* cell instance $21777 m0 *1 57.105,174.72
X$21777 227 642 228 644 645 cell_1rw
* cell instance $21778 r0 *1 57.105,174.72
X$21778 227 643 228 644 645 cell_1rw
* cell instance $21779 r0 *1 57.81,87.36
X$21779 229 322 230 644 645 cell_1rw
* cell instance $21780 m0 *1 57.81,90.09
X$21780 229 581 230 644 645 cell_1rw
* cell instance $21781 r0 *1 57.81,90.09
X$21781 229 580 230 644 645 cell_1rw
* cell instance $21782 m0 *1 57.81,92.82
X$21782 229 583 230 644 645 cell_1rw
* cell instance $21783 r0 *1 57.81,92.82
X$21783 229 582 230 644 645 cell_1rw
* cell instance $21784 m0 *1 57.81,95.55
X$21784 229 584 230 644 645 cell_1rw
* cell instance $21785 r0 *1 57.81,95.55
X$21785 229 585 230 644 645 cell_1rw
* cell instance $21786 m0 *1 57.81,98.28
X$21786 229 586 230 644 645 cell_1rw
* cell instance $21787 r0 *1 57.81,98.28
X$21787 229 587 230 644 645 cell_1rw
* cell instance $21788 m0 *1 57.81,101.01
X$21788 229 588 230 644 645 cell_1rw
* cell instance $21789 r0 *1 57.81,101.01
X$21789 229 589 230 644 645 cell_1rw
* cell instance $21790 m0 *1 57.81,103.74
X$21790 229 590 230 644 645 cell_1rw
* cell instance $21791 r0 *1 57.81,103.74
X$21791 229 591 230 644 645 cell_1rw
* cell instance $21792 m0 *1 57.81,106.47
X$21792 229 593 230 644 645 cell_1rw
* cell instance $21793 r0 *1 57.81,106.47
X$21793 229 592 230 644 645 cell_1rw
* cell instance $21794 m0 *1 57.81,109.2
X$21794 229 594 230 644 645 cell_1rw
* cell instance $21795 r0 *1 57.81,109.2
X$21795 229 595 230 644 645 cell_1rw
* cell instance $21796 m0 *1 57.81,111.93
X$21796 229 597 230 644 645 cell_1rw
* cell instance $21797 r0 *1 57.81,111.93
X$21797 229 596 230 644 645 cell_1rw
* cell instance $21798 m0 *1 57.81,114.66
X$21798 229 598 230 644 645 cell_1rw
* cell instance $21799 r0 *1 57.81,114.66
X$21799 229 599 230 644 645 cell_1rw
* cell instance $21800 m0 *1 57.81,117.39
X$21800 229 600 230 644 645 cell_1rw
* cell instance $21801 r0 *1 57.81,117.39
X$21801 229 601 230 644 645 cell_1rw
* cell instance $21802 m0 *1 57.81,120.12
X$21802 229 602 230 644 645 cell_1rw
* cell instance $21803 r0 *1 57.81,120.12
X$21803 229 603 230 644 645 cell_1rw
* cell instance $21804 m0 *1 57.81,122.85
X$21804 229 604 230 644 645 cell_1rw
* cell instance $21805 r0 *1 57.81,122.85
X$21805 229 605 230 644 645 cell_1rw
* cell instance $21806 m0 *1 57.81,125.58
X$21806 229 606 230 644 645 cell_1rw
* cell instance $21807 r0 *1 57.81,125.58
X$21807 229 607 230 644 645 cell_1rw
* cell instance $21808 m0 *1 57.81,128.31
X$21808 229 609 230 644 645 cell_1rw
* cell instance $21809 r0 *1 57.81,128.31
X$21809 229 608 230 644 645 cell_1rw
* cell instance $21810 m0 *1 57.81,131.04
X$21810 229 610 230 644 645 cell_1rw
* cell instance $21811 r0 *1 57.81,131.04
X$21811 229 611 230 644 645 cell_1rw
* cell instance $21812 m0 *1 57.81,133.77
X$21812 229 612 230 644 645 cell_1rw
* cell instance $21813 r0 *1 57.81,133.77
X$21813 229 613 230 644 645 cell_1rw
* cell instance $21814 m0 *1 57.81,136.5
X$21814 229 615 230 644 645 cell_1rw
* cell instance $21815 m0 *1 57.81,139.23
X$21815 229 617 230 644 645 cell_1rw
* cell instance $21816 r0 *1 57.81,136.5
X$21816 229 614 230 644 645 cell_1rw
* cell instance $21817 m0 *1 57.81,141.96
X$21817 229 618 230 644 645 cell_1rw
* cell instance $21818 r0 *1 57.81,139.23
X$21818 229 616 230 644 645 cell_1rw
* cell instance $21819 r0 *1 57.81,141.96
X$21819 229 619 230 644 645 cell_1rw
* cell instance $21820 m0 *1 57.81,144.69
X$21820 229 620 230 644 645 cell_1rw
* cell instance $21821 m0 *1 57.81,147.42
X$21821 229 622 230 644 645 cell_1rw
* cell instance $21822 r0 *1 57.81,144.69
X$21822 229 621 230 644 645 cell_1rw
* cell instance $21823 r0 *1 57.81,147.42
X$21823 229 623 230 644 645 cell_1rw
* cell instance $21824 m0 *1 57.81,150.15
X$21824 229 624 230 644 645 cell_1rw
* cell instance $21825 m0 *1 57.81,152.88
X$21825 229 626 230 644 645 cell_1rw
* cell instance $21826 r0 *1 57.81,150.15
X$21826 229 625 230 644 645 cell_1rw
* cell instance $21827 r0 *1 57.81,152.88
X$21827 229 627 230 644 645 cell_1rw
* cell instance $21828 m0 *1 57.81,155.61
X$21828 229 628 230 644 645 cell_1rw
* cell instance $21829 r0 *1 57.81,155.61
X$21829 229 629 230 644 645 cell_1rw
* cell instance $21830 m0 *1 57.81,158.34
X$21830 229 630 230 644 645 cell_1rw
* cell instance $21831 r0 *1 57.81,158.34
X$21831 229 631 230 644 645 cell_1rw
* cell instance $21832 m0 *1 57.81,161.07
X$21832 229 632 230 644 645 cell_1rw
* cell instance $21833 r0 *1 57.81,161.07
X$21833 229 633 230 644 645 cell_1rw
* cell instance $21834 m0 *1 57.81,163.8
X$21834 229 634 230 644 645 cell_1rw
* cell instance $21835 r0 *1 57.81,163.8
X$21835 229 635 230 644 645 cell_1rw
* cell instance $21836 m0 *1 57.81,166.53
X$21836 229 637 230 644 645 cell_1rw
* cell instance $21837 r0 *1 57.81,166.53
X$21837 229 636 230 644 645 cell_1rw
* cell instance $21838 m0 *1 57.81,169.26
X$21838 229 639 230 644 645 cell_1rw
* cell instance $21839 r0 *1 57.81,169.26
X$21839 229 638 230 644 645 cell_1rw
* cell instance $21840 m0 *1 57.81,171.99
X$21840 229 640 230 644 645 cell_1rw
* cell instance $21841 r0 *1 57.81,171.99
X$21841 229 641 230 644 645 cell_1rw
* cell instance $21842 m0 *1 57.81,174.72
X$21842 229 642 230 644 645 cell_1rw
* cell instance $21843 r0 *1 57.81,174.72
X$21843 229 643 230 644 645 cell_1rw
* cell instance $21844 r0 *1 58.515,87.36
X$21844 231 322 232 644 645 cell_1rw
* cell instance $21845 m0 *1 58.515,90.09
X$21845 231 581 232 644 645 cell_1rw
* cell instance $21846 r0 *1 58.515,90.09
X$21846 231 580 232 644 645 cell_1rw
* cell instance $21847 m0 *1 58.515,92.82
X$21847 231 583 232 644 645 cell_1rw
* cell instance $21848 r0 *1 58.515,92.82
X$21848 231 582 232 644 645 cell_1rw
* cell instance $21849 m0 *1 58.515,95.55
X$21849 231 584 232 644 645 cell_1rw
* cell instance $21850 r0 *1 58.515,95.55
X$21850 231 585 232 644 645 cell_1rw
* cell instance $21851 m0 *1 58.515,98.28
X$21851 231 586 232 644 645 cell_1rw
* cell instance $21852 r0 *1 58.515,98.28
X$21852 231 587 232 644 645 cell_1rw
* cell instance $21853 m0 *1 58.515,101.01
X$21853 231 588 232 644 645 cell_1rw
* cell instance $21854 r0 *1 58.515,101.01
X$21854 231 589 232 644 645 cell_1rw
* cell instance $21855 m0 *1 58.515,103.74
X$21855 231 590 232 644 645 cell_1rw
* cell instance $21856 r0 *1 58.515,103.74
X$21856 231 591 232 644 645 cell_1rw
* cell instance $21857 m0 *1 58.515,106.47
X$21857 231 593 232 644 645 cell_1rw
* cell instance $21858 r0 *1 58.515,106.47
X$21858 231 592 232 644 645 cell_1rw
* cell instance $21859 m0 *1 58.515,109.2
X$21859 231 594 232 644 645 cell_1rw
* cell instance $21860 r0 *1 58.515,109.2
X$21860 231 595 232 644 645 cell_1rw
* cell instance $21861 m0 *1 58.515,111.93
X$21861 231 597 232 644 645 cell_1rw
* cell instance $21862 r0 *1 58.515,111.93
X$21862 231 596 232 644 645 cell_1rw
* cell instance $21863 m0 *1 58.515,114.66
X$21863 231 598 232 644 645 cell_1rw
* cell instance $21864 r0 *1 58.515,114.66
X$21864 231 599 232 644 645 cell_1rw
* cell instance $21865 m0 *1 58.515,117.39
X$21865 231 600 232 644 645 cell_1rw
* cell instance $21866 r0 *1 58.515,117.39
X$21866 231 601 232 644 645 cell_1rw
* cell instance $21867 m0 *1 58.515,120.12
X$21867 231 602 232 644 645 cell_1rw
* cell instance $21868 r0 *1 58.515,120.12
X$21868 231 603 232 644 645 cell_1rw
* cell instance $21869 m0 *1 58.515,122.85
X$21869 231 604 232 644 645 cell_1rw
* cell instance $21870 r0 *1 58.515,122.85
X$21870 231 605 232 644 645 cell_1rw
* cell instance $21871 m0 *1 58.515,125.58
X$21871 231 606 232 644 645 cell_1rw
* cell instance $21872 m0 *1 58.515,128.31
X$21872 231 609 232 644 645 cell_1rw
* cell instance $21873 r0 *1 58.515,125.58
X$21873 231 607 232 644 645 cell_1rw
* cell instance $21874 r0 *1 58.515,128.31
X$21874 231 608 232 644 645 cell_1rw
* cell instance $21875 m0 *1 58.515,131.04
X$21875 231 610 232 644 645 cell_1rw
* cell instance $21876 r0 *1 58.515,131.04
X$21876 231 611 232 644 645 cell_1rw
* cell instance $21877 m0 *1 58.515,133.77
X$21877 231 612 232 644 645 cell_1rw
* cell instance $21878 r0 *1 58.515,133.77
X$21878 231 613 232 644 645 cell_1rw
* cell instance $21879 m0 *1 58.515,136.5
X$21879 231 615 232 644 645 cell_1rw
* cell instance $21880 r0 *1 58.515,136.5
X$21880 231 614 232 644 645 cell_1rw
* cell instance $21881 m0 *1 58.515,139.23
X$21881 231 617 232 644 645 cell_1rw
* cell instance $21882 r0 *1 58.515,139.23
X$21882 231 616 232 644 645 cell_1rw
* cell instance $21883 m0 *1 58.515,141.96
X$21883 231 618 232 644 645 cell_1rw
* cell instance $21884 r0 *1 58.515,141.96
X$21884 231 619 232 644 645 cell_1rw
* cell instance $21885 m0 *1 58.515,144.69
X$21885 231 620 232 644 645 cell_1rw
* cell instance $21886 r0 *1 58.515,144.69
X$21886 231 621 232 644 645 cell_1rw
* cell instance $21887 m0 *1 58.515,147.42
X$21887 231 622 232 644 645 cell_1rw
* cell instance $21888 r0 *1 58.515,147.42
X$21888 231 623 232 644 645 cell_1rw
* cell instance $21889 m0 *1 58.515,150.15
X$21889 231 624 232 644 645 cell_1rw
* cell instance $21890 r0 *1 58.515,150.15
X$21890 231 625 232 644 645 cell_1rw
* cell instance $21891 m0 *1 58.515,152.88
X$21891 231 626 232 644 645 cell_1rw
* cell instance $21892 r0 *1 58.515,152.88
X$21892 231 627 232 644 645 cell_1rw
* cell instance $21893 m0 *1 58.515,155.61
X$21893 231 628 232 644 645 cell_1rw
* cell instance $21894 m0 *1 58.515,158.34
X$21894 231 630 232 644 645 cell_1rw
* cell instance $21895 r0 *1 58.515,155.61
X$21895 231 629 232 644 645 cell_1rw
* cell instance $21896 m0 *1 58.515,161.07
X$21896 231 632 232 644 645 cell_1rw
* cell instance $21897 r0 *1 58.515,158.34
X$21897 231 631 232 644 645 cell_1rw
* cell instance $21898 r0 *1 58.515,161.07
X$21898 231 633 232 644 645 cell_1rw
* cell instance $21899 m0 *1 58.515,163.8
X$21899 231 634 232 644 645 cell_1rw
* cell instance $21900 r0 *1 58.515,163.8
X$21900 231 635 232 644 645 cell_1rw
* cell instance $21901 m0 *1 58.515,166.53
X$21901 231 637 232 644 645 cell_1rw
* cell instance $21902 r0 *1 58.515,166.53
X$21902 231 636 232 644 645 cell_1rw
* cell instance $21903 m0 *1 58.515,169.26
X$21903 231 639 232 644 645 cell_1rw
* cell instance $21904 r0 *1 58.515,169.26
X$21904 231 638 232 644 645 cell_1rw
* cell instance $21905 m0 *1 58.515,171.99
X$21905 231 640 232 644 645 cell_1rw
* cell instance $21906 r0 *1 58.515,171.99
X$21906 231 641 232 644 645 cell_1rw
* cell instance $21907 m0 *1 58.515,174.72
X$21907 231 642 232 644 645 cell_1rw
* cell instance $21908 r0 *1 58.515,174.72
X$21908 231 643 232 644 645 cell_1rw
* cell instance $21909 r0 *1 59.22,87.36
X$21909 233 322 234 644 645 cell_1rw
* cell instance $21910 m0 *1 59.22,90.09
X$21910 233 581 234 644 645 cell_1rw
* cell instance $21911 m0 *1 59.22,92.82
X$21911 233 583 234 644 645 cell_1rw
* cell instance $21912 r0 *1 59.22,90.09
X$21912 233 580 234 644 645 cell_1rw
* cell instance $21913 r0 *1 59.22,92.82
X$21913 233 582 234 644 645 cell_1rw
* cell instance $21914 m0 *1 59.22,95.55
X$21914 233 584 234 644 645 cell_1rw
* cell instance $21915 r0 *1 59.22,95.55
X$21915 233 585 234 644 645 cell_1rw
* cell instance $21916 m0 *1 59.22,98.28
X$21916 233 586 234 644 645 cell_1rw
* cell instance $21917 m0 *1 59.22,101.01
X$21917 233 588 234 644 645 cell_1rw
* cell instance $21918 r0 *1 59.22,98.28
X$21918 233 587 234 644 645 cell_1rw
* cell instance $21919 m0 *1 59.22,103.74
X$21919 233 590 234 644 645 cell_1rw
* cell instance $21920 r0 *1 59.22,101.01
X$21920 233 589 234 644 645 cell_1rw
* cell instance $21921 r0 *1 59.22,103.74
X$21921 233 591 234 644 645 cell_1rw
* cell instance $21922 m0 *1 59.22,106.47
X$21922 233 593 234 644 645 cell_1rw
* cell instance $21923 r0 *1 59.22,106.47
X$21923 233 592 234 644 645 cell_1rw
* cell instance $21924 m0 *1 59.22,109.2
X$21924 233 594 234 644 645 cell_1rw
* cell instance $21925 r0 *1 59.22,109.2
X$21925 233 595 234 644 645 cell_1rw
* cell instance $21926 m0 *1 59.22,111.93
X$21926 233 597 234 644 645 cell_1rw
* cell instance $21927 r0 *1 59.22,111.93
X$21927 233 596 234 644 645 cell_1rw
* cell instance $21928 m0 *1 59.22,114.66
X$21928 233 598 234 644 645 cell_1rw
* cell instance $21929 r0 *1 59.22,114.66
X$21929 233 599 234 644 645 cell_1rw
* cell instance $21930 m0 *1 59.22,117.39
X$21930 233 600 234 644 645 cell_1rw
* cell instance $21931 r0 *1 59.22,117.39
X$21931 233 601 234 644 645 cell_1rw
* cell instance $21932 m0 *1 59.22,120.12
X$21932 233 602 234 644 645 cell_1rw
* cell instance $21933 r0 *1 59.22,120.12
X$21933 233 603 234 644 645 cell_1rw
* cell instance $21934 m0 *1 59.22,122.85
X$21934 233 604 234 644 645 cell_1rw
* cell instance $21935 r0 *1 59.22,122.85
X$21935 233 605 234 644 645 cell_1rw
* cell instance $21936 m0 *1 59.22,125.58
X$21936 233 606 234 644 645 cell_1rw
* cell instance $21937 r0 *1 59.22,125.58
X$21937 233 607 234 644 645 cell_1rw
* cell instance $21938 m0 *1 59.22,128.31
X$21938 233 609 234 644 645 cell_1rw
* cell instance $21939 r0 *1 59.22,128.31
X$21939 233 608 234 644 645 cell_1rw
* cell instance $21940 m0 *1 59.22,131.04
X$21940 233 610 234 644 645 cell_1rw
* cell instance $21941 m0 *1 59.22,133.77
X$21941 233 612 234 644 645 cell_1rw
* cell instance $21942 r0 *1 59.22,131.04
X$21942 233 611 234 644 645 cell_1rw
* cell instance $21943 r0 *1 59.22,133.77
X$21943 233 613 234 644 645 cell_1rw
* cell instance $21944 m0 *1 59.22,136.5
X$21944 233 615 234 644 645 cell_1rw
* cell instance $21945 r0 *1 59.22,136.5
X$21945 233 614 234 644 645 cell_1rw
* cell instance $21946 m0 *1 59.22,139.23
X$21946 233 617 234 644 645 cell_1rw
* cell instance $21947 r0 *1 59.22,139.23
X$21947 233 616 234 644 645 cell_1rw
* cell instance $21948 m0 *1 59.22,141.96
X$21948 233 618 234 644 645 cell_1rw
* cell instance $21949 r0 *1 59.22,141.96
X$21949 233 619 234 644 645 cell_1rw
* cell instance $21950 m0 *1 59.22,144.69
X$21950 233 620 234 644 645 cell_1rw
* cell instance $21951 r0 *1 59.22,144.69
X$21951 233 621 234 644 645 cell_1rw
* cell instance $21952 m0 *1 59.22,147.42
X$21952 233 622 234 644 645 cell_1rw
* cell instance $21953 r0 *1 59.22,147.42
X$21953 233 623 234 644 645 cell_1rw
* cell instance $21954 m0 *1 59.22,150.15
X$21954 233 624 234 644 645 cell_1rw
* cell instance $21955 r0 *1 59.22,150.15
X$21955 233 625 234 644 645 cell_1rw
* cell instance $21956 m0 *1 59.22,152.88
X$21956 233 626 234 644 645 cell_1rw
* cell instance $21957 r0 *1 59.22,152.88
X$21957 233 627 234 644 645 cell_1rw
* cell instance $21958 m0 *1 59.22,155.61
X$21958 233 628 234 644 645 cell_1rw
* cell instance $21959 r0 *1 59.22,155.61
X$21959 233 629 234 644 645 cell_1rw
* cell instance $21960 m0 *1 59.22,158.34
X$21960 233 630 234 644 645 cell_1rw
* cell instance $21961 r0 *1 59.22,158.34
X$21961 233 631 234 644 645 cell_1rw
* cell instance $21962 m0 *1 59.22,161.07
X$21962 233 632 234 644 645 cell_1rw
* cell instance $21963 r0 *1 59.22,161.07
X$21963 233 633 234 644 645 cell_1rw
* cell instance $21964 m0 *1 59.22,163.8
X$21964 233 634 234 644 645 cell_1rw
* cell instance $21965 r0 *1 59.22,163.8
X$21965 233 635 234 644 645 cell_1rw
* cell instance $21966 m0 *1 59.22,166.53
X$21966 233 637 234 644 645 cell_1rw
* cell instance $21967 m0 *1 59.22,169.26
X$21967 233 639 234 644 645 cell_1rw
* cell instance $21968 r0 *1 59.22,166.53
X$21968 233 636 234 644 645 cell_1rw
* cell instance $21969 r0 *1 59.22,169.26
X$21969 233 638 234 644 645 cell_1rw
* cell instance $21970 m0 *1 59.22,171.99
X$21970 233 640 234 644 645 cell_1rw
* cell instance $21971 r0 *1 59.22,171.99
X$21971 233 641 234 644 645 cell_1rw
* cell instance $21972 m0 *1 59.22,174.72
X$21972 233 642 234 644 645 cell_1rw
* cell instance $21973 r0 *1 59.22,174.72
X$21973 233 643 234 644 645 cell_1rw
* cell instance $21974 r0 *1 59.925,87.36
X$21974 235 322 236 644 645 cell_1rw
* cell instance $21975 m0 *1 59.925,90.09
X$21975 235 581 236 644 645 cell_1rw
* cell instance $21976 r0 *1 59.925,90.09
X$21976 235 580 236 644 645 cell_1rw
* cell instance $21977 m0 *1 59.925,92.82
X$21977 235 583 236 644 645 cell_1rw
* cell instance $21978 r0 *1 59.925,92.82
X$21978 235 582 236 644 645 cell_1rw
* cell instance $21979 m0 *1 59.925,95.55
X$21979 235 584 236 644 645 cell_1rw
* cell instance $21980 r0 *1 59.925,95.55
X$21980 235 585 236 644 645 cell_1rw
* cell instance $21981 m0 *1 59.925,98.28
X$21981 235 586 236 644 645 cell_1rw
* cell instance $21982 r0 *1 59.925,98.28
X$21982 235 587 236 644 645 cell_1rw
* cell instance $21983 m0 *1 59.925,101.01
X$21983 235 588 236 644 645 cell_1rw
* cell instance $21984 r0 *1 59.925,101.01
X$21984 235 589 236 644 645 cell_1rw
* cell instance $21985 m0 *1 59.925,103.74
X$21985 235 590 236 644 645 cell_1rw
* cell instance $21986 r0 *1 59.925,103.74
X$21986 235 591 236 644 645 cell_1rw
* cell instance $21987 m0 *1 59.925,106.47
X$21987 235 593 236 644 645 cell_1rw
* cell instance $21988 r0 *1 59.925,106.47
X$21988 235 592 236 644 645 cell_1rw
* cell instance $21989 m0 *1 59.925,109.2
X$21989 235 594 236 644 645 cell_1rw
* cell instance $21990 m0 *1 59.925,111.93
X$21990 235 597 236 644 645 cell_1rw
* cell instance $21991 r0 *1 59.925,109.2
X$21991 235 595 236 644 645 cell_1rw
* cell instance $21992 m0 *1 59.925,114.66
X$21992 235 598 236 644 645 cell_1rw
* cell instance $21993 r0 *1 59.925,111.93
X$21993 235 596 236 644 645 cell_1rw
* cell instance $21994 r0 *1 59.925,114.66
X$21994 235 599 236 644 645 cell_1rw
* cell instance $21995 m0 *1 59.925,117.39
X$21995 235 600 236 644 645 cell_1rw
* cell instance $21996 r0 *1 59.925,117.39
X$21996 235 601 236 644 645 cell_1rw
* cell instance $21997 m0 *1 59.925,120.12
X$21997 235 602 236 644 645 cell_1rw
* cell instance $21998 r0 *1 59.925,120.12
X$21998 235 603 236 644 645 cell_1rw
* cell instance $21999 m0 *1 59.925,122.85
X$21999 235 604 236 644 645 cell_1rw
* cell instance $22000 m0 *1 59.925,125.58
X$22000 235 606 236 644 645 cell_1rw
* cell instance $22001 r0 *1 59.925,122.85
X$22001 235 605 236 644 645 cell_1rw
* cell instance $22002 r0 *1 59.925,125.58
X$22002 235 607 236 644 645 cell_1rw
* cell instance $22003 m0 *1 59.925,128.31
X$22003 235 609 236 644 645 cell_1rw
* cell instance $22004 r0 *1 59.925,128.31
X$22004 235 608 236 644 645 cell_1rw
* cell instance $22005 m0 *1 59.925,131.04
X$22005 235 610 236 644 645 cell_1rw
* cell instance $22006 r0 *1 59.925,131.04
X$22006 235 611 236 644 645 cell_1rw
* cell instance $22007 m0 *1 59.925,133.77
X$22007 235 612 236 644 645 cell_1rw
* cell instance $22008 r0 *1 59.925,133.77
X$22008 235 613 236 644 645 cell_1rw
* cell instance $22009 m0 *1 59.925,136.5
X$22009 235 615 236 644 645 cell_1rw
* cell instance $22010 m0 *1 59.925,139.23
X$22010 235 617 236 644 645 cell_1rw
* cell instance $22011 r0 *1 59.925,136.5
X$22011 235 614 236 644 645 cell_1rw
* cell instance $22012 r0 *1 59.925,139.23
X$22012 235 616 236 644 645 cell_1rw
* cell instance $22013 m0 *1 59.925,141.96
X$22013 235 618 236 644 645 cell_1rw
* cell instance $22014 r0 *1 59.925,141.96
X$22014 235 619 236 644 645 cell_1rw
* cell instance $22015 m0 *1 59.925,144.69
X$22015 235 620 236 644 645 cell_1rw
* cell instance $22016 r0 *1 59.925,144.69
X$22016 235 621 236 644 645 cell_1rw
* cell instance $22017 m0 *1 59.925,147.42
X$22017 235 622 236 644 645 cell_1rw
* cell instance $22018 r0 *1 59.925,147.42
X$22018 235 623 236 644 645 cell_1rw
* cell instance $22019 m0 *1 59.925,150.15
X$22019 235 624 236 644 645 cell_1rw
* cell instance $22020 r0 *1 59.925,150.15
X$22020 235 625 236 644 645 cell_1rw
* cell instance $22021 m0 *1 59.925,152.88
X$22021 235 626 236 644 645 cell_1rw
* cell instance $22022 r0 *1 59.925,152.88
X$22022 235 627 236 644 645 cell_1rw
* cell instance $22023 m0 *1 59.925,155.61
X$22023 235 628 236 644 645 cell_1rw
* cell instance $22024 r0 *1 59.925,155.61
X$22024 235 629 236 644 645 cell_1rw
* cell instance $22025 m0 *1 59.925,158.34
X$22025 235 630 236 644 645 cell_1rw
* cell instance $22026 r0 *1 59.925,158.34
X$22026 235 631 236 644 645 cell_1rw
* cell instance $22027 m0 *1 59.925,161.07
X$22027 235 632 236 644 645 cell_1rw
* cell instance $22028 r0 *1 59.925,161.07
X$22028 235 633 236 644 645 cell_1rw
* cell instance $22029 m0 *1 59.925,163.8
X$22029 235 634 236 644 645 cell_1rw
* cell instance $22030 r0 *1 59.925,163.8
X$22030 235 635 236 644 645 cell_1rw
* cell instance $22031 m0 *1 59.925,166.53
X$22031 235 637 236 644 645 cell_1rw
* cell instance $22032 r0 *1 59.925,166.53
X$22032 235 636 236 644 645 cell_1rw
* cell instance $22033 m0 *1 59.925,169.26
X$22033 235 639 236 644 645 cell_1rw
* cell instance $22034 r0 *1 59.925,169.26
X$22034 235 638 236 644 645 cell_1rw
* cell instance $22035 m0 *1 59.925,171.99
X$22035 235 640 236 644 645 cell_1rw
* cell instance $22036 r0 *1 59.925,171.99
X$22036 235 641 236 644 645 cell_1rw
* cell instance $22037 m0 *1 59.925,174.72
X$22037 235 642 236 644 645 cell_1rw
* cell instance $22038 r0 *1 59.925,174.72
X$22038 235 643 236 644 645 cell_1rw
* cell instance $22039 r0 *1 60.63,87.36
X$22039 237 322 238 644 645 cell_1rw
* cell instance $22040 m0 *1 60.63,90.09
X$22040 237 581 238 644 645 cell_1rw
* cell instance $22041 r0 *1 60.63,90.09
X$22041 237 580 238 644 645 cell_1rw
* cell instance $22042 m0 *1 60.63,92.82
X$22042 237 583 238 644 645 cell_1rw
* cell instance $22043 r0 *1 60.63,92.82
X$22043 237 582 238 644 645 cell_1rw
* cell instance $22044 m0 *1 60.63,95.55
X$22044 237 584 238 644 645 cell_1rw
* cell instance $22045 r0 *1 60.63,95.55
X$22045 237 585 238 644 645 cell_1rw
* cell instance $22046 m0 *1 60.63,98.28
X$22046 237 586 238 644 645 cell_1rw
* cell instance $22047 r0 *1 60.63,98.28
X$22047 237 587 238 644 645 cell_1rw
* cell instance $22048 m0 *1 60.63,101.01
X$22048 237 588 238 644 645 cell_1rw
* cell instance $22049 r0 *1 60.63,101.01
X$22049 237 589 238 644 645 cell_1rw
* cell instance $22050 m0 *1 60.63,103.74
X$22050 237 590 238 644 645 cell_1rw
* cell instance $22051 r0 *1 60.63,103.74
X$22051 237 591 238 644 645 cell_1rw
* cell instance $22052 m0 *1 60.63,106.47
X$22052 237 593 238 644 645 cell_1rw
* cell instance $22053 r0 *1 60.63,106.47
X$22053 237 592 238 644 645 cell_1rw
* cell instance $22054 m0 *1 60.63,109.2
X$22054 237 594 238 644 645 cell_1rw
* cell instance $22055 r0 *1 60.63,109.2
X$22055 237 595 238 644 645 cell_1rw
* cell instance $22056 m0 *1 60.63,111.93
X$22056 237 597 238 644 645 cell_1rw
* cell instance $22057 r0 *1 60.63,111.93
X$22057 237 596 238 644 645 cell_1rw
* cell instance $22058 m0 *1 60.63,114.66
X$22058 237 598 238 644 645 cell_1rw
* cell instance $22059 r0 *1 60.63,114.66
X$22059 237 599 238 644 645 cell_1rw
* cell instance $22060 m0 *1 60.63,117.39
X$22060 237 600 238 644 645 cell_1rw
* cell instance $22061 r0 *1 60.63,117.39
X$22061 237 601 238 644 645 cell_1rw
* cell instance $22062 m0 *1 60.63,120.12
X$22062 237 602 238 644 645 cell_1rw
* cell instance $22063 r0 *1 60.63,120.12
X$22063 237 603 238 644 645 cell_1rw
* cell instance $22064 m0 *1 60.63,122.85
X$22064 237 604 238 644 645 cell_1rw
* cell instance $22065 r0 *1 60.63,122.85
X$22065 237 605 238 644 645 cell_1rw
* cell instance $22066 m0 *1 60.63,125.58
X$22066 237 606 238 644 645 cell_1rw
* cell instance $22067 r0 *1 60.63,125.58
X$22067 237 607 238 644 645 cell_1rw
* cell instance $22068 m0 *1 60.63,128.31
X$22068 237 609 238 644 645 cell_1rw
* cell instance $22069 m0 *1 60.63,131.04
X$22069 237 610 238 644 645 cell_1rw
* cell instance $22070 r0 *1 60.63,128.31
X$22070 237 608 238 644 645 cell_1rw
* cell instance $22071 r0 *1 60.63,131.04
X$22071 237 611 238 644 645 cell_1rw
* cell instance $22072 m0 *1 60.63,133.77
X$22072 237 612 238 644 645 cell_1rw
* cell instance $22073 r0 *1 60.63,133.77
X$22073 237 613 238 644 645 cell_1rw
* cell instance $22074 m0 *1 60.63,136.5
X$22074 237 615 238 644 645 cell_1rw
* cell instance $22075 r0 *1 60.63,136.5
X$22075 237 614 238 644 645 cell_1rw
* cell instance $22076 m0 *1 60.63,139.23
X$22076 237 617 238 644 645 cell_1rw
* cell instance $22077 r0 *1 60.63,139.23
X$22077 237 616 238 644 645 cell_1rw
* cell instance $22078 m0 *1 60.63,141.96
X$22078 237 618 238 644 645 cell_1rw
* cell instance $22079 r0 *1 60.63,141.96
X$22079 237 619 238 644 645 cell_1rw
* cell instance $22080 m0 *1 60.63,144.69
X$22080 237 620 238 644 645 cell_1rw
* cell instance $22081 r0 *1 60.63,144.69
X$22081 237 621 238 644 645 cell_1rw
* cell instance $22082 m0 *1 60.63,147.42
X$22082 237 622 238 644 645 cell_1rw
* cell instance $22083 m0 *1 60.63,150.15
X$22083 237 624 238 644 645 cell_1rw
* cell instance $22084 r0 *1 60.63,147.42
X$22084 237 623 238 644 645 cell_1rw
* cell instance $22085 r0 *1 60.63,150.15
X$22085 237 625 238 644 645 cell_1rw
* cell instance $22086 m0 *1 60.63,152.88
X$22086 237 626 238 644 645 cell_1rw
* cell instance $22087 r0 *1 60.63,152.88
X$22087 237 627 238 644 645 cell_1rw
* cell instance $22088 m0 *1 60.63,155.61
X$22088 237 628 238 644 645 cell_1rw
* cell instance $22089 r0 *1 60.63,155.61
X$22089 237 629 238 644 645 cell_1rw
* cell instance $22090 m0 *1 60.63,158.34
X$22090 237 630 238 644 645 cell_1rw
* cell instance $22091 r0 *1 60.63,158.34
X$22091 237 631 238 644 645 cell_1rw
* cell instance $22092 m0 *1 60.63,161.07
X$22092 237 632 238 644 645 cell_1rw
* cell instance $22093 r0 *1 60.63,161.07
X$22093 237 633 238 644 645 cell_1rw
* cell instance $22094 m0 *1 60.63,163.8
X$22094 237 634 238 644 645 cell_1rw
* cell instance $22095 r0 *1 60.63,163.8
X$22095 237 635 238 644 645 cell_1rw
* cell instance $22096 m0 *1 60.63,166.53
X$22096 237 637 238 644 645 cell_1rw
* cell instance $22097 r0 *1 60.63,166.53
X$22097 237 636 238 644 645 cell_1rw
* cell instance $22098 m0 *1 60.63,169.26
X$22098 237 639 238 644 645 cell_1rw
* cell instance $22099 r0 *1 60.63,169.26
X$22099 237 638 238 644 645 cell_1rw
* cell instance $22100 m0 *1 60.63,171.99
X$22100 237 640 238 644 645 cell_1rw
* cell instance $22101 r0 *1 60.63,171.99
X$22101 237 641 238 644 645 cell_1rw
* cell instance $22102 m0 *1 60.63,174.72
X$22102 237 642 238 644 645 cell_1rw
* cell instance $22103 r0 *1 60.63,174.72
X$22103 237 643 238 644 645 cell_1rw
* cell instance $22104 m0 *1 61.335,90.09
X$22104 239 581 240 644 645 cell_1rw
* cell instance $22105 r0 *1 61.335,87.36
X$22105 239 322 240 644 645 cell_1rw
* cell instance $22106 r0 *1 61.335,90.09
X$22106 239 580 240 644 645 cell_1rw
* cell instance $22107 m0 *1 61.335,92.82
X$22107 239 583 240 644 645 cell_1rw
* cell instance $22108 r0 *1 61.335,92.82
X$22108 239 582 240 644 645 cell_1rw
* cell instance $22109 m0 *1 61.335,95.55
X$22109 239 584 240 644 645 cell_1rw
* cell instance $22110 r0 *1 61.335,95.55
X$22110 239 585 240 644 645 cell_1rw
* cell instance $22111 m0 *1 61.335,98.28
X$22111 239 586 240 644 645 cell_1rw
* cell instance $22112 r0 *1 61.335,98.28
X$22112 239 587 240 644 645 cell_1rw
* cell instance $22113 m0 *1 61.335,101.01
X$22113 239 588 240 644 645 cell_1rw
* cell instance $22114 r0 *1 61.335,101.01
X$22114 239 589 240 644 645 cell_1rw
* cell instance $22115 m0 *1 61.335,103.74
X$22115 239 590 240 644 645 cell_1rw
* cell instance $22116 r0 *1 61.335,103.74
X$22116 239 591 240 644 645 cell_1rw
* cell instance $22117 m0 *1 61.335,106.47
X$22117 239 593 240 644 645 cell_1rw
* cell instance $22118 m0 *1 61.335,109.2
X$22118 239 594 240 644 645 cell_1rw
* cell instance $22119 r0 *1 61.335,106.47
X$22119 239 592 240 644 645 cell_1rw
* cell instance $22120 r0 *1 61.335,109.2
X$22120 239 595 240 644 645 cell_1rw
* cell instance $22121 m0 *1 61.335,111.93
X$22121 239 597 240 644 645 cell_1rw
* cell instance $22122 r0 *1 61.335,111.93
X$22122 239 596 240 644 645 cell_1rw
* cell instance $22123 m0 *1 61.335,114.66
X$22123 239 598 240 644 645 cell_1rw
* cell instance $22124 r0 *1 61.335,114.66
X$22124 239 599 240 644 645 cell_1rw
* cell instance $22125 m0 *1 61.335,117.39
X$22125 239 600 240 644 645 cell_1rw
* cell instance $22126 r0 *1 61.335,117.39
X$22126 239 601 240 644 645 cell_1rw
* cell instance $22127 m0 *1 61.335,120.12
X$22127 239 602 240 644 645 cell_1rw
* cell instance $22128 r0 *1 61.335,120.12
X$22128 239 603 240 644 645 cell_1rw
* cell instance $22129 m0 *1 61.335,122.85
X$22129 239 604 240 644 645 cell_1rw
* cell instance $22130 r0 *1 61.335,122.85
X$22130 239 605 240 644 645 cell_1rw
* cell instance $22131 m0 *1 61.335,125.58
X$22131 239 606 240 644 645 cell_1rw
* cell instance $22132 r0 *1 61.335,125.58
X$22132 239 607 240 644 645 cell_1rw
* cell instance $22133 m0 *1 61.335,128.31
X$22133 239 609 240 644 645 cell_1rw
* cell instance $22134 r0 *1 61.335,128.31
X$22134 239 608 240 644 645 cell_1rw
* cell instance $22135 m0 *1 61.335,131.04
X$22135 239 610 240 644 645 cell_1rw
* cell instance $22136 m0 *1 61.335,133.77
X$22136 239 612 240 644 645 cell_1rw
* cell instance $22137 r0 *1 61.335,131.04
X$22137 239 611 240 644 645 cell_1rw
* cell instance $22138 m0 *1 61.335,136.5
X$22138 239 615 240 644 645 cell_1rw
* cell instance $22139 r0 *1 61.335,133.77
X$22139 239 613 240 644 645 cell_1rw
* cell instance $22140 m0 *1 61.335,139.23
X$22140 239 617 240 644 645 cell_1rw
* cell instance $22141 r0 *1 61.335,136.5
X$22141 239 614 240 644 645 cell_1rw
* cell instance $22142 r0 *1 61.335,139.23
X$22142 239 616 240 644 645 cell_1rw
* cell instance $22143 m0 *1 61.335,141.96
X$22143 239 618 240 644 645 cell_1rw
* cell instance $22144 r0 *1 61.335,141.96
X$22144 239 619 240 644 645 cell_1rw
* cell instance $22145 m0 *1 61.335,144.69
X$22145 239 620 240 644 645 cell_1rw
* cell instance $22146 r0 *1 61.335,144.69
X$22146 239 621 240 644 645 cell_1rw
* cell instance $22147 m0 *1 61.335,147.42
X$22147 239 622 240 644 645 cell_1rw
* cell instance $22148 r0 *1 61.335,147.42
X$22148 239 623 240 644 645 cell_1rw
* cell instance $22149 m0 *1 61.335,150.15
X$22149 239 624 240 644 645 cell_1rw
* cell instance $22150 r0 *1 61.335,150.15
X$22150 239 625 240 644 645 cell_1rw
* cell instance $22151 m0 *1 61.335,152.88
X$22151 239 626 240 644 645 cell_1rw
* cell instance $22152 r0 *1 61.335,152.88
X$22152 239 627 240 644 645 cell_1rw
* cell instance $22153 m0 *1 61.335,155.61
X$22153 239 628 240 644 645 cell_1rw
* cell instance $22154 r0 *1 61.335,155.61
X$22154 239 629 240 644 645 cell_1rw
* cell instance $22155 m0 *1 61.335,158.34
X$22155 239 630 240 644 645 cell_1rw
* cell instance $22156 r0 *1 61.335,158.34
X$22156 239 631 240 644 645 cell_1rw
* cell instance $22157 m0 *1 61.335,161.07
X$22157 239 632 240 644 645 cell_1rw
* cell instance $22158 r0 *1 61.335,161.07
X$22158 239 633 240 644 645 cell_1rw
* cell instance $22159 m0 *1 61.335,163.8
X$22159 239 634 240 644 645 cell_1rw
* cell instance $22160 r0 *1 61.335,163.8
X$22160 239 635 240 644 645 cell_1rw
* cell instance $22161 m0 *1 61.335,166.53
X$22161 239 637 240 644 645 cell_1rw
* cell instance $22162 m0 *1 61.335,169.26
X$22162 239 639 240 644 645 cell_1rw
* cell instance $22163 r0 *1 61.335,166.53
X$22163 239 636 240 644 645 cell_1rw
* cell instance $22164 r0 *1 61.335,169.26
X$22164 239 638 240 644 645 cell_1rw
* cell instance $22165 m0 *1 61.335,171.99
X$22165 239 640 240 644 645 cell_1rw
* cell instance $22166 r0 *1 61.335,171.99
X$22166 239 641 240 644 645 cell_1rw
* cell instance $22167 m0 *1 61.335,174.72
X$22167 239 642 240 644 645 cell_1rw
* cell instance $22168 r0 *1 61.335,174.72
X$22168 239 643 240 644 645 cell_1rw
* cell instance $22169 r0 *1 62.04,87.36
X$22169 241 322 242 644 645 cell_1rw
* cell instance $22170 m0 *1 62.04,90.09
X$22170 241 581 242 644 645 cell_1rw
* cell instance $22171 r0 *1 62.04,90.09
X$22171 241 580 242 644 645 cell_1rw
* cell instance $22172 m0 *1 62.04,92.82
X$22172 241 583 242 644 645 cell_1rw
* cell instance $22173 r0 *1 62.04,92.82
X$22173 241 582 242 644 645 cell_1rw
* cell instance $22174 m0 *1 62.04,95.55
X$22174 241 584 242 644 645 cell_1rw
* cell instance $22175 r0 *1 62.04,95.55
X$22175 241 585 242 644 645 cell_1rw
* cell instance $22176 m0 *1 62.04,98.28
X$22176 241 586 242 644 645 cell_1rw
* cell instance $22177 r0 *1 62.04,98.28
X$22177 241 587 242 644 645 cell_1rw
* cell instance $22178 m0 *1 62.04,101.01
X$22178 241 588 242 644 645 cell_1rw
* cell instance $22179 r0 *1 62.04,101.01
X$22179 241 589 242 644 645 cell_1rw
* cell instance $22180 m0 *1 62.04,103.74
X$22180 241 590 242 644 645 cell_1rw
* cell instance $22181 r0 *1 62.04,103.74
X$22181 241 591 242 644 645 cell_1rw
* cell instance $22182 m0 *1 62.04,106.47
X$22182 241 593 242 644 645 cell_1rw
* cell instance $22183 r0 *1 62.04,106.47
X$22183 241 592 242 644 645 cell_1rw
* cell instance $22184 m0 *1 62.04,109.2
X$22184 241 594 242 644 645 cell_1rw
* cell instance $22185 r0 *1 62.04,109.2
X$22185 241 595 242 644 645 cell_1rw
* cell instance $22186 m0 *1 62.04,111.93
X$22186 241 597 242 644 645 cell_1rw
* cell instance $22187 r0 *1 62.04,111.93
X$22187 241 596 242 644 645 cell_1rw
* cell instance $22188 m0 *1 62.04,114.66
X$22188 241 598 242 644 645 cell_1rw
* cell instance $22189 r0 *1 62.04,114.66
X$22189 241 599 242 644 645 cell_1rw
* cell instance $22190 m0 *1 62.04,117.39
X$22190 241 600 242 644 645 cell_1rw
* cell instance $22191 r0 *1 62.04,117.39
X$22191 241 601 242 644 645 cell_1rw
* cell instance $22192 m0 *1 62.04,120.12
X$22192 241 602 242 644 645 cell_1rw
* cell instance $22193 r0 *1 62.04,120.12
X$22193 241 603 242 644 645 cell_1rw
* cell instance $22194 m0 *1 62.04,122.85
X$22194 241 604 242 644 645 cell_1rw
* cell instance $22195 r0 *1 62.04,122.85
X$22195 241 605 242 644 645 cell_1rw
* cell instance $22196 m0 *1 62.04,125.58
X$22196 241 606 242 644 645 cell_1rw
* cell instance $22197 r0 *1 62.04,125.58
X$22197 241 607 242 644 645 cell_1rw
* cell instance $22198 m0 *1 62.04,128.31
X$22198 241 609 242 644 645 cell_1rw
* cell instance $22199 r0 *1 62.04,128.31
X$22199 241 608 242 644 645 cell_1rw
* cell instance $22200 m0 *1 62.04,131.04
X$22200 241 610 242 644 645 cell_1rw
* cell instance $22201 r0 *1 62.04,131.04
X$22201 241 611 242 644 645 cell_1rw
* cell instance $22202 m0 *1 62.04,133.77
X$22202 241 612 242 644 645 cell_1rw
* cell instance $22203 r0 *1 62.04,133.77
X$22203 241 613 242 644 645 cell_1rw
* cell instance $22204 m0 *1 62.04,136.5
X$22204 241 615 242 644 645 cell_1rw
* cell instance $22205 r0 *1 62.04,136.5
X$22205 241 614 242 644 645 cell_1rw
* cell instance $22206 m0 *1 62.04,139.23
X$22206 241 617 242 644 645 cell_1rw
* cell instance $22207 m0 *1 62.04,141.96
X$22207 241 618 242 644 645 cell_1rw
* cell instance $22208 r0 *1 62.04,139.23
X$22208 241 616 242 644 645 cell_1rw
* cell instance $22209 r0 *1 62.04,141.96
X$22209 241 619 242 644 645 cell_1rw
* cell instance $22210 m0 *1 62.04,144.69
X$22210 241 620 242 644 645 cell_1rw
* cell instance $22211 r0 *1 62.04,144.69
X$22211 241 621 242 644 645 cell_1rw
* cell instance $22212 m0 *1 62.04,147.42
X$22212 241 622 242 644 645 cell_1rw
* cell instance $22213 r0 *1 62.04,147.42
X$22213 241 623 242 644 645 cell_1rw
* cell instance $22214 m0 *1 62.04,150.15
X$22214 241 624 242 644 645 cell_1rw
* cell instance $22215 r0 *1 62.04,150.15
X$22215 241 625 242 644 645 cell_1rw
* cell instance $22216 m0 *1 62.04,152.88
X$22216 241 626 242 644 645 cell_1rw
* cell instance $22217 r0 *1 62.04,152.88
X$22217 241 627 242 644 645 cell_1rw
* cell instance $22218 m0 *1 62.04,155.61
X$22218 241 628 242 644 645 cell_1rw
* cell instance $22219 r0 *1 62.04,155.61
X$22219 241 629 242 644 645 cell_1rw
* cell instance $22220 m0 *1 62.04,158.34
X$22220 241 630 242 644 645 cell_1rw
* cell instance $22221 m0 *1 62.04,161.07
X$22221 241 632 242 644 645 cell_1rw
* cell instance $22222 r0 *1 62.04,158.34
X$22222 241 631 242 644 645 cell_1rw
* cell instance $22223 r0 *1 62.04,161.07
X$22223 241 633 242 644 645 cell_1rw
* cell instance $22224 m0 *1 62.04,163.8
X$22224 241 634 242 644 645 cell_1rw
* cell instance $22225 r0 *1 62.04,163.8
X$22225 241 635 242 644 645 cell_1rw
* cell instance $22226 m0 *1 62.04,166.53
X$22226 241 637 242 644 645 cell_1rw
* cell instance $22227 r0 *1 62.04,166.53
X$22227 241 636 242 644 645 cell_1rw
* cell instance $22228 m0 *1 62.04,169.26
X$22228 241 639 242 644 645 cell_1rw
* cell instance $22229 r0 *1 62.04,169.26
X$22229 241 638 242 644 645 cell_1rw
* cell instance $22230 m0 *1 62.04,171.99
X$22230 241 640 242 644 645 cell_1rw
* cell instance $22231 r0 *1 62.04,171.99
X$22231 241 641 242 644 645 cell_1rw
* cell instance $22232 m0 *1 62.04,174.72
X$22232 241 642 242 644 645 cell_1rw
* cell instance $22233 r0 *1 62.04,174.72
X$22233 241 643 242 644 645 cell_1rw
* cell instance $22234 r0 *1 62.745,87.36
X$22234 243 322 244 644 645 cell_1rw
* cell instance $22235 m0 *1 62.745,90.09
X$22235 243 581 244 644 645 cell_1rw
* cell instance $22236 r0 *1 62.745,90.09
X$22236 243 580 244 644 645 cell_1rw
* cell instance $22237 m0 *1 62.745,92.82
X$22237 243 583 244 644 645 cell_1rw
* cell instance $22238 m0 *1 62.745,95.55
X$22238 243 584 244 644 645 cell_1rw
* cell instance $22239 r0 *1 62.745,92.82
X$22239 243 582 244 644 645 cell_1rw
* cell instance $22240 r0 *1 62.745,95.55
X$22240 243 585 244 644 645 cell_1rw
* cell instance $22241 m0 *1 62.745,98.28
X$22241 243 586 244 644 645 cell_1rw
* cell instance $22242 r0 *1 62.745,98.28
X$22242 243 587 244 644 645 cell_1rw
* cell instance $22243 m0 *1 62.745,101.01
X$22243 243 588 244 644 645 cell_1rw
* cell instance $22244 m0 *1 62.745,103.74
X$22244 243 590 244 644 645 cell_1rw
* cell instance $22245 r0 *1 62.745,101.01
X$22245 243 589 244 644 645 cell_1rw
* cell instance $22246 r0 *1 62.745,103.74
X$22246 243 591 244 644 645 cell_1rw
* cell instance $22247 m0 *1 62.745,106.47
X$22247 243 593 244 644 645 cell_1rw
* cell instance $22248 r0 *1 62.745,106.47
X$22248 243 592 244 644 645 cell_1rw
* cell instance $22249 m0 *1 62.745,109.2
X$22249 243 594 244 644 645 cell_1rw
* cell instance $22250 r0 *1 62.745,109.2
X$22250 243 595 244 644 645 cell_1rw
* cell instance $22251 m0 *1 62.745,111.93
X$22251 243 597 244 644 645 cell_1rw
* cell instance $22252 r0 *1 62.745,111.93
X$22252 243 596 244 644 645 cell_1rw
* cell instance $22253 m0 *1 62.745,114.66
X$22253 243 598 244 644 645 cell_1rw
* cell instance $22254 r0 *1 62.745,114.66
X$22254 243 599 244 644 645 cell_1rw
* cell instance $22255 m0 *1 62.745,117.39
X$22255 243 600 244 644 645 cell_1rw
* cell instance $22256 r0 *1 62.745,117.39
X$22256 243 601 244 644 645 cell_1rw
* cell instance $22257 m0 *1 62.745,120.12
X$22257 243 602 244 644 645 cell_1rw
* cell instance $22258 m0 *1 62.745,122.85
X$22258 243 604 244 644 645 cell_1rw
* cell instance $22259 r0 *1 62.745,120.12
X$22259 243 603 244 644 645 cell_1rw
* cell instance $22260 r0 *1 62.745,122.85
X$22260 243 605 244 644 645 cell_1rw
* cell instance $22261 m0 *1 62.745,125.58
X$22261 243 606 244 644 645 cell_1rw
* cell instance $22262 r0 *1 62.745,125.58
X$22262 243 607 244 644 645 cell_1rw
* cell instance $22263 m0 *1 62.745,128.31
X$22263 243 609 244 644 645 cell_1rw
* cell instance $22264 r0 *1 62.745,128.31
X$22264 243 608 244 644 645 cell_1rw
* cell instance $22265 m0 *1 62.745,131.04
X$22265 243 610 244 644 645 cell_1rw
* cell instance $22266 r0 *1 62.745,131.04
X$22266 243 611 244 644 645 cell_1rw
* cell instance $22267 m0 *1 62.745,133.77
X$22267 243 612 244 644 645 cell_1rw
* cell instance $22268 r0 *1 62.745,133.77
X$22268 243 613 244 644 645 cell_1rw
* cell instance $22269 m0 *1 62.745,136.5
X$22269 243 615 244 644 645 cell_1rw
* cell instance $22270 r0 *1 62.745,136.5
X$22270 243 614 244 644 645 cell_1rw
* cell instance $22271 m0 *1 62.745,139.23
X$22271 243 617 244 644 645 cell_1rw
* cell instance $22272 r0 *1 62.745,139.23
X$22272 243 616 244 644 645 cell_1rw
* cell instance $22273 m0 *1 62.745,141.96
X$22273 243 618 244 644 645 cell_1rw
* cell instance $22274 r0 *1 62.745,141.96
X$22274 243 619 244 644 645 cell_1rw
* cell instance $22275 m0 *1 62.745,144.69
X$22275 243 620 244 644 645 cell_1rw
* cell instance $22276 m0 *1 62.745,147.42
X$22276 243 622 244 644 645 cell_1rw
* cell instance $22277 r0 *1 62.745,144.69
X$22277 243 621 244 644 645 cell_1rw
* cell instance $22278 m0 *1 62.745,150.15
X$22278 243 624 244 644 645 cell_1rw
* cell instance $22279 r0 *1 62.745,147.42
X$22279 243 623 244 644 645 cell_1rw
* cell instance $22280 r0 *1 62.745,150.15
X$22280 243 625 244 644 645 cell_1rw
* cell instance $22281 m0 *1 62.745,152.88
X$22281 243 626 244 644 645 cell_1rw
* cell instance $22282 r0 *1 62.745,152.88
X$22282 243 627 244 644 645 cell_1rw
* cell instance $22283 m0 *1 62.745,155.61
X$22283 243 628 244 644 645 cell_1rw
* cell instance $22284 r0 *1 62.745,155.61
X$22284 243 629 244 644 645 cell_1rw
* cell instance $22285 m0 *1 62.745,158.34
X$22285 243 630 244 644 645 cell_1rw
* cell instance $22286 r0 *1 62.745,158.34
X$22286 243 631 244 644 645 cell_1rw
* cell instance $22287 m0 *1 62.745,161.07
X$22287 243 632 244 644 645 cell_1rw
* cell instance $22288 m0 *1 62.745,163.8
X$22288 243 634 244 644 645 cell_1rw
* cell instance $22289 r0 *1 62.745,161.07
X$22289 243 633 244 644 645 cell_1rw
* cell instance $22290 r0 *1 62.745,163.8
X$22290 243 635 244 644 645 cell_1rw
* cell instance $22291 m0 *1 62.745,166.53
X$22291 243 637 244 644 645 cell_1rw
* cell instance $22292 r0 *1 62.745,166.53
X$22292 243 636 244 644 645 cell_1rw
* cell instance $22293 m0 *1 62.745,169.26
X$22293 243 639 244 644 645 cell_1rw
* cell instance $22294 r0 *1 62.745,169.26
X$22294 243 638 244 644 645 cell_1rw
* cell instance $22295 m0 *1 62.745,171.99
X$22295 243 640 244 644 645 cell_1rw
* cell instance $22296 m0 *1 62.745,174.72
X$22296 243 642 244 644 645 cell_1rw
* cell instance $22297 r0 *1 62.745,171.99
X$22297 243 641 244 644 645 cell_1rw
* cell instance $22298 r0 *1 62.745,174.72
X$22298 243 643 244 644 645 cell_1rw
* cell instance $22299 r0 *1 63.45,87.36
X$22299 245 322 246 644 645 cell_1rw
* cell instance $22300 m0 *1 63.45,90.09
X$22300 245 581 246 644 645 cell_1rw
* cell instance $22301 r0 *1 63.45,90.09
X$22301 245 580 246 644 645 cell_1rw
* cell instance $22302 m0 *1 63.45,92.82
X$22302 245 583 246 644 645 cell_1rw
* cell instance $22303 m0 *1 63.45,95.55
X$22303 245 584 246 644 645 cell_1rw
* cell instance $22304 r0 *1 63.45,92.82
X$22304 245 582 246 644 645 cell_1rw
* cell instance $22305 r0 *1 63.45,95.55
X$22305 245 585 246 644 645 cell_1rw
* cell instance $22306 m0 *1 63.45,98.28
X$22306 245 586 246 644 645 cell_1rw
* cell instance $22307 r0 *1 63.45,98.28
X$22307 245 587 246 644 645 cell_1rw
* cell instance $22308 m0 *1 63.45,101.01
X$22308 245 588 246 644 645 cell_1rw
* cell instance $22309 r0 *1 63.45,101.01
X$22309 245 589 246 644 645 cell_1rw
* cell instance $22310 m0 *1 63.45,103.74
X$22310 245 590 246 644 645 cell_1rw
* cell instance $22311 m0 *1 63.45,106.47
X$22311 245 593 246 644 645 cell_1rw
* cell instance $22312 r0 *1 63.45,103.74
X$22312 245 591 246 644 645 cell_1rw
* cell instance $22313 r0 *1 63.45,106.47
X$22313 245 592 246 644 645 cell_1rw
* cell instance $22314 m0 *1 63.45,109.2
X$22314 245 594 246 644 645 cell_1rw
* cell instance $22315 r0 *1 63.45,109.2
X$22315 245 595 246 644 645 cell_1rw
* cell instance $22316 m0 *1 63.45,111.93
X$22316 245 597 246 644 645 cell_1rw
* cell instance $22317 r0 *1 63.45,111.93
X$22317 245 596 246 644 645 cell_1rw
* cell instance $22318 m0 *1 63.45,114.66
X$22318 245 598 246 644 645 cell_1rw
* cell instance $22319 m0 *1 63.45,117.39
X$22319 245 600 246 644 645 cell_1rw
* cell instance $22320 r0 *1 63.45,114.66
X$22320 245 599 246 644 645 cell_1rw
* cell instance $22321 m0 *1 63.45,120.12
X$22321 245 602 246 644 645 cell_1rw
* cell instance $22322 r0 *1 63.45,117.39
X$22322 245 601 246 644 645 cell_1rw
* cell instance $22323 r0 *1 63.45,120.12
X$22323 245 603 246 644 645 cell_1rw
* cell instance $22324 m0 *1 63.45,122.85
X$22324 245 604 246 644 645 cell_1rw
* cell instance $22325 r0 *1 63.45,122.85
X$22325 245 605 246 644 645 cell_1rw
* cell instance $22326 m0 *1 63.45,125.58
X$22326 245 606 246 644 645 cell_1rw
* cell instance $22327 r0 *1 63.45,125.58
X$22327 245 607 246 644 645 cell_1rw
* cell instance $22328 m0 *1 63.45,128.31
X$22328 245 609 246 644 645 cell_1rw
* cell instance $22329 r0 *1 63.45,128.31
X$22329 245 608 246 644 645 cell_1rw
* cell instance $22330 m0 *1 63.45,131.04
X$22330 245 610 246 644 645 cell_1rw
* cell instance $22331 r0 *1 63.45,131.04
X$22331 245 611 246 644 645 cell_1rw
* cell instance $22332 m0 *1 63.45,133.77
X$22332 245 612 246 644 645 cell_1rw
* cell instance $22333 m0 *1 63.45,136.5
X$22333 245 615 246 644 645 cell_1rw
* cell instance $22334 r0 *1 63.45,133.77
X$22334 245 613 246 644 645 cell_1rw
* cell instance $22335 r0 *1 63.45,136.5
X$22335 245 614 246 644 645 cell_1rw
* cell instance $22336 m0 *1 63.45,139.23
X$22336 245 617 246 644 645 cell_1rw
* cell instance $22337 r0 *1 63.45,139.23
X$22337 245 616 246 644 645 cell_1rw
* cell instance $22338 m0 *1 63.45,141.96
X$22338 245 618 246 644 645 cell_1rw
* cell instance $22339 r0 *1 63.45,141.96
X$22339 245 619 246 644 645 cell_1rw
* cell instance $22340 m0 *1 63.45,144.69
X$22340 245 620 246 644 645 cell_1rw
* cell instance $22341 r0 *1 63.45,144.69
X$22341 245 621 246 644 645 cell_1rw
* cell instance $22342 m0 *1 63.45,147.42
X$22342 245 622 246 644 645 cell_1rw
* cell instance $22343 m0 *1 63.45,150.15
X$22343 245 624 246 644 645 cell_1rw
* cell instance $22344 r0 *1 63.45,147.42
X$22344 245 623 246 644 645 cell_1rw
* cell instance $22345 r0 *1 63.45,150.15
X$22345 245 625 246 644 645 cell_1rw
* cell instance $22346 m0 *1 63.45,152.88
X$22346 245 626 246 644 645 cell_1rw
* cell instance $22347 r0 *1 63.45,152.88
X$22347 245 627 246 644 645 cell_1rw
* cell instance $22348 m0 *1 63.45,155.61
X$22348 245 628 246 644 645 cell_1rw
* cell instance $22349 r0 *1 63.45,155.61
X$22349 245 629 246 644 645 cell_1rw
* cell instance $22350 m0 *1 63.45,158.34
X$22350 245 630 246 644 645 cell_1rw
* cell instance $22351 m0 *1 63.45,161.07
X$22351 245 632 246 644 645 cell_1rw
* cell instance $22352 r0 *1 63.45,158.34
X$22352 245 631 246 644 645 cell_1rw
* cell instance $22353 m0 *1 63.45,163.8
X$22353 245 634 246 644 645 cell_1rw
* cell instance $22354 r0 *1 63.45,161.07
X$22354 245 633 246 644 645 cell_1rw
* cell instance $22355 m0 *1 63.45,166.53
X$22355 245 637 246 644 645 cell_1rw
* cell instance $22356 r0 *1 63.45,163.8
X$22356 245 635 246 644 645 cell_1rw
* cell instance $22357 r0 *1 63.45,166.53
X$22357 245 636 246 644 645 cell_1rw
* cell instance $22358 m0 *1 63.45,169.26
X$22358 245 639 246 644 645 cell_1rw
* cell instance $22359 m0 *1 63.45,171.99
X$22359 245 640 246 644 645 cell_1rw
* cell instance $22360 r0 *1 63.45,169.26
X$22360 245 638 246 644 645 cell_1rw
* cell instance $22361 r0 *1 63.45,171.99
X$22361 245 641 246 644 645 cell_1rw
* cell instance $22362 m0 *1 63.45,174.72
X$22362 245 642 246 644 645 cell_1rw
* cell instance $22363 r0 *1 63.45,174.72
X$22363 245 643 246 644 645 cell_1rw
* cell instance $22364 r0 *1 64.155,87.36
X$22364 247 322 248 644 645 cell_1rw
* cell instance $22365 m0 *1 64.155,90.09
X$22365 247 581 248 644 645 cell_1rw
* cell instance $22366 r0 *1 64.155,90.09
X$22366 247 580 248 644 645 cell_1rw
* cell instance $22367 m0 *1 64.155,92.82
X$22367 247 583 248 644 645 cell_1rw
* cell instance $22368 r0 *1 64.155,92.82
X$22368 247 582 248 644 645 cell_1rw
* cell instance $22369 m0 *1 64.155,95.55
X$22369 247 584 248 644 645 cell_1rw
* cell instance $22370 r0 *1 64.155,95.55
X$22370 247 585 248 644 645 cell_1rw
* cell instance $22371 m0 *1 64.155,98.28
X$22371 247 586 248 644 645 cell_1rw
* cell instance $22372 r0 *1 64.155,98.28
X$22372 247 587 248 644 645 cell_1rw
* cell instance $22373 m0 *1 64.155,101.01
X$22373 247 588 248 644 645 cell_1rw
* cell instance $22374 r0 *1 64.155,101.01
X$22374 247 589 248 644 645 cell_1rw
* cell instance $22375 m0 *1 64.155,103.74
X$22375 247 590 248 644 645 cell_1rw
* cell instance $22376 m0 *1 64.155,106.47
X$22376 247 593 248 644 645 cell_1rw
* cell instance $22377 r0 *1 64.155,103.74
X$22377 247 591 248 644 645 cell_1rw
* cell instance $22378 r0 *1 64.155,106.47
X$22378 247 592 248 644 645 cell_1rw
* cell instance $22379 m0 *1 64.155,109.2
X$22379 247 594 248 644 645 cell_1rw
* cell instance $22380 r0 *1 64.155,109.2
X$22380 247 595 248 644 645 cell_1rw
* cell instance $22381 m0 *1 64.155,111.93
X$22381 247 597 248 644 645 cell_1rw
* cell instance $22382 r0 *1 64.155,111.93
X$22382 247 596 248 644 645 cell_1rw
* cell instance $22383 m0 *1 64.155,114.66
X$22383 247 598 248 644 645 cell_1rw
* cell instance $22384 r0 *1 64.155,114.66
X$22384 247 599 248 644 645 cell_1rw
* cell instance $22385 m0 *1 64.155,117.39
X$22385 247 600 248 644 645 cell_1rw
* cell instance $22386 r0 *1 64.155,117.39
X$22386 247 601 248 644 645 cell_1rw
* cell instance $22387 m0 *1 64.155,120.12
X$22387 247 602 248 644 645 cell_1rw
* cell instance $22388 r0 *1 64.155,120.12
X$22388 247 603 248 644 645 cell_1rw
* cell instance $22389 m0 *1 64.155,122.85
X$22389 247 604 248 644 645 cell_1rw
* cell instance $22390 r0 *1 64.155,122.85
X$22390 247 605 248 644 645 cell_1rw
* cell instance $22391 m0 *1 64.155,125.58
X$22391 247 606 248 644 645 cell_1rw
* cell instance $22392 r0 *1 64.155,125.58
X$22392 247 607 248 644 645 cell_1rw
* cell instance $22393 m0 *1 64.155,128.31
X$22393 247 609 248 644 645 cell_1rw
* cell instance $22394 r0 *1 64.155,128.31
X$22394 247 608 248 644 645 cell_1rw
* cell instance $22395 m0 *1 64.155,131.04
X$22395 247 610 248 644 645 cell_1rw
* cell instance $22396 r0 *1 64.155,131.04
X$22396 247 611 248 644 645 cell_1rw
* cell instance $22397 m0 *1 64.155,133.77
X$22397 247 612 248 644 645 cell_1rw
* cell instance $22398 r0 *1 64.155,133.77
X$22398 247 613 248 644 645 cell_1rw
* cell instance $22399 m0 *1 64.155,136.5
X$22399 247 615 248 644 645 cell_1rw
* cell instance $22400 r0 *1 64.155,136.5
X$22400 247 614 248 644 645 cell_1rw
* cell instance $22401 m0 *1 64.155,139.23
X$22401 247 617 248 644 645 cell_1rw
* cell instance $22402 m0 *1 64.155,141.96
X$22402 247 618 248 644 645 cell_1rw
* cell instance $22403 r0 *1 64.155,139.23
X$22403 247 616 248 644 645 cell_1rw
* cell instance $22404 r0 *1 64.155,141.96
X$22404 247 619 248 644 645 cell_1rw
* cell instance $22405 m0 *1 64.155,144.69
X$22405 247 620 248 644 645 cell_1rw
* cell instance $22406 r0 *1 64.155,144.69
X$22406 247 621 248 644 645 cell_1rw
* cell instance $22407 m0 *1 64.155,147.42
X$22407 247 622 248 644 645 cell_1rw
* cell instance $22408 r0 *1 64.155,147.42
X$22408 247 623 248 644 645 cell_1rw
* cell instance $22409 m0 *1 64.155,150.15
X$22409 247 624 248 644 645 cell_1rw
* cell instance $22410 r0 *1 64.155,150.15
X$22410 247 625 248 644 645 cell_1rw
* cell instance $22411 m0 *1 64.155,152.88
X$22411 247 626 248 644 645 cell_1rw
* cell instance $22412 r0 *1 64.155,152.88
X$22412 247 627 248 644 645 cell_1rw
* cell instance $22413 m0 *1 64.155,155.61
X$22413 247 628 248 644 645 cell_1rw
* cell instance $22414 r0 *1 64.155,155.61
X$22414 247 629 248 644 645 cell_1rw
* cell instance $22415 m0 *1 64.155,158.34
X$22415 247 630 248 644 645 cell_1rw
* cell instance $22416 r0 *1 64.155,158.34
X$22416 247 631 248 644 645 cell_1rw
* cell instance $22417 m0 *1 64.155,161.07
X$22417 247 632 248 644 645 cell_1rw
* cell instance $22418 r0 *1 64.155,161.07
X$22418 247 633 248 644 645 cell_1rw
* cell instance $22419 m0 *1 64.155,163.8
X$22419 247 634 248 644 645 cell_1rw
* cell instance $22420 r0 *1 64.155,163.8
X$22420 247 635 248 644 645 cell_1rw
* cell instance $22421 m0 *1 64.155,166.53
X$22421 247 637 248 644 645 cell_1rw
* cell instance $22422 r0 *1 64.155,166.53
X$22422 247 636 248 644 645 cell_1rw
* cell instance $22423 m0 *1 64.155,169.26
X$22423 247 639 248 644 645 cell_1rw
* cell instance $22424 m0 *1 64.155,171.99
X$22424 247 640 248 644 645 cell_1rw
* cell instance $22425 r0 *1 64.155,169.26
X$22425 247 638 248 644 645 cell_1rw
* cell instance $22426 r0 *1 64.155,171.99
X$22426 247 641 248 644 645 cell_1rw
* cell instance $22427 m0 *1 64.155,174.72
X$22427 247 642 248 644 645 cell_1rw
* cell instance $22428 r0 *1 64.155,174.72
X$22428 247 643 248 644 645 cell_1rw
* cell instance $22429 r0 *1 64.86,87.36
X$22429 249 322 250 644 645 cell_1rw
* cell instance $22430 m0 *1 64.86,90.09
X$22430 249 581 250 644 645 cell_1rw
* cell instance $22431 r0 *1 64.86,90.09
X$22431 249 580 250 644 645 cell_1rw
* cell instance $22432 m0 *1 64.86,92.82
X$22432 249 583 250 644 645 cell_1rw
* cell instance $22433 r0 *1 64.86,92.82
X$22433 249 582 250 644 645 cell_1rw
* cell instance $22434 m0 *1 64.86,95.55
X$22434 249 584 250 644 645 cell_1rw
* cell instance $22435 r0 *1 64.86,95.55
X$22435 249 585 250 644 645 cell_1rw
* cell instance $22436 m0 *1 64.86,98.28
X$22436 249 586 250 644 645 cell_1rw
* cell instance $22437 r0 *1 64.86,98.28
X$22437 249 587 250 644 645 cell_1rw
* cell instance $22438 m0 *1 64.86,101.01
X$22438 249 588 250 644 645 cell_1rw
* cell instance $22439 r0 *1 64.86,101.01
X$22439 249 589 250 644 645 cell_1rw
* cell instance $22440 m0 *1 64.86,103.74
X$22440 249 590 250 644 645 cell_1rw
* cell instance $22441 r0 *1 64.86,103.74
X$22441 249 591 250 644 645 cell_1rw
* cell instance $22442 m0 *1 64.86,106.47
X$22442 249 593 250 644 645 cell_1rw
* cell instance $22443 r0 *1 64.86,106.47
X$22443 249 592 250 644 645 cell_1rw
* cell instance $22444 m0 *1 64.86,109.2
X$22444 249 594 250 644 645 cell_1rw
* cell instance $22445 r0 *1 64.86,109.2
X$22445 249 595 250 644 645 cell_1rw
* cell instance $22446 m0 *1 64.86,111.93
X$22446 249 597 250 644 645 cell_1rw
* cell instance $22447 r0 *1 64.86,111.93
X$22447 249 596 250 644 645 cell_1rw
* cell instance $22448 m0 *1 64.86,114.66
X$22448 249 598 250 644 645 cell_1rw
* cell instance $22449 r0 *1 64.86,114.66
X$22449 249 599 250 644 645 cell_1rw
* cell instance $22450 m0 *1 64.86,117.39
X$22450 249 600 250 644 645 cell_1rw
* cell instance $22451 r0 *1 64.86,117.39
X$22451 249 601 250 644 645 cell_1rw
* cell instance $22452 m0 *1 64.86,120.12
X$22452 249 602 250 644 645 cell_1rw
* cell instance $22453 r0 *1 64.86,120.12
X$22453 249 603 250 644 645 cell_1rw
* cell instance $22454 m0 *1 64.86,122.85
X$22454 249 604 250 644 645 cell_1rw
* cell instance $22455 r0 *1 64.86,122.85
X$22455 249 605 250 644 645 cell_1rw
* cell instance $22456 m0 *1 64.86,125.58
X$22456 249 606 250 644 645 cell_1rw
* cell instance $22457 r0 *1 64.86,125.58
X$22457 249 607 250 644 645 cell_1rw
* cell instance $22458 m0 *1 64.86,128.31
X$22458 249 609 250 644 645 cell_1rw
* cell instance $22459 r0 *1 64.86,128.31
X$22459 249 608 250 644 645 cell_1rw
* cell instance $22460 m0 *1 64.86,131.04
X$22460 249 610 250 644 645 cell_1rw
* cell instance $22461 r0 *1 64.86,131.04
X$22461 249 611 250 644 645 cell_1rw
* cell instance $22462 m0 *1 64.86,133.77
X$22462 249 612 250 644 645 cell_1rw
* cell instance $22463 r0 *1 64.86,133.77
X$22463 249 613 250 644 645 cell_1rw
* cell instance $22464 m0 *1 64.86,136.5
X$22464 249 615 250 644 645 cell_1rw
* cell instance $22465 r0 *1 64.86,136.5
X$22465 249 614 250 644 645 cell_1rw
* cell instance $22466 m0 *1 64.86,139.23
X$22466 249 617 250 644 645 cell_1rw
* cell instance $22467 m0 *1 64.86,141.96
X$22467 249 618 250 644 645 cell_1rw
* cell instance $22468 r0 *1 64.86,139.23
X$22468 249 616 250 644 645 cell_1rw
* cell instance $22469 r0 *1 64.86,141.96
X$22469 249 619 250 644 645 cell_1rw
* cell instance $22470 m0 *1 64.86,144.69
X$22470 249 620 250 644 645 cell_1rw
* cell instance $22471 m0 *1 64.86,147.42
X$22471 249 622 250 644 645 cell_1rw
* cell instance $22472 r0 *1 64.86,144.69
X$22472 249 621 250 644 645 cell_1rw
* cell instance $22473 r0 *1 64.86,147.42
X$22473 249 623 250 644 645 cell_1rw
* cell instance $22474 m0 *1 64.86,150.15
X$22474 249 624 250 644 645 cell_1rw
* cell instance $22475 m0 *1 64.86,152.88
X$22475 249 626 250 644 645 cell_1rw
* cell instance $22476 r0 *1 64.86,150.15
X$22476 249 625 250 644 645 cell_1rw
* cell instance $22477 r0 *1 64.86,152.88
X$22477 249 627 250 644 645 cell_1rw
* cell instance $22478 m0 *1 64.86,155.61
X$22478 249 628 250 644 645 cell_1rw
* cell instance $22479 r0 *1 64.86,155.61
X$22479 249 629 250 644 645 cell_1rw
* cell instance $22480 m0 *1 64.86,158.34
X$22480 249 630 250 644 645 cell_1rw
* cell instance $22481 m0 *1 64.86,161.07
X$22481 249 632 250 644 645 cell_1rw
* cell instance $22482 r0 *1 64.86,158.34
X$22482 249 631 250 644 645 cell_1rw
* cell instance $22483 r0 *1 64.86,161.07
X$22483 249 633 250 644 645 cell_1rw
* cell instance $22484 m0 *1 64.86,163.8
X$22484 249 634 250 644 645 cell_1rw
* cell instance $22485 r0 *1 64.86,163.8
X$22485 249 635 250 644 645 cell_1rw
* cell instance $22486 m0 *1 64.86,166.53
X$22486 249 637 250 644 645 cell_1rw
* cell instance $22487 r0 *1 64.86,166.53
X$22487 249 636 250 644 645 cell_1rw
* cell instance $22488 m0 *1 64.86,169.26
X$22488 249 639 250 644 645 cell_1rw
* cell instance $22489 r0 *1 64.86,169.26
X$22489 249 638 250 644 645 cell_1rw
* cell instance $22490 m0 *1 64.86,171.99
X$22490 249 640 250 644 645 cell_1rw
* cell instance $22491 r0 *1 64.86,171.99
X$22491 249 641 250 644 645 cell_1rw
* cell instance $22492 m0 *1 64.86,174.72
X$22492 249 642 250 644 645 cell_1rw
* cell instance $22493 r0 *1 64.86,174.72
X$22493 249 643 250 644 645 cell_1rw
* cell instance $22494 r0 *1 65.565,87.36
X$22494 251 322 252 644 645 cell_1rw
* cell instance $22495 m0 *1 65.565,90.09
X$22495 251 581 252 644 645 cell_1rw
* cell instance $22496 m0 *1 65.565,92.82
X$22496 251 583 252 644 645 cell_1rw
* cell instance $22497 r0 *1 65.565,90.09
X$22497 251 580 252 644 645 cell_1rw
* cell instance $22498 r0 *1 65.565,92.82
X$22498 251 582 252 644 645 cell_1rw
* cell instance $22499 m0 *1 65.565,95.55
X$22499 251 584 252 644 645 cell_1rw
* cell instance $22500 r0 *1 65.565,95.55
X$22500 251 585 252 644 645 cell_1rw
* cell instance $22501 m0 *1 65.565,98.28
X$22501 251 586 252 644 645 cell_1rw
* cell instance $22502 r0 *1 65.565,98.28
X$22502 251 587 252 644 645 cell_1rw
* cell instance $22503 m0 *1 65.565,101.01
X$22503 251 588 252 644 645 cell_1rw
* cell instance $22504 r0 *1 65.565,101.01
X$22504 251 589 252 644 645 cell_1rw
* cell instance $22505 m0 *1 65.565,103.74
X$22505 251 590 252 644 645 cell_1rw
* cell instance $22506 r0 *1 65.565,103.74
X$22506 251 591 252 644 645 cell_1rw
* cell instance $22507 m0 *1 65.565,106.47
X$22507 251 593 252 644 645 cell_1rw
* cell instance $22508 r0 *1 65.565,106.47
X$22508 251 592 252 644 645 cell_1rw
* cell instance $22509 m0 *1 65.565,109.2
X$22509 251 594 252 644 645 cell_1rw
* cell instance $22510 r0 *1 65.565,109.2
X$22510 251 595 252 644 645 cell_1rw
* cell instance $22511 m0 *1 65.565,111.93
X$22511 251 597 252 644 645 cell_1rw
* cell instance $22512 r0 *1 65.565,111.93
X$22512 251 596 252 644 645 cell_1rw
* cell instance $22513 m0 *1 65.565,114.66
X$22513 251 598 252 644 645 cell_1rw
* cell instance $22514 m0 *1 65.565,117.39
X$22514 251 600 252 644 645 cell_1rw
* cell instance $22515 r0 *1 65.565,114.66
X$22515 251 599 252 644 645 cell_1rw
* cell instance $22516 r0 *1 65.565,117.39
X$22516 251 601 252 644 645 cell_1rw
* cell instance $22517 m0 *1 65.565,120.12
X$22517 251 602 252 644 645 cell_1rw
* cell instance $22518 r0 *1 65.565,120.12
X$22518 251 603 252 644 645 cell_1rw
* cell instance $22519 m0 *1 65.565,122.85
X$22519 251 604 252 644 645 cell_1rw
* cell instance $22520 r0 *1 65.565,122.85
X$22520 251 605 252 644 645 cell_1rw
* cell instance $22521 m0 *1 65.565,125.58
X$22521 251 606 252 644 645 cell_1rw
* cell instance $22522 r0 *1 65.565,125.58
X$22522 251 607 252 644 645 cell_1rw
* cell instance $22523 m0 *1 65.565,128.31
X$22523 251 609 252 644 645 cell_1rw
* cell instance $22524 r0 *1 65.565,128.31
X$22524 251 608 252 644 645 cell_1rw
* cell instance $22525 m0 *1 65.565,131.04
X$22525 251 610 252 644 645 cell_1rw
* cell instance $22526 r0 *1 65.565,131.04
X$22526 251 611 252 644 645 cell_1rw
* cell instance $22527 m0 *1 65.565,133.77
X$22527 251 612 252 644 645 cell_1rw
* cell instance $22528 r0 *1 65.565,133.77
X$22528 251 613 252 644 645 cell_1rw
* cell instance $22529 m0 *1 65.565,136.5
X$22529 251 615 252 644 645 cell_1rw
* cell instance $22530 r0 *1 65.565,136.5
X$22530 251 614 252 644 645 cell_1rw
* cell instance $22531 m0 *1 65.565,139.23
X$22531 251 617 252 644 645 cell_1rw
* cell instance $22532 r0 *1 65.565,139.23
X$22532 251 616 252 644 645 cell_1rw
* cell instance $22533 m0 *1 65.565,141.96
X$22533 251 618 252 644 645 cell_1rw
* cell instance $22534 r0 *1 65.565,141.96
X$22534 251 619 252 644 645 cell_1rw
* cell instance $22535 m0 *1 65.565,144.69
X$22535 251 620 252 644 645 cell_1rw
* cell instance $22536 r0 *1 65.565,144.69
X$22536 251 621 252 644 645 cell_1rw
* cell instance $22537 m0 *1 65.565,147.42
X$22537 251 622 252 644 645 cell_1rw
* cell instance $22538 m0 *1 65.565,150.15
X$22538 251 624 252 644 645 cell_1rw
* cell instance $22539 r0 *1 65.565,147.42
X$22539 251 623 252 644 645 cell_1rw
* cell instance $22540 m0 *1 65.565,152.88
X$22540 251 626 252 644 645 cell_1rw
* cell instance $22541 r0 *1 65.565,150.15
X$22541 251 625 252 644 645 cell_1rw
* cell instance $22542 r0 *1 65.565,152.88
X$22542 251 627 252 644 645 cell_1rw
* cell instance $22543 m0 *1 65.565,155.61
X$22543 251 628 252 644 645 cell_1rw
* cell instance $22544 r0 *1 65.565,155.61
X$22544 251 629 252 644 645 cell_1rw
* cell instance $22545 m0 *1 65.565,158.34
X$22545 251 630 252 644 645 cell_1rw
* cell instance $22546 r0 *1 65.565,158.34
X$22546 251 631 252 644 645 cell_1rw
* cell instance $22547 m0 *1 65.565,161.07
X$22547 251 632 252 644 645 cell_1rw
* cell instance $22548 r0 *1 65.565,161.07
X$22548 251 633 252 644 645 cell_1rw
* cell instance $22549 m0 *1 65.565,163.8
X$22549 251 634 252 644 645 cell_1rw
* cell instance $22550 m0 *1 65.565,166.53
X$22550 251 637 252 644 645 cell_1rw
* cell instance $22551 r0 *1 65.565,163.8
X$22551 251 635 252 644 645 cell_1rw
* cell instance $22552 r0 *1 65.565,166.53
X$22552 251 636 252 644 645 cell_1rw
* cell instance $22553 m0 *1 65.565,169.26
X$22553 251 639 252 644 645 cell_1rw
* cell instance $22554 r0 *1 65.565,169.26
X$22554 251 638 252 644 645 cell_1rw
* cell instance $22555 m0 *1 65.565,171.99
X$22555 251 640 252 644 645 cell_1rw
* cell instance $22556 r0 *1 65.565,171.99
X$22556 251 641 252 644 645 cell_1rw
* cell instance $22557 m0 *1 65.565,174.72
X$22557 251 642 252 644 645 cell_1rw
* cell instance $22558 r0 *1 65.565,174.72
X$22558 251 643 252 644 645 cell_1rw
* cell instance $22559 r0 *1 66.27,87.36
X$22559 253 322 254 644 645 cell_1rw
* cell instance $22560 m0 *1 66.27,90.09
X$22560 253 581 254 644 645 cell_1rw
* cell instance $22561 r0 *1 66.27,90.09
X$22561 253 580 254 644 645 cell_1rw
* cell instance $22562 m0 *1 66.27,92.82
X$22562 253 583 254 644 645 cell_1rw
* cell instance $22563 r0 *1 66.27,92.82
X$22563 253 582 254 644 645 cell_1rw
* cell instance $22564 m0 *1 66.27,95.55
X$22564 253 584 254 644 645 cell_1rw
* cell instance $22565 r0 *1 66.27,95.55
X$22565 253 585 254 644 645 cell_1rw
* cell instance $22566 m0 *1 66.27,98.28
X$22566 253 586 254 644 645 cell_1rw
* cell instance $22567 r0 *1 66.27,98.28
X$22567 253 587 254 644 645 cell_1rw
* cell instance $22568 m0 *1 66.27,101.01
X$22568 253 588 254 644 645 cell_1rw
* cell instance $22569 r0 *1 66.27,101.01
X$22569 253 589 254 644 645 cell_1rw
* cell instance $22570 m0 *1 66.27,103.74
X$22570 253 590 254 644 645 cell_1rw
* cell instance $22571 r0 *1 66.27,103.74
X$22571 253 591 254 644 645 cell_1rw
* cell instance $22572 m0 *1 66.27,106.47
X$22572 253 593 254 644 645 cell_1rw
* cell instance $22573 r0 *1 66.27,106.47
X$22573 253 592 254 644 645 cell_1rw
* cell instance $22574 m0 *1 66.27,109.2
X$22574 253 594 254 644 645 cell_1rw
* cell instance $22575 m0 *1 66.27,111.93
X$22575 253 597 254 644 645 cell_1rw
* cell instance $22576 r0 *1 66.27,109.2
X$22576 253 595 254 644 645 cell_1rw
* cell instance $22577 r0 *1 66.27,111.93
X$22577 253 596 254 644 645 cell_1rw
* cell instance $22578 m0 *1 66.27,114.66
X$22578 253 598 254 644 645 cell_1rw
* cell instance $22579 r0 *1 66.27,114.66
X$22579 253 599 254 644 645 cell_1rw
* cell instance $22580 m0 *1 66.27,117.39
X$22580 253 600 254 644 645 cell_1rw
* cell instance $22581 m0 *1 66.27,120.12
X$22581 253 602 254 644 645 cell_1rw
* cell instance $22582 r0 *1 66.27,117.39
X$22582 253 601 254 644 645 cell_1rw
* cell instance $22583 r0 *1 66.27,120.12
X$22583 253 603 254 644 645 cell_1rw
* cell instance $22584 m0 *1 66.27,122.85
X$22584 253 604 254 644 645 cell_1rw
* cell instance $22585 r0 *1 66.27,122.85
X$22585 253 605 254 644 645 cell_1rw
* cell instance $22586 m0 *1 66.27,125.58
X$22586 253 606 254 644 645 cell_1rw
* cell instance $22587 r0 *1 66.27,125.58
X$22587 253 607 254 644 645 cell_1rw
* cell instance $22588 m0 *1 66.27,128.31
X$22588 253 609 254 644 645 cell_1rw
* cell instance $22589 r0 *1 66.27,128.31
X$22589 253 608 254 644 645 cell_1rw
* cell instance $22590 m0 *1 66.27,131.04
X$22590 253 610 254 644 645 cell_1rw
* cell instance $22591 r0 *1 66.27,131.04
X$22591 253 611 254 644 645 cell_1rw
* cell instance $22592 m0 *1 66.27,133.77
X$22592 253 612 254 644 645 cell_1rw
* cell instance $22593 r0 *1 66.27,133.77
X$22593 253 613 254 644 645 cell_1rw
* cell instance $22594 m0 *1 66.27,136.5
X$22594 253 615 254 644 645 cell_1rw
* cell instance $22595 r0 *1 66.27,136.5
X$22595 253 614 254 644 645 cell_1rw
* cell instance $22596 m0 *1 66.27,139.23
X$22596 253 617 254 644 645 cell_1rw
* cell instance $22597 m0 *1 66.27,141.96
X$22597 253 618 254 644 645 cell_1rw
* cell instance $22598 r0 *1 66.27,139.23
X$22598 253 616 254 644 645 cell_1rw
* cell instance $22599 r0 *1 66.27,141.96
X$22599 253 619 254 644 645 cell_1rw
* cell instance $22600 m0 *1 66.27,144.69
X$22600 253 620 254 644 645 cell_1rw
* cell instance $22601 r0 *1 66.27,144.69
X$22601 253 621 254 644 645 cell_1rw
* cell instance $22602 m0 *1 66.27,147.42
X$22602 253 622 254 644 645 cell_1rw
* cell instance $22603 r0 *1 66.27,147.42
X$22603 253 623 254 644 645 cell_1rw
* cell instance $22604 m0 *1 66.27,150.15
X$22604 253 624 254 644 645 cell_1rw
* cell instance $22605 r0 *1 66.27,150.15
X$22605 253 625 254 644 645 cell_1rw
* cell instance $22606 m0 *1 66.27,152.88
X$22606 253 626 254 644 645 cell_1rw
* cell instance $22607 m0 *1 66.27,155.61
X$22607 253 628 254 644 645 cell_1rw
* cell instance $22608 r0 *1 66.27,152.88
X$22608 253 627 254 644 645 cell_1rw
* cell instance $22609 m0 *1 66.27,158.34
X$22609 253 630 254 644 645 cell_1rw
* cell instance $22610 r0 *1 66.27,155.61
X$22610 253 629 254 644 645 cell_1rw
* cell instance $22611 r0 *1 66.27,158.34
X$22611 253 631 254 644 645 cell_1rw
* cell instance $22612 m0 *1 66.27,161.07
X$22612 253 632 254 644 645 cell_1rw
* cell instance $22613 r0 *1 66.27,161.07
X$22613 253 633 254 644 645 cell_1rw
* cell instance $22614 m0 *1 66.27,163.8
X$22614 253 634 254 644 645 cell_1rw
* cell instance $22615 m0 *1 66.27,166.53
X$22615 253 637 254 644 645 cell_1rw
* cell instance $22616 r0 *1 66.27,163.8
X$22616 253 635 254 644 645 cell_1rw
* cell instance $22617 r0 *1 66.27,166.53
X$22617 253 636 254 644 645 cell_1rw
* cell instance $22618 m0 *1 66.27,169.26
X$22618 253 639 254 644 645 cell_1rw
* cell instance $22619 r0 *1 66.27,169.26
X$22619 253 638 254 644 645 cell_1rw
* cell instance $22620 m0 *1 66.27,171.99
X$22620 253 640 254 644 645 cell_1rw
* cell instance $22621 r0 *1 66.27,171.99
X$22621 253 641 254 644 645 cell_1rw
* cell instance $22622 m0 *1 66.27,174.72
X$22622 253 642 254 644 645 cell_1rw
* cell instance $22623 r0 *1 66.27,174.72
X$22623 253 643 254 644 645 cell_1rw
* cell instance $22624 m0 *1 66.975,90.09
X$22624 255 581 256 644 645 cell_1rw
* cell instance $22625 r0 *1 66.975,87.36
X$22625 255 322 256 644 645 cell_1rw
* cell instance $22626 r0 *1 66.975,90.09
X$22626 255 580 256 644 645 cell_1rw
* cell instance $22627 m0 *1 66.975,92.82
X$22627 255 583 256 644 645 cell_1rw
* cell instance $22628 r0 *1 66.975,92.82
X$22628 255 582 256 644 645 cell_1rw
* cell instance $22629 m0 *1 66.975,95.55
X$22629 255 584 256 644 645 cell_1rw
* cell instance $22630 r0 *1 66.975,95.55
X$22630 255 585 256 644 645 cell_1rw
* cell instance $22631 m0 *1 66.975,98.28
X$22631 255 586 256 644 645 cell_1rw
* cell instance $22632 r0 *1 66.975,98.28
X$22632 255 587 256 644 645 cell_1rw
* cell instance $22633 m0 *1 66.975,101.01
X$22633 255 588 256 644 645 cell_1rw
* cell instance $22634 m0 *1 66.975,103.74
X$22634 255 590 256 644 645 cell_1rw
* cell instance $22635 r0 *1 66.975,101.01
X$22635 255 589 256 644 645 cell_1rw
* cell instance $22636 r0 *1 66.975,103.74
X$22636 255 591 256 644 645 cell_1rw
* cell instance $22637 m0 *1 66.975,106.47
X$22637 255 593 256 644 645 cell_1rw
* cell instance $22638 r0 *1 66.975,106.47
X$22638 255 592 256 644 645 cell_1rw
* cell instance $22639 m0 *1 66.975,109.2
X$22639 255 594 256 644 645 cell_1rw
* cell instance $22640 r0 *1 66.975,109.2
X$22640 255 595 256 644 645 cell_1rw
* cell instance $22641 m0 *1 66.975,111.93
X$22641 255 597 256 644 645 cell_1rw
* cell instance $22642 r0 *1 66.975,111.93
X$22642 255 596 256 644 645 cell_1rw
* cell instance $22643 m0 *1 66.975,114.66
X$22643 255 598 256 644 645 cell_1rw
* cell instance $22644 r0 *1 66.975,114.66
X$22644 255 599 256 644 645 cell_1rw
* cell instance $22645 m0 *1 66.975,117.39
X$22645 255 600 256 644 645 cell_1rw
* cell instance $22646 r0 *1 66.975,117.39
X$22646 255 601 256 644 645 cell_1rw
* cell instance $22647 m0 *1 66.975,120.12
X$22647 255 602 256 644 645 cell_1rw
* cell instance $22648 r0 *1 66.975,120.12
X$22648 255 603 256 644 645 cell_1rw
* cell instance $22649 m0 *1 66.975,122.85
X$22649 255 604 256 644 645 cell_1rw
* cell instance $22650 r0 *1 66.975,122.85
X$22650 255 605 256 644 645 cell_1rw
* cell instance $22651 m0 *1 66.975,125.58
X$22651 255 606 256 644 645 cell_1rw
* cell instance $22652 r0 *1 66.975,125.58
X$22652 255 607 256 644 645 cell_1rw
* cell instance $22653 m0 *1 66.975,128.31
X$22653 255 609 256 644 645 cell_1rw
* cell instance $22654 r0 *1 66.975,128.31
X$22654 255 608 256 644 645 cell_1rw
* cell instance $22655 m0 *1 66.975,131.04
X$22655 255 610 256 644 645 cell_1rw
* cell instance $22656 r0 *1 66.975,131.04
X$22656 255 611 256 644 645 cell_1rw
* cell instance $22657 m0 *1 66.975,133.77
X$22657 255 612 256 644 645 cell_1rw
* cell instance $22658 r0 *1 66.975,133.77
X$22658 255 613 256 644 645 cell_1rw
* cell instance $22659 m0 *1 66.975,136.5
X$22659 255 615 256 644 645 cell_1rw
* cell instance $22660 r0 *1 66.975,136.5
X$22660 255 614 256 644 645 cell_1rw
* cell instance $22661 m0 *1 66.975,139.23
X$22661 255 617 256 644 645 cell_1rw
* cell instance $22662 r0 *1 66.975,139.23
X$22662 255 616 256 644 645 cell_1rw
* cell instance $22663 m0 *1 66.975,141.96
X$22663 255 618 256 644 645 cell_1rw
* cell instance $22664 r0 *1 66.975,141.96
X$22664 255 619 256 644 645 cell_1rw
* cell instance $22665 m0 *1 66.975,144.69
X$22665 255 620 256 644 645 cell_1rw
* cell instance $22666 r0 *1 66.975,144.69
X$22666 255 621 256 644 645 cell_1rw
* cell instance $22667 m0 *1 66.975,147.42
X$22667 255 622 256 644 645 cell_1rw
* cell instance $22668 m0 *1 66.975,150.15
X$22668 255 624 256 644 645 cell_1rw
* cell instance $22669 r0 *1 66.975,147.42
X$22669 255 623 256 644 645 cell_1rw
* cell instance $22670 r0 *1 66.975,150.15
X$22670 255 625 256 644 645 cell_1rw
* cell instance $22671 m0 *1 66.975,152.88
X$22671 255 626 256 644 645 cell_1rw
* cell instance $22672 r0 *1 66.975,152.88
X$22672 255 627 256 644 645 cell_1rw
* cell instance $22673 m0 *1 66.975,155.61
X$22673 255 628 256 644 645 cell_1rw
* cell instance $22674 m0 *1 66.975,158.34
X$22674 255 630 256 644 645 cell_1rw
* cell instance $22675 r0 *1 66.975,155.61
X$22675 255 629 256 644 645 cell_1rw
* cell instance $22676 r0 *1 66.975,158.34
X$22676 255 631 256 644 645 cell_1rw
* cell instance $22677 m0 *1 66.975,161.07
X$22677 255 632 256 644 645 cell_1rw
* cell instance $22678 m0 *1 66.975,163.8
X$22678 255 634 256 644 645 cell_1rw
* cell instance $22679 r0 *1 66.975,161.07
X$22679 255 633 256 644 645 cell_1rw
* cell instance $22680 r0 *1 66.975,163.8
X$22680 255 635 256 644 645 cell_1rw
* cell instance $22681 m0 *1 66.975,166.53
X$22681 255 637 256 644 645 cell_1rw
* cell instance $22682 r0 *1 66.975,166.53
X$22682 255 636 256 644 645 cell_1rw
* cell instance $22683 m0 *1 66.975,169.26
X$22683 255 639 256 644 645 cell_1rw
* cell instance $22684 m0 *1 66.975,171.99
X$22684 255 640 256 644 645 cell_1rw
* cell instance $22685 r0 *1 66.975,169.26
X$22685 255 638 256 644 645 cell_1rw
* cell instance $22686 m0 *1 66.975,174.72
X$22686 255 642 256 644 645 cell_1rw
* cell instance $22687 r0 *1 66.975,171.99
X$22687 255 641 256 644 645 cell_1rw
* cell instance $22688 r0 *1 66.975,174.72
X$22688 255 643 256 644 645 cell_1rw
* cell instance $22689 m0 *1 67.68,90.09
X$22689 257 581 258 644 645 cell_1rw
* cell instance $22690 r0 *1 67.68,87.36
X$22690 257 322 258 644 645 cell_1rw
* cell instance $22691 r0 *1 67.68,90.09
X$22691 257 580 258 644 645 cell_1rw
* cell instance $22692 m0 *1 67.68,92.82
X$22692 257 583 258 644 645 cell_1rw
* cell instance $22693 m0 *1 67.68,95.55
X$22693 257 584 258 644 645 cell_1rw
* cell instance $22694 r0 *1 67.68,92.82
X$22694 257 582 258 644 645 cell_1rw
* cell instance $22695 m0 *1 67.68,98.28
X$22695 257 586 258 644 645 cell_1rw
* cell instance $22696 r0 *1 67.68,95.55
X$22696 257 585 258 644 645 cell_1rw
* cell instance $22697 r0 *1 67.68,98.28
X$22697 257 587 258 644 645 cell_1rw
* cell instance $22698 m0 *1 67.68,101.01
X$22698 257 588 258 644 645 cell_1rw
* cell instance $22699 r0 *1 67.68,101.01
X$22699 257 589 258 644 645 cell_1rw
* cell instance $22700 m0 *1 67.68,103.74
X$22700 257 590 258 644 645 cell_1rw
* cell instance $22701 r0 *1 67.68,103.74
X$22701 257 591 258 644 645 cell_1rw
* cell instance $22702 m0 *1 67.68,106.47
X$22702 257 593 258 644 645 cell_1rw
* cell instance $22703 r0 *1 67.68,106.47
X$22703 257 592 258 644 645 cell_1rw
* cell instance $22704 m0 *1 67.68,109.2
X$22704 257 594 258 644 645 cell_1rw
* cell instance $22705 r0 *1 67.68,109.2
X$22705 257 595 258 644 645 cell_1rw
* cell instance $22706 m0 *1 67.68,111.93
X$22706 257 597 258 644 645 cell_1rw
* cell instance $22707 r0 *1 67.68,111.93
X$22707 257 596 258 644 645 cell_1rw
* cell instance $22708 m0 *1 67.68,114.66
X$22708 257 598 258 644 645 cell_1rw
* cell instance $22709 r0 *1 67.68,114.66
X$22709 257 599 258 644 645 cell_1rw
* cell instance $22710 m0 *1 67.68,117.39
X$22710 257 600 258 644 645 cell_1rw
* cell instance $22711 r0 *1 67.68,117.39
X$22711 257 601 258 644 645 cell_1rw
* cell instance $22712 m0 *1 67.68,120.12
X$22712 257 602 258 644 645 cell_1rw
* cell instance $22713 r0 *1 67.68,120.12
X$22713 257 603 258 644 645 cell_1rw
* cell instance $22714 m0 *1 67.68,122.85
X$22714 257 604 258 644 645 cell_1rw
* cell instance $22715 r0 *1 67.68,122.85
X$22715 257 605 258 644 645 cell_1rw
* cell instance $22716 m0 *1 67.68,125.58
X$22716 257 606 258 644 645 cell_1rw
* cell instance $22717 m0 *1 67.68,128.31
X$22717 257 609 258 644 645 cell_1rw
* cell instance $22718 r0 *1 67.68,125.58
X$22718 257 607 258 644 645 cell_1rw
* cell instance $22719 r0 *1 67.68,128.31
X$22719 257 608 258 644 645 cell_1rw
* cell instance $22720 m0 *1 67.68,131.04
X$22720 257 610 258 644 645 cell_1rw
* cell instance $22721 r0 *1 67.68,131.04
X$22721 257 611 258 644 645 cell_1rw
* cell instance $22722 m0 *1 67.68,133.77
X$22722 257 612 258 644 645 cell_1rw
* cell instance $22723 r0 *1 67.68,133.77
X$22723 257 613 258 644 645 cell_1rw
* cell instance $22724 m0 *1 67.68,136.5
X$22724 257 615 258 644 645 cell_1rw
* cell instance $22725 r0 *1 67.68,136.5
X$22725 257 614 258 644 645 cell_1rw
* cell instance $22726 m0 *1 67.68,139.23
X$22726 257 617 258 644 645 cell_1rw
* cell instance $22727 r0 *1 67.68,139.23
X$22727 257 616 258 644 645 cell_1rw
* cell instance $22728 m0 *1 67.68,141.96
X$22728 257 618 258 644 645 cell_1rw
* cell instance $22729 r0 *1 67.68,141.96
X$22729 257 619 258 644 645 cell_1rw
* cell instance $22730 m0 *1 67.68,144.69
X$22730 257 620 258 644 645 cell_1rw
* cell instance $22731 m0 *1 67.68,147.42
X$22731 257 622 258 644 645 cell_1rw
* cell instance $22732 r0 *1 67.68,144.69
X$22732 257 621 258 644 645 cell_1rw
* cell instance $22733 m0 *1 67.68,150.15
X$22733 257 624 258 644 645 cell_1rw
* cell instance $22734 r0 *1 67.68,147.42
X$22734 257 623 258 644 645 cell_1rw
* cell instance $22735 m0 *1 67.68,152.88
X$22735 257 626 258 644 645 cell_1rw
* cell instance $22736 r0 *1 67.68,150.15
X$22736 257 625 258 644 645 cell_1rw
* cell instance $22737 r0 *1 67.68,152.88
X$22737 257 627 258 644 645 cell_1rw
* cell instance $22738 m0 *1 67.68,155.61
X$22738 257 628 258 644 645 cell_1rw
* cell instance $22739 m0 *1 67.68,158.34
X$22739 257 630 258 644 645 cell_1rw
* cell instance $22740 r0 *1 67.68,155.61
X$22740 257 629 258 644 645 cell_1rw
* cell instance $22741 r0 *1 67.68,158.34
X$22741 257 631 258 644 645 cell_1rw
* cell instance $22742 m0 *1 67.68,161.07
X$22742 257 632 258 644 645 cell_1rw
* cell instance $22743 m0 *1 67.68,163.8
X$22743 257 634 258 644 645 cell_1rw
* cell instance $22744 r0 *1 67.68,161.07
X$22744 257 633 258 644 645 cell_1rw
* cell instance $22745 r0 *1 67.68,163.8
X$22745 257 635 258 644 645 cell_1rw
* cell instance $22746 m0 *1 67.68,166.53
X$22746 257 637 258 644 645 cell_1rw
* cell instance $22747 m0 *1 67.68,169.26
X$22747 257 639 258 644 645 cell_1rw
* cell instance $22748 r0 *1 67.68,166.53
X$22748 257 636 258 644 645 cell_1rw
* cell instance $22749 r0 *1 67.68,169.26
X$22749 257 638 258 644 645 cell_1rw
* cell instance $22750 m0 *1 67.68,171.99
X$22750 257 640 258 644 645 cell_1rw
* cell instance $22751 r0 *1 67.68,171.99
X$22751 257 641 258 644 645 cell_1rw
* cell instance $22752 m0 *1 67.68,174.72
X$22752 257 642 258 644 645 cell_1rw
* cell instance $22753 r0 *1 67.68,174.72
X$22753 257 643 258 644 645 cell_1rw
* cell instance $22754 r0 *1 68.385,87.36
X$22754 259 322 260 644 645 cell_1rw
* cell instance $22755 m0 *1 68.385,90.09
X$22755 259 581 260 644 645 cell_1rw
* cell instance $22756 m0 *1 68.385,92.82
X$22756 259 583 260 644 645 cell_1rw
* cell instance $22757 r0 *1 68.385,90.09
X$22757 259 580 260 644 645 cell_1rw
* cell instance $22758 r0 *1 68.385,92.82
X$22758 259 582 260 644 645 cell_1rw
* cell instance $22759 m0 *1 68.385,95.55
X$22759 259 584 260 644 645 cell_1rw
* cell instance $22760 m0 *1 68.385,98.28
X$22760 259 586 260 644 645 cell_1rw
* cell instance $22761 r0 *1 68.385,95.55
X$22761 259 585 260 644 645 cell_1rw
* cell instance $22762 m0 *1 68.385,101.01
X$22762 259 588 260 644 645 cell_1rw
* cell instance $22763 r0 *1 68.385,98.28
X$22763 259 587 260 644 645 cell_1rw
* cell instance $22764 r0 *1 68.385,101.01
X$22764 259 589 260 644 645 cell_1rw
* cell instance $22765 m0 *1 68.385,103.74
X$22765 259 590 260 644 645 cell_1rw
* cell instance $22766 m0 *1 68.385,106.47
X$22766 259 593 260 644 645 cell_1rw
* cell instance $22767 r0 *1 68.385,103.74
X$22767 259 591 260 644 645 cell_1rw
* cell instance $22768 r0 *1 68.385,106.47
X$22768 259 592 260 644 645 cell_1rw
* cell instance $22769 m0 *1 68.385,109.2
X$22769 259 594 260 644 645 cell_1rw
* cell instance $22770 r0 *1 68.385,109.2
X$22770 259 595 260 644 645 cell_1rw
* cell instance $22771 m0 *1 68.385,111.93
X$22771 259 597 260 644 645 cell_1rw
* cell instance $22772 r0 *1 68.385,111.93
X$22772 259 596 260 644 645 cell_1rw
* cell instance $22773 m0 *1 68.385,114.66
X$22773 259 598 260 644 645 cell_1rw
* cell instance $22774 r0 *1 68.385,114.66
X$22774 259 599 260 644 645 cell_1rw
* cell instance $22775 m0 *1 68.385,117.39
X$22775 259 600 260 644 645 cell_1rw
* cell instance $22776 r0 *1 68.385,117.39
X$22776 259 601 260 644 645 cell_1rw
* cell instance $22777 m0 *1 68.385,120.12
X$22777 259 602 260 644 645 cell_1rw
* cell instance $22778 r0 *1 68.385,120.12
X$22778 259 603 260 644 645 cell_1rw
* cell instance $22779 m0 *1 68.385,122.85
X$22779 259 604 260 644 645 cell_1rw
* cell instance $22780 r0 *1 68.385,122.85
X$22780 259 605 260 644 645 cell_1rw
* cell instance $22781 m0 *1 68.385,125.58
X$22781 259 606 260 644 645 cell_1rw
* cell instance $22782 r0 *1 68.385,125.58
X$22782 259 607 260 644 645 cell_1rw
* cell instance $22783 m0 *1 68.385,128.31
X$22783 259 609 260 644 645 cell_1rw
* cell instance $22784 m0 *1 68.385,131.04
X$22784 259 610 260 644 645 cell_1rw
* cell instance $22785 r0 *1 68.385,128.31
X$22785 259 608 260 644 645 cell_1rw
* cell instance $22786 r0 *1 68.385,131.04
X$22786 259 611 260 644 645 cell_1rw
* cell instance $22787 m0 *1 68.385,133.77
X$22787 259 612 260 644 645 cell_1rw
* cell instance $22788 r0 *1 68.385,133.77
X$22788 259 613 260 644 645 cell_1rw
* cell instance $22789 m0 *1 68.385,136.5
X$22789 259 615 260 644 645 cell_1rw
* cell instance $22790 m0 *1 68.385,139.23
X$22790 259 617 260 644 645 cell_1rw
* cell instance $22791 r0 *1 68.385,136.5
X$22791 259 614 260 644 645 cell_1rw
* cell instance $22792 r0 *1 68.385,139.23
X$22792 259 616 260 644 645 cell_1rw
* cell instance $22793 m0 *1 68.385,141.96
X$22793 259 618 260 644 645 cell_1rw
* cell instance $22794 r0 *1 68.385,141.96
X$22794 259 619 260 644 645 cell_1rw
* cell instance $22795 m0 *1 68.385,144.69
X$22795 259 620 260 644 645 cell_1rw
* cell instance $22796 r0 *1 68.385,144.69
X$22796 259 621 260 644 645 cell_1rw
* cell instance $22797 m0 *1 68.385,147.42
X$22797 259 622 260 644 645 cell_1rw
* cell instance $22798 m0 *1 68.385,150.15
X$22798 259 624 260 644 645 cell_1rw
* cell instance $22799 r0 *1 68.385,147.42
X$22799 259 623 260 644 645 cell_1rw
* cell instance $22800 r0 *1 68.385,150.15
X$22800 259 625 260 644 645 cell_1rw
* cell instance $22801 m0 *1 68.385,152.88
X$22801 259 626 260 644 645 cell_1rw
* cell instance $22802 m0 *1 68.385,155.61
X$22802 259 628 260 644 645 cell_1rw
* cell instance $22803 r0 *1 68.385,152.88
X$22803 259 627 260 644 645 cell_1rw
* cell instance $22804 r0 *1 68.385,155.61
X$22804 259 629 260 644 645 cell_1rw
* cell instance $22805 m0 *1 68.385,158.34
X$22805 259 630 260 644 645 cell_1rw
* cell instance $22806 m0 *1 68.385,161.07
X$22806 259 632 260 644 645 cell_1rw
* cell instance $22807 r0 *1 68.385,158.34
X$22807 259 631 260 644 645 cell_1rw
* cell instance $22808 r0 *1 68.385,161.07
X$22808 259 633 260 644 645 cell_1rw
* cell instance $22809 m0 *1 68.385,163.8
X$22809 259 634 260 644 645 cell_1rw
* cell instance $22810 r0 *1 68.385,163.8
X$22810 259 635 260 644 645 cell_1rw
* cell instance $22811 m0 *1 68.385,166.53
X$22811 259 637 260 644 645 cell_1rw
* cell instance $22812 m0 *1 68.385,169.26
X$22812 259 639 260 644 645 cell_1rw
* cell instance $22813 r0 *1 68.385,166.53
X$22813 259 636 260 644 645 cell_1rw
* cell instance $22814 m0 *1 68.385,171.99
X$22814 259 640 260 644 645 cell_1rw
* cell instance $22815 r0 *1 68.385,169.26
X$22815 259 638 260 644 645 cell_1rw
* cell instance $22816 m0 *1 68.385,174.72
X$22816 259 642 260 644 645 cell_1rw
* cell instance $22817 r0 *1 68.385,171.99
X$22817 259 641 260 644 645 cell_1rw
* cell instance $22818 r0 *1 68.385,174.72
X$22818 259 643 260 644 645 cell_1rw
* cell instance $22819 r0 *1 69.09,87.36
X$22819 261 322 262 644 645 cell_1rw
* cell instance $22820 m0 *1 69.09,90.09
X$22820 261 581 262 644 645 cell_1rw
* cell instance $22821 r0 *1 69.09,90.09
X$22821 261 580 262 644 645 cell_1rw
* cell instance $22822 m0 *1 69.09,92.82
X$22822 261 583 262 644 645 cell_1rw
* cell instance $22823 r0 *1 69.09,92.82
X$22823 261 582 262 644 645 cell_1rw
* cell instance $22824 m0 *1 69.09,95.55
X$22824 261 584 262 644 645 cell_1rw
* cell instance $22825 r0 *1 69.09,95.55
X$22825 261 585 262 644 645 cell_1rw
* cell instance $22826 m0 *1 69.09,98.28
X$22826 261 586 262 644 645 cell_1rw
* cell instance $22827 r0 *1 69.09,98.28
X$22827 261 587 262 644 645 cell_1rw
* cell instance $22828 m0 *1 69.09,101.01
X$22828 261 588 262 644 645 cell_1rw
* cell instance $22829 r0 *1 69.09,101.01
X$22829 261 589 262 644 645 cell_1rw
* cell instance $22830 m0 *1 69.09,103.74
X$22830 261 590 262 644 645 cell_1rw
* cell instance $22831 r0 *1 69.09,103.74
X$22831 261 591 262 644 645 cell_1rw
* cell instance $22832 m0 *1 69.09,106.47
X$22832 261 593 262 644 645 cell_1rw
* cell instance $22833 r0 *1 69.09,106.47
X$22833 261 592 262 644 645 cell_1rw
* cell instance $22834 m0 *1 69.09,109.2
X$22834 261 594 262 644 645 cell_1rw
* cell instance $22835 r0 *1 69.09,109.2
X$22835 261 595 262 644 645 cell_1rw
* cell instance $22836 m0 *1 69.09,111.93
X$22836 261 597 262 644 645 cell_1rw
* cell instance $22837 r0 *1 69.09,111.93
X$22837 261 596 262 644 645 cell_1rw
* cell instance $22838 m0 *1 69.09,114.66
X$22838 261 598 262 644 645 cell_1rw
* cell instance $22839 r0 *1 69.09,114.66
X$22839 261 599 262 644 645 cell_1rw
* cell instance $22840 m0 *1 69.09,117.39
X$22840 261 600 262 644 645 cell_1rw
* cell instance $22841 r0 *1 69.09,117.39
X$22841 261 601 262 644 645 cell_1rw
* cell instance $22842 m0 *1 69.09,120.12
X$22842 261 602 262 644 645 cell_1rw
* cell instance $22843 r0 *1 69.09,120.12
X$22843 261 603 262 644 645 cell_1rw
* cell instance $22844 m0 *1 69.09,122.85
X$22844 261 604 262 644 645 cell_1rw
* cell instance $22845 r0 *1 69.09,122.85
X$22845 261 605 262 644 645 cell_1rw
* cell instance $22846 m0 *1 69.09,125.58
X$22846 261 606 262 644 645 cell_1rw
* cell instance $22847 r0 *1 69.09,125.58
X$22847 261 607 262 644 645 cell_1rw
* cell instance $22848 m0 *1 69.09,128.31
X$22848 261 609 262 644 645 cell_1rw
* cell instance $22849 r0 *1 69.09,128.31
X$22849 261 608 262 644 645 cell_1rw
* cell instance $22850 m0 *1 69.09,131.04
X$22850 261 610 262 644 645 cell_1rw
* cell instance $22851 m0 *1 69.09,133.77
X$22851 261 612 262 644 645 cell_1rw
* cell instance $22852 r0 *1 69.09,131.04
X$22852 261 611 262 644 645 cell_1rw
* cell instance $22853 r0 *1 69.09,133.77
X$22853 261 613 262 644 645 cell_1rw
* cell instance $22854 m0 *1 69.09,136.5
X$22854 261 615 262 644 645 cell_1rw
* cell instance $22855 r0 *1 69.09,136.5
X$22855 261 614 262 644 645 cell_1rw
* cell instance $22856 m0 *1 69.09,139.23
X$22856 261 617 262 644 645 cell_1rw
* cell instance $22857 m0 *1 69.09,141.96
X$22857 261 618 262 644 645 cell_1rw
* cell instance $22858 r0 *1 69.09,139.23
X$22858 261 616 262 644 645 cell_1rw
* cell instance $22859 r0 *1 69.09,141.96
X$22859 261 619 262 644 645 cell_1rw
* cell instance $22860 m0 *1 69.09,144.69
X$22860 261 620 262 644 645 cell_1rw
* cell instance $22861 m0 *1 69.09,147.42
X$22861 261 622 262 644 645 cell_1rw
* cell instance $22862 r0 *1 69.09,144.69
X$22862 261 621 262 644 645 cell_1rw
* cell instance $22863 m0 *1 69.09,150.15
X$22863 261 624 262 644 645 cell_1rw
* cell instance $22864 r0 *1 69.09,147.42
X$22864 261 623 262 644 645 cell_1rw
* cell instance $22865 r0 *1 69.09,150.15
X$22865 261 625 262 644 645 cell_1rw
* cell instance $22866 m0 *1 69.09,152.88
X$22866 261 626 262 644 645 cell_1rw
* cell instance $22867 r0 *1 69.09,152.88
X$22867 261 627 262 644 645 cell_1rw
* cell instance $22868 m0 *1 69.09,155.61
X$22868 261 628 262 644 645 cell_1rw
* cell instance $22869 r0 *1 69.09,155.61
X$22869 261 629 262 644 645 cell_1rw
* cell instance $22870 m0 *1 69.09,158.34
X$22870 261 630 262 644 645 cell_1rw
* cell instance $22871 r0 *1 69.09,158.34
X$22871 261 631 262 644 645 cell_1rw
* cell instance $22872 m0 *1 69.09,161.07
X$22872 261 632 262 644 645 cell_1rw
* cell instance $22873 m0 *1 69.09,163.8
X$22873 261 634 262 644 645 cell_1rw
* cell instance $22874 r0 *1 69.09,161.07
X$22874 261 633 262 644 645 cell_1rw
* cell instance $22875 r0 *1 69.09,163.8
X$22875 261 635 262 644 645 cell_1rw
* cell instance $22876 m0 *1 69.09,166.53
X$22876 261 637 262 644 645 cell_1rw
* cell instance $22877 r0 *1 69.09,166.53
X$22877 261 636 262 644 645 cell_1rw
* cell instance $22878 m0 *1 69.09,169.26
X$22878 261 639 262 644 645 cell_1rw
* cell instance $22879 r0 *1 69.09,169.26
X$22879 261 638 262 644 645 cell_1rw
* cell instance $22880 m0 *1 69.09,171.99
X$22880 261 640 262 644 645 cell_1rw
* cell instance $22881 r0 *1 69.09,171.99
X$22881 261 641 262 644 645 cell_1rw
* cell instance $22882 m0 *1 69.09,174.72
X$22882 261 642 262 644 645 cell_1rw
* cell instance $22883 r0 *1 69.09,174.72
X$22883 261 643 262 644 645 cell_1rw
* cell instance $22884 r0 *1 69.795,87.36
X$22884 263 322 264 644 645 cell_1rw
* cell instance $22885 m0 *1 69.795,90.09
X$22885 263 581 264 644 645 cell_1rw
* cell instance $22886 r0 *1 69.795,90.09
X$22886 263 580 264 644 645 cell_1rw
* cell instance $22887 m0 *1 69.795,92.82
X$22887 263 583 264 644 645 cell_1rw
* cell instance $22888 m0 *1 69.795,95.55
X$22888 263 584 264 644 645 cell_1rw
* cell instance $22889 r0 *1 69.795,92.82
X$22889 263 582 264 644 645 cell_1rw
* cell instance $22890 m0 *1 69.795,98.28
X$22890 263 586 264 644 645 cell_1rw
* cell instance $22891 r0 *1 69.795,95.55
X$22891 263 585 264 644 645 cell_1rw
* cell instance $22892 r0 *1 69.795,98.28
X$22892 263 587 264 644 645 cell_1rw
* cell instance $22893 m0 *1 69.795,101.01
X$22893 263 588 264 644 645 cell_1rw
* cell instance $22894 r0 *1 69.795,101.01
X$22894 263 589 264 644 645 cell_1rw
* cell instance $22895 m0 *1 69.795,103.74
X$22895 263 590 264 644 645 cell_1rw
* cell instance $22896 r0 *1 69.795,103.74
X$22896 263 591 264 644 645 cell_1rw
* cell instance $22897 m0 *1 69.795,106.47
X$22897 263 593 264 644 645 cell_1rw
* cell instance $22898 m0 *1 69.795,109.2
X$22898 263 594 264 644 645 cell_1rw
* cell instance $22899 r0 *1 69.795,106.47
X$22899 263 592 264 644 645 cell_1rw
* cell instance $22900 m0 *1 69.795,111.93
X$22900 263 597 264 644 645 cell_1rw
* cell instance $22901 r0 *1 69.795,109.2
X$22901 263 595 264 644 645 cell_1rw
* cell instance $22902 r0 *1 69.795,111.93
X$22902 263 596 264 644 645 cell_1rw
* cell instance $22903 m0 *1 69.795,114.66
X$22903 263 598 264 644 645 cell_1rw
* cell instance $22904 r0 *1 69.795,114.66
X$22904 263 599 264 644 645 cell_1rw
* cell instance $22905 m0 *1 69.795,117.39
X$22905 263 600 264 644 645 cell_1rw
* cell instance $22906 r0 *1 69.795,117.39
X$22906 263 601 264 644 645 cell_1rw
* cell instance $22907 m0 *1 69.795,120.12
X$22907 263 602 264 644 645 cell_1rw
* cell instance $22908 r0 *1 69.795,120.12
X$22908 263 603 264 644 645 cell_1rw
* cell instance $22909 m0 *1 69.795,122.85
X$22909 263 604 264 644 645 cell_1rw
* cell instance $22910 m0 *1 69.795,125.58
X$22910 263 606 264 644 645 cell_1rw
* cell instance $22911 r0 *1 69.795,122.85
X$22911 263 605 264 644 645 cell_1rw
* cell instance $22912 r0 *1 69.795,125.58
X$22912 263 607 264 644 645 cell_1rw
* cell instance $22913 m0 *1 69.795,128.31
X$22913 263 609 264 644 645 cell_1rw
* cell instance $22914 m0 *1 69.795,131.04
X$22914 263 610 264 644 645 cell_1rw
* cell instance $22915 r0 *1 69.795,128.31
X$22915 263 608 264 644 645 cell_1rw
* cell instance $22916 r0 *1 69.795,131.04
X$22916 263 611 264 644 645 cell_1rw
* cell instance $22917 m0 *1 69.795,133.77
X$22917 263 612 264 644 645 cell_1rw
* cell instance $22918 r0 *1 69.795,133.77
X$22918 263 613 264 644 645 cell_1rw
* cell instance $22919 m0 *1 69.795,136.5
X$22919 263 615 264 644 645 cell_1rw
* cell instance $22920 m0 *1 69.795,139.23
X$22920 263 617 264 644 645 cell_1rw
* cell instance $22921 r0 *1 69.795,136.5
X$22921 263 614 264 644 645 cell_1rw
* cell instance $22922 r0 *1 69.795,139.23
X$22922 263 616 264 644 645 cell_1rw
* cell instance $22923 m0 *1 69.795,141.96
X$22923 263 618 264 644 645 cell_1rw
* cell instance $22924 m0 *1 69.795,144.69
X$22924 263 620 264 644 645 cell_1rw
* cell instance $22925 r0 *1 69.795,141.96
X$22925 263 619 264 644 645 cell_1rw
* cell instance $22926 r0 *1 69.795,144.69
X$22926 263 621 264 644 645 cell_1rw
* cell instance $22927 m0 *1 69.795,147.42
X$22927 263 622 264 644 645 cell_1rw
* cell instance $22928 r0 *1 69.795,147.42
X$22928 263 623 264 644 645 cell_1rw
* cell instance $22929 m0 *1 69.795,150.15
X$22929 263 624 264 644 645 cell_1rw
* cell instance $22930 r0 *1 69.795,150.15
X$22930 263 625 264 644 645 cell_1rw
* cell instance $22931 m0 *1 69.795,152.88
X$22931 263 626 264 644 645 cell_1rw
* cell instance $22932 m0 *1 69.795,155.61
X$22932 263 628 264 644 645 cell_1rw
* cell instance $22933 r0 *1 69.795,152.88
X$22933 263 627 264 644 645 cell_1rw
* cell instance $22934 m0 *1 69.795,158.34
X$22934 263 630 264 644 645 cell_1rw
* cell instance $22935 r0 *1 69.795,155.61
X$22935 263 629 264 644 645 cell_1rw
* cell instance $22936 r0 *1 69.795,158.34
X$22936 263 631 264 644 645 cell_1rw
* cell instance $22937 m0 *1 69.795,161.07
X$22937 263 632 264 644 645 cell_1rw
* cell instance $22938 r0 *1 69.795,161.07
X$22938 263 633 264 644 645 cell_1rw
* cell instance $22939 m0 *1 69.795,163.8
X$22939 263 634 264 644 645 cell_1rw
* cell instance $22940 r0 *1 69.795,163.8
X$22940 263 635 264 644 645 cell_1rw
* cell instance $22941 m0 *1 69.795,166.53
X$22941 263 637 264 644 645 cell_1rw
* cell instance $22942 r0 *1 69.795,166.53
X$22942 263 636 264 644 645 cell_1rw
* cell instance $22943 m0 *1 69.795,169.26
X$22943 263 639 264 644 645 cell_1rw
* cell instance $22944 r0 *1 69.795,169.26
X$22944 263 638 264 644 645 cell_1rw
* cell instance $22945 m0 *1 69.795,171.99
X$22945 263 640 264 644 645 cell_1rw
* cell instance $22946 r0 *1 69.795,171.99
X$22946 263 641 264 644 645 cell_1rw
* cell instance $22947 m0 *1 69.795,174.72
X$22947 263 642 264 644 645 cell_1rw
* cell instance $22948 r0 *1 69.795,174.72
X$22948 263 643 264 644 645 cell_1rw
* cell instance $22949 m0 *1 70.5,90.09
X$22949 265 581 266 644 645 cell_1rw
* cell instance $22950 r0 *1 70.5,87.36
X$22950 265 322 266 644 645 cell_1rw
* cell instance $22951 r0 *1 70.5,90.09
X$22951 265 580 266 644 645 cell_1rw
* cell instance $22952 m0 *1 70.5,92.82
X$22952 265 583 266 644 645 cell_1rw
* cell instance $22953 m0 *1 70.5,95.55
X$22953 265 584 266 644 645 cell_1rw
* cell instance $22954 r0 *1 70.5,92.82
X$22954 265 582 266 644 645 cell_1rw
* cell instance $22955 r0 *1 70.5,95.55
X$22955 265 585 266 644 645 cell_1rw
* cell instance $22956 m0 *1 70.5,98.28
X$22956 265 586 266 644 645 cell_1rw
* cell instance $22957 m0 *1 70.5,101.01
X$22957 265 588 266 644 645 cell_1rw
* cell instance $22958 r0 *1 70.5,98.28
X$22958 265 587 266 644 645 cell_1rw
* cell instance $22959 m0 *1 70.5,103.74
X$22959 265 590 266 644 645 cell_1rw
* cell instance $22960 r0 *1 70.5,101.01
X$22960 265 589 266 644 645 cell_1rw
* cell instance $22961 r0 *1 70.5,103.74
X$22961 265 591 266 644 645 cell_1rw
* cell instance $22962 m0 *1 70.5,106.47
X$22962 265 593 266 644 645 cell_1rw
* cell instance $22963 r0 *1 70.5,106.47
X$22963 265 592 266 644 645 cell_1rw
* cell instance $22964 m0 *1 70.5,109.2
X$22964 265 594 266 644 645 cell_1rw
* cell instance $22965 r0 *1 70.5,109.2
X$22965 265 595 266 644 645 cell_1rw
* cell instance $22966 m0 *1 70.5,111.93
X$22966 265 597 266 644 645 cell_1rw
* cell instance $22967 r0 *1 70.5,111.93
X$22967 265 596 266 644 645 cell_1rw
* cell instance $22968 m0 *1 70.5,114.66
X$22968 265 598 266 644 645 cell_1rw
* cell instance $22969 r0 *1 70.5,114.66
X$22969 265 599 266 644 645 cell_1rw
* cell instance $22970 m0 *1 70.5,117.39
X$22970 265 600 266 644 645 cell_1rw
* cell instance $22971 r0 *1 70.5,117.39
X$22971 265 601 266 644 645 cell_1rw
* cell instance $22972 m0 *1 70.5,120.12
X$22972 265 602 266 644 645 cell_1rw
* cell instance $22973 r0 *1 70.5,120.12
X$22973 265 603 266 644 645 cell_1rw
* cell instance $22974 m0 *1 70.5,122.85
X$22974 265 604 266 644 645 cell_1rw
* cell instance $22975 r0 *1 70.5,122.85
X$22975 265 605 266 644 645 cell_1rw
* cell instance $22976 m0 *1 70.5,125.58
X$22976 265 606 266 644 645 cell_1rw
* cell instance $22977 r0 *1 70.5,125.58
X$22977 265 607 266 644 645 cell_1rw
* cell instance $22978 m0 *1 70.5,128.31
X$22978 265 609 266 644 645 cell_1rw
* cell instance $22979 r0 *1 70.5,128.31
X$22979 265 608 266 644 645 cell_1rw
* cell instance $22980 m0 *1 70.5,131.04
X$22980 265 610 266 644 645 cell_1rw
* cell instance $22981 r0 *1 70.5,131.04
X$22981 265 611 266 644 645 cell_1rw
* cell instance $22982 m0 *1 70.5,133.77
X$22982 265 612 266 644 645 cell_1rw
* cell instance $22983 m0 *1 70.5,136.5
X$22983 265 615 266 644 645 cell_1rw
* cell instance $22984 r0 *1 70.5,133.77
X$22984 265 613 266 644 645 cell_1rw
* cell instance $22985 r0 *1 70.5,136.5
X$22985 265 614 266 644 645 cell_1rw
* cell instance $22986 m0 *1 70.5,139.23
X$22986 265 617 266 644 645 cell_1rw
* cell instance $22987 r0 *1 70.5,139.23
X$22987 265 616 266 644 645 cell_1rw
* cell instance $22988 m0 *1 70.5,141.96
X$22988 265 618 266 644 645 cell_1rw
* cell instance $22989 m0 *1 70.5,144.69
X$22989 265 620 266 644 645 cell_1rw
* cell instance $22990 r0 *1 70.5,141.96
X$22990 265 619 266 644 645 cell_1rw
* cell instance $22991 r0 *1 70.5,144.69
X$22991 265 621 266 644 645 cell_1rw
* cell instance $22992 m0 *1 70.5,147.42
X$22992 265 622 266 644 645 cell_1rw
* cell instance $22993 r0 *1 70.5,147.42
X$22993 265 623 266 644 645 cell_1rw
* cell instance $22994 m0 *1 70.5,150.15
X$22994 265 624 266 644 645 cell_1rw
* cell instance $22995 r0 *1 70.5,150.15
X$22995 265 625 266 644 645 cell_1rw
* cell instance $22996 m0 *1 70.5,152.88
X$22996 265 626 266 644 645 cell_1rw
* cell instance $22997 r0 *1 70.5,152.88
X$22997 265 627 266 644 645 cell_1rw
* cell instance $22998 m0 *1 70.5,155.61
X$22998 265 628 266 644 645 cell_1rw
* cell instance $22999 r0 *1 70.5,155.61
X$22999 265 629 266 644 645 cell_1rw
* cell instance $23000 m0 *1 70.5,158.34
X$23000 265 630 266 644 645 cell_1rw
* cell instance $23001 r0 *1 70.5,158.34
X$23001 265 631 266 644 645 cell_1rw
* cell instance $23002 m0 *1 70.5,161.07
X$23002 265 632 266 644 645 cell_1rw
* cell instance $23003 r0 *1 70.5,161.07
X$23003 265 633 266 644 645 cell_1rw
* cell instance $23004 m0 *1 70.5,163.8
X$23004 265 634 266 644 645 cell_1rw
* cell instance $23005 r0 *1 70.5,163.8
X$23005 265 635 266 644 645 cell_1rw
* cell instance $23006 m0 *1 70.5,166.53
X$23006 265 637 266 644 645 cell_1rw
* cell instance $23007 r0 *1 70.5,166.53
X$23007 265 636 266 644 645 cell_1rw
* cell instance $23008 m0 *1 70.5,169.26
X$23008 265 639 266 644 645 cell_1rw
* cell instance $23009 r0 *1 70.5,169.26
X$23009 265 638 266 644 645 cell_1rw
* cell instance $23010 m0 *1 70.5,171.99
X$23010 265 640 266 644 645 cell_1rw
* cell instance $23011 r0 *1 70.5,171.99
X$23011 265 641 266 644 645 cell_1rw
* cell instance $23012 m0 *1 70.5,174.72
X$23012 265 642 266 644 645 cell_1rw
* cell instance $23013 r0 *1 70.5,174.72
X$23013 265 643 266 644 645 cell_1rw
* cell instance $23014 r0 *1 71.205,87.36
X$23014 267 322 268 644 645 cell_1rw
* cell instance $23015 m0 *1 71.205,90.09
X$23015 267 581 268 644 645 cell_1rw
* cell instance $23016 r0 *1 71.205,90.09
X$23016 267 580 268 644 645 cell_1rw
* cell instance $23017 m0 *1 71.205,92.82
X$23017 267 583 268 644 645 cell_1rw
* cell instance $23018 r0 *1 71.205,92.82
X$23018 267 582 268 644 645 cell_1rw
* cell instance $23019 m0 *1 71.205,95.55
X$23019 267 584 268 644 645 cell_1rw
* cell instance $23020 r0 *1 71.205,95.55
X$23020 267 585 268 644 645 cell_1rw
* cell instance $23021 m0 *1 71.205,98.28
X$23021 267 586 268 644 645 cell_1rw
* cell instance $23022 r0 *1 71.205,98.28
X$23022 267 587 268 644 645 cell_1rw
* cell instance $23023 m0 *1 71.205,101.01
X$23023 267 588 268 644 645 cell_1rw
* cell instance $23024 r0 *1 71.205,101.01
X$23024 267 589 268 644 645 cell_1rw
* cell instance $23025 m0 *1 71.205,103.74
X$23025 267 590 268 644 645 cell_1rw
* cell instance $23026 r0 *1 71.205,103.74
X$23026 267 591 268 644 645 cell_1rw
* cell instance $23027 m0 *1 71.205,106.47
X$23027 267 593 268 644 645 cell_1rw
* cell instance $23028 r0 *1 71.205,106.47
X$23028 267 592 268 644 645 cell_1rw
* cell instance $23029 m0 *1 71.205,109.2
X$23029 267 594 268 644 645 cell_1rw
* cell instance $23030 m0 *1 71.205,111.93
X$23030 267 597 268 644 645 cell_1rw
* cell instance $23031 r0 *1 71.205,109.2
X$23031 267 595 268 644 645 cell_1rw
* cell instance $23032 r0 *1 71.205,111.93
X$23032 267 596 268 644 645 cell_1rw
* cell instance $23033 m0 *1 71.205,114.66
X$23033 267 598 268 644 645 cell_1rw
* cell instance $23034 r0 *1 71.205,114.66
X$23034 267 599 268 644 645 cell_1rw
* cell instance $23035 m0 *1 71.205,117.39
X$23035 267 600 268 644 645 cell_1rw
* cell instance $23036 r0 *1 71.205,117.39
X$23036 267 601 268 644 645 cell_1rw
* cell instance $23037 m0 *1 71.205,120.12
X$23037 267 602 268 644 645 cell_1rw
* cell instance $23038 r0 *1 71.205,120.12
X$23038 267 603 268 644 645 cell_1rw
* cell instance $23039 m0 *1 71.205,122.85
X$23039 267 604 268 644 645 cell_1rw
* cell instance $23040 r0 *1 71.205,122.85
X$23040 267 605 268 644 645 cell_1rw
* cell instance $23041 m0 *1 71.205,125.58
X$23041 267 606 268 644 645 cell_1rw
* cell instance $23042 r0 *1 71.205,125.58
X$23042 267 607 268 644 645 cell_1rw
* cell instance $23043 m0 *1 71.205,128.31
X$23043 267 609 268 644 645 cell_1rw
* cell instance $23044 r0 *1 71.205,128.31
X$23044 267 608 268 644 645 cell_1rw
* cell instance $23045 m0 *1 71.205,131.04
X$23045 267 610 268 644 645 cell_1rw
* cell instance $23046 r0 *1 71.205,131.04
X$23046 267 611 268 644 645 cell_1rw
* cell instance $23047 m0 *1 71.205,133.77
X$23047 267 612 268 644 645 cell_1rw
* cell instance $23048 r0 *1 71.205,133.77
X$23048 267 613 268 644 645 cell_1rw
* cell instance $23049 m0 *1 71.205,136.5
X$23049 267 615 268 644 645 cell_1rw
* cell instance $23050 r0 *1 71.205,136.5
X$23050 267 614 268 644 645 cell_1rw
* cell instance $23051 m0 *1 71.205,139.23
X$23051 267 617 268 644 645 cell_1rw
* cell instance $23052 r0 *1 71.205,139.23
X$23052 267 616 268 644 645 cell_1rw
* cell instance $23053 m0 *1 71.205,141.96
X$23053 267 618 268 644 645 cell_1rw
* cell instance $23054 r0 *1 71.205,141.96
X$23054 267 619 268 644 645 cell_1rw
* cell instance $23055 m0 *1 71.205,144.69
X$23055 267 620 268 644 645 cell_1rw
* cell instance $23056 r0 *1 71.205,144.69
X$23056 267 621 268 644 645 cell_1rw
* cell instance $23057 m0 *1 71.205,147.42
X$23057 267 622 268 644 645 cell_1rw
* cell instance $23058 r0 *1 71.205,147.42
X$23058 267 623 268 644 645 cell_1rw
* cell instance $23059 m0 *1 71.205,150.15
X$23059 267 624 268 644 645 cell_1rw
* cell instance $23060 r0 *1 71.205,150.15
X$23060 267 625 268 644 645 cell_1rw
* cell instance $23061 m0 *1 71.205,152.88
X$23061 267 626 268 644 645 cell_1rw
* cell instance $23062 r0 *1 71.205,152.88
X$23062 267 627 268 644 645 cell_1rw
* cell instance $23063 m0 *1 71.205,155.61
X$23063 267 628 268 644 645 cell_1rw
* cell instance $23064 r0 *1 71.205,155.61
X$23064 267 629 268 644 645 cell_1rw
* cell instance $23065 m0 *1 71.205,158.34
X$23065 267 630 268 644 645 cell_1rw
* cell instance $23066 m0 *1 71.205,161.07
X$23066 267 632 268 644 645 cell_1rw
* cell instance $23067 r0 *1 71.205,158.34
X$23067 267 631 268 644 645 cell_1rw
* cell instance $23068 r0 *1 71.205,161.07
X$23068 267 633 268 644 645 cell_1rw
* cell instance $23069 m0 *1 71.205,163.8
X$23069 267 634 268 644 645 cell_1rw
* cell instance $23070 r0 *1 71.205,163.8
X$23070 267 635 268 644 645 cell_1rw
* cell instance $23071 m0 *1 71.205,166.53
X$23071 267 637 268 644 645 cell_1rw
* cell instance $23072 r0 *1 71.205,166.53
X$23072 267 636 268 644 645 cell_1rw
* cell instance $23073 m0 *1 71.205,169.26
X$23073 267 639 268 644 645 cell_1rw
* cell instance $23074 r0 *1 71.205,169.26
X$23074 267 638 268 644 645 cell_1rw
* cell instance $23075 m0 *1 71.205,171.99
X$23075 267 640 268 644 645 cell_1rw
* cell instance $23076 r0 *1 71.205,171.99
X$23076 267 641 268 644 645 cell_1rw
* cell instance $23077 m0 *1 71.205,174.72
X$23077 267 642 268 644 645 cell_1rw
* cell instance $23078 r0 *1 71.205,174.72
X$23078 267 643 268 644 645 cell_1rw
* cell instance $23079 r0 *1 71.91,87.36
X$23079 269 322 270 644 645 cell_1rw
* cell instance $23080 m0 *1 71.91,90.09
X$23080 269 581 270 644 645 cell_1rw
* cell instance $23081 m0 *1 71.91,92.82
X$23081 269 583 270 644 645 cell_1rw
* cell instance $23082 r0 *1 71.91,90.09
X$23082 269 580 270 644 645 cell_1rw
* cell instance $23083 r0 *1 71.91,92.82
X$23083 269 582 270 644 645 cell_1rw
* cell instance $23084 m0 *1 71.91,95.55
X$23084 269 584 270 644 645 cell_1rw
* cell instance $23085 m0 *1 71.91,98.28
X$23085 269 586 270 644 645 cell_1rw
* cell instance $23086 r0 *1 71.91,95.55
X$23086 269 585 270 644 645 cell_1rw
* cell instance $23087 m0 *1 71.91,101.01
X$23087 269 588 270 644 645 cell_1rw
* cell instance $23088 r0 *1 71.91,98.28
X$23088 269 587 270 644 645 cell_1rw
* cell instance $23089 r0 *1 71.91,101.01
X$23089 269 589 270 644 645 cell_1rw
* cell instance $23090 m0 *1 71.91,103.74
X$23090 269 590 270 644 645 cell_1rw
* cell instance $23091 m0 *1 71.91,106.47
X$23091 269 593 270 644 645 cell_1rw
* cell instance $23092 r0 *1 71.91,103.74
X$23092 269 591 270 644 645 cell_1rw
* cell instance $23093 r0 *1 71.91,106.47
X$23093 269 592 270 644 645 cell_1rw
* cell instance $23094 m0 *1 71.91,109.2
X$23094 269 594 270 644 645 cell_1rw
* cell instance $23095 r0 *1 71.91,109.2
X$23095 269 595 270 644 645 cell_1rw
* cell instance $23096 m0 *1 71.91,111.93
X$23096 269 597 270 644 645 cell_1rw
* cell instance $23097 r0 *1 71.91,111.93
X$23097 269 596 270 644 645 cell_1rw
* cell instance $23098 m0 *1 71.91,114.66
X$23098 269 598 270 644 645 cell_1rw
* cell instance $23099 r0 *1 71.91,114.66
X$23099 269 599 270 644 645 cell_1rw
* cell instance $23100 m0 *1 71.91,117.39
X$23100 269 600 270 644 645 cell_1rw
* cell instance $23101 r0 *1 71.91,117.39
X$23101 269 601 270 644 645 cell_1rw
* cell instance $23102 m0 *1 71.91,120.12
X$23102 269 602 270 644 645 cell_1rw
* cell instance $23103 r0 *1 71.91,120.12
X$23103 269 603 270 644 645 cell_1rw
* cell instance $23104 m0 *1 71.91,122.85
X$23104 269 604 270 644 645 cell_1rw
* cell instance $23105 r0 *1 71.91,122.85
X$23105 269 605 270 644 645 cell_1rw
* cell instance $23106 m0 *1 71.91,125.58
X$23106 269 606 270 644 645 cell_1rw
* cell instance $23107 m0 *1 71.91,128.31
X$23107 269 609 270 644 645 cell_1rw
* cell instance $23108 r0 *1 71.91,125.58
X$23108 269 607 270 644 645 cell_1rw
* cell instance $23109 r0 *1 71.91,128.31
X$23109 269 608 270 644 645 cell_1rw
* cell instance $23110 m0 *1 71.91,131.04
X$23110 269 610 270 644 645 cell_1rw
* cell instance $23111 m0 *1 71.91,133.77
X$23111 269 612 270 644 645 cell_1rw
* cell instance $23112 r0 *1 71.91,131.04
X$23112 269 611 270 644 645 cell_1rw
* cell instance $23113 r0 *1 71.91,133.77
X$23113 269 613 270 644 645 cell_1rw
* cell instance $23114 m0 *1 71.91,136.5
X$23114 269 615 270 644 645 cell_1rw
* cell instance $23115 r0 *1 71.91,136.5
X$23115 269 614 270 644 645 cell_1rw
* cell instance $23116 m0 *1 71.91,139.23
X$23116 269 617 270 644 645 cell_1rw
* cell instance $23117 r0 *1 71.91,139.23
X$23117 269 616 270 644 645 cell_1rw
* cell instance $23118 m0 *1 71.91,141.96
X$23118 269 618 270 644 645 cell_1rw
* cell instance $23119 r0 *1 71.91,141.96
X$23119 269 619 270 644 645 cell_1rw
* cell instance $23120 m0 *1 71.91,144.69
X$23120 269 620 270 644 645 cell_1rw
* cell instance $23121 r0 *1 71.91,144.69
X$23121 269 621 270 644 645 cell_1rw
* cell instance $23122 m0 *1 71.91,147.42
X$23122 269 622 270 644 645 cell_1rw
* cell instance $23123 m0 *1 71.91,150.15
X$23123 269 624 270 644 645 cell_1rw
* cell instance $23124 r0 *1 71.91,147.42
X$23124 269 623 270 644 645 cell_1rw
* cell instance $23125 m0 *1 71.91,152.88
X$23125 269 626 270 644 645 cell_1rw
* cell instance $23126 r0 *1 71.91,150.15
X$23126 269 625 270 644 645 cell_1rw
* cell instance $23127 r0 *1 71.91,152.88
X$23127 269 627 270 644 645 cell_1rw
* cell instance $23128 m0 *1 71.91,155.61
X$23128 269 628 270 644 645 cell_1rw
* cell instance $23129 r0 *1 71.91,155.61
X$23129 269 629 270 644 645 cell_1rw
* cell instance $23130 m0 *1 71.91,158.34
X$23130 269 630 270 644 645 cell_1rw
* cell instance $23131 r0 *1 71.91,158.34
X$23131 269 631 270 644 645 cell_1rw
* cell instance $23132 m0 *1 71.91,161.07
X$23132 269 632 270 644 645 cell_1rw
* cell instance $23133 m0 *1 71.91,163.8
X$23133 269 634 270 644 645 cell_1rw
* cell instance $23134 r0 *1 71.91,161.07
X$23134 269 633 270 644 645 cell_1rw
* cell instance $23135 m0 *1 71.91,166.53
X$23135 269 637 270 644 645 cell_1rw
* cell instance $23136 r0 *1 71.91,163.8
X$23136 269 635 270 644 645 cell_1rw
* cell instance $23137 r0 *1 71.91,166.53
X$23137 269 636 270 644 645 cell_1rw
* cell instance $23138 m0 *1 71.91,169.26
X$23138 269 639 270 644 645 cell_1rw
* cell instance $23139 m0 *1 71.91,171.99
X$23139 269 640 270 644 645 cell_1rw
* cell instance $23140 r0 *1 71.91,169.26
X$23140 269 638 270 644 645 cell_1rw
* cell instance $23141 m0 *1 71.91,174.72
X$23141 269 642 270 644 645 cell_1rw
* cell instance $23142 r0 *1 71.91,171.99
X$23142 269 641 270 644 645 cell_1rw
* cell instance $23143 r0 *1 71.91,174.72
X$23143 269 643 270 644 645 cell_1rw
* cell instance $23144 m0 *1 72.615,90.09
X$23144 271 581 272 644 645 cell_1rw
* cell instance $23145 r0 *1 72.615,87.36
X$23145 271 322 272 644 645 cell_1rw
* cell instance $23146 r0 *1 72.615,90.09
X$23146 271 580 272 644 645 cell_1rw
* cell instance $23147 m0 *1 72.615,92.82
X$23147 271 583 272 644 645 cell_1rw
* cell instance $23148 r0 *1 72.615,92.82
X$23148 271 582 272 644 645 cell_1rw
* cell instance $23149 m0 *1 72.615,95.55
X$23149 271 584 272 644 645 cell_1rw
* cell instance $23150 r0 *1 72.615,95.55
X$23150 271 585 272 644 645 cell_1rw
* cell instance $23151 m0 *1 72.615,98.28
X$23151 271 586 272 644 645 cell_1rw
* cell instance $23152 r0 *1 72.615,98.28
X$23152 271 587 272 644 645 cell_1rw
* cell instance $23153 m0 *1 72.615,101.01
X$23153 271 588 272 644 645 cell_1rw
* cell instance $23154 r0 *1 72.615,101.01
X$23154 271 589 272 644 645 cell_1rw
* cell instance $23155 m0 *1 72.615,103.74
X$23155 271 590 272 644 645 cell_1rw
* cell instance $23156 r0 *1 72.615,103.74
X$23156 271 591 272 644 645 cell_1rw
* cell instance $23157 m0 *1 72.615,106.47
X$23157 271 593 272 644 645 cell_1rw
* cell instance $23158 r0 *1 72.615,106.47
X$23158 271 592 272 644 645 cell_1rw
* cell instance $23159 m0 *1 72.615,109.2
X$23159 271 594 272 644 645 cell_1rw
* cell instance $23160 r0 *1 72.615,109.2
X$23160 271 595 272 644 645 cell_1rw
* cell instance $23161 m0 *1 72.615,111.93
X$23161 271 597 272 644 645 cell_1rw
* cell instance $23162 r0 *1 72.615,111.93
X$23162 271 596 272 644 645 cell_1rw
* cell instance $23163 m0 *1 72.615,114.66
X$23163 271 598 272 644 645 cell_1rw
* cell instance $23164 r0 *1 72.615,114.66
X$23164 271 599 272 644 645 cell_1rw
* cell instance $23165 m0 *1 72.615,117.39
X$23165 271 600 272 644 645 cell_1rw
* cell instance $23166 r0 *1 72.615,117.39
X$23166 271 601 272 644 645 cell_1rw
* cell instance $23167 m0 *1 72.615,120.12
X$23167 271 602 272 644 645 cell_1rw
* cell instance $23168 r0 *1 72.615,120.12
X$23168 271 603 272 644 645 cell_1rw
* cell instance $23169 m0 *1 72.615,122.85
X$23169 271 604 272 644 645 cell_1rw
* cell instance $23170 r0 *1 72.615,122.85
X$23170 271 605 272 644 645 cell_1rw
* cell instance $23171 m0 *1 72.615,125.58
X$23171 271 606 272 644 645 cell_1rw
* cell instance $23172 r0 *1 72.615,125.58
X$23172 271 607 272 644 645 cell_1rw
* cell instance $23173 m0 *1 72.615,128.31
X$23173 271 609 272 644 645 cell_1rw
* cell instance $23174 r0 *1 72.615,128.31
X$23174 271 608 272 644 645 cell_1rw
* cell instance $23175 m0 *1 72.615,131.04
X$23175 271 610 272 644 645 cell_1rw
* cell instance $23176 r0 *1 72.615,131.04
X$23176 271 611 272 644 645 cell_1rw
* cell instance $23177 m0 *1 72.615,133.77
X$23177 271 612 272 644 645 cell_1rw
* cell instance $23178 r0 *1 72.615,133.77
X$23178 271 613 272 644 645 cell_1rw
* cell instance $23179 m0 *1 72.615,136.5
X$23179 271 615 272 644 645 cell_1rw
* cell instance $23180 r0 *1 72.615,136.5
X$23180 271 614 272 644 645 cell_1rw
* cell instance $23181 m0 *1 72.615,139.23
X$23181 271 617 272 644 645 cell_1rw
* cell instance $23182 m0 *1 72.615,141.96
X$23182 271 618 272 644 645 cell_1rw
* cell instance $23183 r0 *1 72.615,139.23
X$23183 271 616 272 644 645 cell_1rw
* cell instance $23184 r0 *1 72.615,141.96
X$23184 271 619 272 644 645 cell_1rw
* cell instance $23185 m0 *1 72.615,144.69
X$23185 271 620 272 644 645 cell_1rw
* cell instance $23186 r0 *1 72.615,144.69
X$23186 271 621 272 644 645 cell_1rw
* cell instance $23187 m0 *1 72.615,147.42
X$23187 271 622 272 644 645 cell_1rw
* cell instance $23188 r0 *1 72.615,147.42
X$23188 271 623 272 644 645 cell_1rw
* cell instance $23189 m0 *1 72.615,150.15
X$23189 271 624 272 644 645 cell_1rw
* cell instance $23190 r0 *1 72.615,150.15
X$23190 271 625 272 644 645 cell_1rw
* cell instance $23191 m0 *1 72.615,152.88
X$23191 271 626 272 644 645 cell_1rw
* cell instance $23192 r0 *1 72.615,152.88
X$23192 271 627 272 644 645 cell_1rw
* cell instance $23193 m0 *1 72.615,155.61
X$23193 271 628 272 644 645 cell_1rw
* cell instance $23194 r0 *1 72.615,155.61
X$23194 271 629 272 644 645 cell_1rw
* cell instance $23195 m0 *1 72.615,158.34
X$23195 271 630 272 644 645 cell_1rw
* cell instance $23196 r0 *1 72.615,158.34
X$23196 271 631 272 644 645 cell_1rw
* cell instance $23197 m0 *1 72.615,161.07
X$23197 271 632 272 644 645 cell_1rw
* cell instance $23198 m0 *1 72.615,163.8
X$23198 271 634 272 644 645 cell_1rw
* cell instance $23199 r0 *1 72.615,161.07
X$23199 271 633 272 644 645 cell_1rw
* cell instance $23200 r0 *1 72.615,163.8
X$23200 271 635 272 644 645 cell_1rw
* cell instance $23201 m0 *1 72.615,166.53
X$23201 271 637 272 644 645 cell_1rw
* cell instance $23202 r0 *1 72.615,166.53
X$23202 271 636 272 644 645 cell_1rw
* cell instance $23203 m0 *1 72.615,169.26
X$23203 271 639 272 644 645 cell_1rw
* cell instance $23204 r0 *1 72.615,169.26
X$23204 271 638 272 644 645 cell_1rw
* cell instance $23205 m0 *1 72.615,171.99
X$23205 271 640 272 644 645 cell_1rw
* cell instance $23206 m0 *1 72.615,174.72
X$23206 271 642 272 644 645 cell_1rw
* cell instance $23207 r0 *1 72.615,171.99
X$23207 271 641 272 644 645 cell_1rw
* cell instance $23208 r0 *1 72.615,174.72
X$23208 271 643 272 644 645 cell_1rw
* cell instance $23209 r0 *1 73.32,87.36
X$23209 273 322 274 644 645 cell_1rw
* cell instance $23210 m0 *1 73.32,90.09
X$23210 273 581 274 644 645 cell_1rw
* cell instance $23211 r0 *1 73.32,90.09
X$23211 273 580 274 644 645 cell_1rw
* cell instance $23212 m0 *1 73.32,92.82
X$23212 273 583 274 644 645 cell_1rw
* cell instance $23213 r0 *1 73.32,92.82
X$23213 273 582 274 644 645 cell_1rw
* cell instance $23214 m0 *1 73.32,95.55
X$23214 273 584 274 644 645 cell_1rw
* cell instance $23215 r0 *1 73.32,95.55
X$23215 273 585 274 644 645 cell_1rw
* cell instance $23216 m0 *1 73.32,98.28
X$23216 273 586 274 644 645 cell_1rw
* cell instance $23217 r0 *1 73.32,98.28
X$23217 273 587 274 644 645 cell_1rw
* cell instance $23218 m0 *1 73.32,101.01
X$23218 273 588 274 644 645 cell_1rw
* cell instance $23219 r0 *1 73.32,101.01
X$23219 273 589 274 644 645 cell_1rw
* cell instance $23220 m0 *1 73.32,103.74
X$23220 273 590 274 644 645 cell_1rw
* cell instance $23221 r0 *1 73.32,103.74
X$23221 273 591 274 644 645 cell_1rw
* cell instance $23222 m0 *1 73.32,106.47
X$23222 273 593 274 644 645 cell_1rw
* cell instance $23223 r0 *1 73.32,106.47
X$23223 273 592 274 644 645 cell_1rw
* cell instance $23224 m0 *1 73.32,109.2
X$23224 273 594 274 644 645 cell_1rw
* cell instance $23225 r0 *1 73.32,109.2
X$23225 273 595 274 644 645 cell_1rw
* cell instance $23226 m0 *1 73.32,111.93
X$23226 273 597 274 644 645 cell_1rw
* cell instance $23227 r0 *1 73.32,111.93
X$23227 273 596 274 644 645 cell_1rw
* cell instance $23228 m0 *1 73.32,114.66
X$23228 273 598 274 644 645 cell_1rw
* cell instance $23229 m0 *1 73.32,117.39
X$23229 273 600 274 644 645 cell_1rw
* cell instance $23230 r0 *1 73.32,114.66
X$23230 273 599 274 644 645 cell_1rw
* cell instance $23231 r0 *1 73.32,117.39
X$23231 273 601 274 644 645 cell_1rw
* cell instance $23232 m0 *1 73.32,120.12
X$23232 273 602 274 644 645 cell_1rw
* cell instance $23233 r0 *1 73.32,120.12
X$23233 273 603 274 644 645 cell_1rw
* cell instance $23234 m0 *1 73.32,122.85
X$23234 273 604 274 644 645 cell_1rw
* cell instance $23235 r0 *1 73.32,122.85
X$23235 273 605 274 644 645 cell_1rw
* cell instance $23236 m0 *1 73.32,125.58
X$23236 273 606 274 644 645 cell_1rw
* cell instance $23237 r0 *1 73.32,125.58
X$23237 273 607 274 644 645 cell_1rw
* cell instance $23238 m0 *1 73.32,128.31
X$23238 273 609 274 644 645 cell_1rw
* cell instance $23239 m0 *1 73.32,131.04
X$23239 273 610 274 644 645 cell_1rw
* cell instance $23240 r0 *1 73.32,128.31
X$23240 273 608 274 644 645 cell_1rw
* cell instance $23241 r0 *1 73.32,131.04
X$23241 273 611 274 644 645 cell_1rw
* cell instance $23242 m0 *1 73.32,133.77
X$23242 273 612 274 644 645 cell_1rw
* cell instance $23243 r0 *1 73.32,133.77
X$23243 273 613 274 644 645 cell_1rw
* cell instance $23244 m0 *1 73.32,136.5
X$23244 273 615 274 644 645 cell_1rw
* cell instance $23245 m0 *1 73.32,139.23
X$23245 273 617 274 644 645 cell_1rw
* cell instance $23246 r0 *1 73.32,136.5
X$23246 273 614 274 644 645 cell_1rw
* cell instance $23247 r0 *1 73.32,139.23
X$23247 273 616 274 644 645 cell_1rw
* cell instance $23248 m0 *1 73.32,141.96
X$23248 273 618 274 644 645 cell_1rw
* cell instance $23249 r0 *1 73.32,141.96
X$23249 273 619 274 644 645 cell_1rw
* cell instance $23250 m0 *1 73.32,144.69
X$23250 273 620 274 644 645 cell_1rw
* cell instance $23251 m0 *1 73.32,147.42
X$23251 273 622 274 644 645 cell_1rw
* cell instance $23252 r0 *1 73.32,144.69
X$23252 273 621 274 644 645 cell_1rw
* cell instance $23253 r0 *1 73.32,147.42
X$23253 273 623 274 644 645 cell_1rw
* cell instance $23254 m0 *1 73.32,150.15
X$23254 273 624 274 644 645 cell_1rw
* cell instance $23255 r0 *1 73.32,150.15
X$23255 273 625 274 644 645 cell_1rw
* cell instance $23256 m0 *1 73.32,152.88
X$23256 273 626 274 644 645 cell_1rw
* cell instance $23257 r0 *1 73.32,152.88
X$23257 273 627 274 644 645 cell_1rw
* cell instance $23258 m0 *1 73.32,155.61
X$23258 273 628 274 644 645 cell_1rw
* cell instance $23259 r0 *1 73.32,155.61
X$23259 273 629 274 644 645 cell_1rw
* cell instance $23260 m0 *1 73.32,158.34
X$23260 273 630 274 644 645 cell_1rw
* cell instance $23261 r0 *1 73.32,158.34
X$23261 273 631 274 644 645 cell_1rw
* cell instance $23262 m0 *1 73.32,161.07
X$23262 273 632 274 644 645 cell_1rw
* cell instance $23263 m0 *1 73.32,163.8
X$23263 273 634 274 644 645 cell_1rw
* cell instance $23264 r0 *1 73.32,161.07
X$23264 273 633 274 644 645 cell_1rw
* cell instance $23265 r0 *1 73.32,163.8
X$23265 273 635 274 644 645 cell_1rw
* cell instance $23266 m0 *1 73.32,166.53
X$23266 273 637 274 644 645 cell_1rw
* cell instance $23267 r0 *1 73.32,166.53
X$23267 273 636 274 644 645 cell_1rw
* cell instance $23268 m0 *1 73.32,169.26
X$23268 273 639 274 644 645 cell_1rw
* cell instance $23269 r0 *1 73.32,169.26
X$23269 273 638 274 644 645 cell_1rw
* cell instance $23270 m0 *1 73.32,171.99
X$23270 273 640 274 644 645 cell_1rw
* cell instance $23271 r0 *1 73.32,171.99
X$23271 273 641 274 644 645 cell_1rw
* cell instance $23272 m0 *1 73.32,174.72
X$23272 273 642 274 644 645 cell_1rw
* cell instance $23273 r0 *1 73.32,174.72
X$23273 273 643 274 644 645 cell_1rw
* cell instance $23274 r0 *1 74.025,87.36
X$23274 275 322 276 644 645 cell_1rw
* cell instance $23275 m0 *1 74.025,90.09
X$23275 275 581 276 644 645 cell_1rw
* cell instance $23276 r0 *1 74.025,90.09
X$23276 275 580 276 644 645 cell_1rw
* cell instance $23277 m0 *1 74.025,92.82
X$23277 275 583 276 644 645 cell_1rw
* cell instance $23278 r0 *1 74.025,92.82
X$23278 275 582 276 644 645 cell_1rw
* cell instance $23279 m0 *1 74.025,95.55
X$23279 275 584 276 644 645 cell_1rw
* cell instance $23280 r0 *1 74.025,95.55
X$23280 275 585 276 644 645 cell_1rw
* cell instance $23281 m0 *1 74.025,98.28
X$23281 275 586 276 644 645 cell_1rw
* cell instance $23282 r0 *1 74.025,98.28
X$23282 275 587 276 644 645 cell_1rw
* cell instance $23283 m0 *1 74.025,101.01
X$23283 275 588 276 644 645 cell_1rw
* cell instance $23284 r0 *1 74.025,101.01
X$23284 275 589 276 644 645 cell_1rw
* cell instance $23285 m0 *1 74.025,103.74
X$23285 275 590 276 644 645 cell_1rw
* cell instance $23286 r0 *1 74.025,103.74
X$23286 275 591 276 644 645 cell_1rw
* cell instance $23287 m0 *1 74.025,106.47
X$23287 275 593 276 644 645 cell_1rw
* cell instance $23288 r0 *1 74.025,106.47
X$23288 275 592 276 644 645 cell_1rw
* cell instance $23289 m0 *1 74.025,109.2
X$23289 275 594 276 644 645 cell_1rw
* cell instance $23290 r0 *1 74.025,109.2
X$23290 275 595 276 644 645 cell_1rw
* cell instance $23291 m0 *1 74.025,111.93
X$23291 275 597 276 644 645 cell_1rw
* cell instance $23292 r0 *1 74.025,111.93
X$23292 275 596 276 644 645 cell_1rw
* cell instance $23293 m0 *1 74.025,114.66
X$23293 275 598 276 644 645 cell_1rw
* cell instance $23294 r0 *1 74.025,114.66
X$23294 275 599 276 644 645 cell_1rw
* cell instance $23295 m0 *1 74.025,117.39
X$23295 275 600 276 644 645 cell_1rw
* cell instance $23296 r0 *1 74.025,117.39
X$23296 275 601 276 644 645 cell_1rw
* cell instance $23297 m0 *1 74.025,120.12
X$23297 275 602 276 644 645 cell_1rw
* cell instance $23298 r0 *1 74.025,120.12
X$23298 275 603 276 644 645 cell_1rw
* cell instance $23299 m0 *1 74.025,122.85
X$23299 275 604 276 644 645 cell_1rw
* cell instance $23300 r0 *1 74.025,122.85
X$23300 275 605 276 644 645 cell_1rw
* cell instance $23301 m0 *1 74.025,125.58
X$23301 275 606 276 644 645 cell_1rw
* cell instance $23302 m0 *1 74.025,128.31
X$23302 275 609 276 644 645 cell_1rw
* cell instance $23303 r0 *1 74.025,125.58
X$23303 275 607 276 644 645 cell_1rw
* cell instance $23304 r0 *1 74.025,128.31
X$23304 275 608 276 644 645 cell_1rw
* cell instance $23305 m0 *1 74.025,131.04
X$23305 275 610 276 644 645 cell_1rw
* cell instance $23306 r0 *1 74.025,131.04
X$23306 275 611 276 644 645 cell_1rw
* cell instance $23307 m0 *1 74.025,133.77
X$23307 275 612 276 644 645 cell_1rw
* cell instance $23308 r0 *1 74.025,133.77
X$23308 275 613 276 644 645 cell_1rw
* cell instance $23309 m0 *1 74.025,136.5
X$23309 275 615 276 644 645 cell_1rw
* cell instance $23310 m0 *1 74.025,139.23
X$23310 275 617 276 644 645 cell_1rw
* cell instance $23311 r0 *1 74.025,136.5
X$23311 275 614 276 644 645 cell_1rw
* cell instance $23312 r0 *1 74.025,139.23
X$23312 275 616 276 644 645 cell_1rw
* cell instance $23313 m0 *1 74.025,141.96
X$23313 275 618 276 644 645 cell_1rw
* cell instance $23314 r0 *1 74.025,141.96
X$23314 275 619 276 644 645 cell_1rw
* cell instance $23315 m0 *1 74.025,144.69
X$23315 275 620 276 644 645 cell_1rw
* cell instance $23316 r0 *1 74.025,144.69
X$23316 275 621 276 644 645 cell_1rw
* cell instance $23317 m0 *1 74.025,147.42
X$23317 275 622 276 644 645 cell_1rw
* cell instance $23318 r0 *1 74.025,147.42
X$23318 275 623 276 644 645 cell_1rw
* cell instance $23319 m0 *1 74.025,150.15
X$23319 275 624 276 644 645 cell_1rw
* cell instance $23320 r0 *1 74.025,150.15
X$23320 275 625 276 644 645 cell_1rw
* cell instance $23321 m0 *1 74.025,152.88
X$23321 275 626 276 644 645 cell_1rw
* cell instance $23322 r0 *1 74.025,152.88
X$23322 275 627 276 644 645 cell_1rw
* cell instance $23323 m0 *1 74.025,155.61
X$23323 275 628 276 644 645 cell_1rw
* cell instance $23324 r0 *1 74.025,155.61
X$23324 275 629 276 644 645 cell_1rw
* cell instance $23325 m0 *1 74.025,158.34
X$23325 275 630 276 644 645 cell_1rw
* cell instance $23326 r0 *1 74.025,158.34
X$23326 275 631 276 644 645 cell_1rw
* cell instance $23327 m0 *1 74.025,161.07
X$23327 275 632 276 644 645 cell_1rw
* cell instance $23328 r0 *1 74.025,161.07
X$23328 275 633 276 644 645 cell_1rw
* cell instance $23329 m0 *1 74.025,163.8
X$23329 275 634 276 644 645 cell_1rw
* cell instance $23330 r0 *1 74.025,163.8
X$23330 275 635 276 644 645 cell_1rw
* cell instance $23331 m0 *1 74.025,166.53
X$23331 275 637 276 644 645 cell_1rw
* cell instance $23332 r0 *1 74.025,166.53
X$23332 275 636 276 644 645 cell_1rw
* cell instance $23333 m0 *1 74.025,169.26
X$23333 275 639 276 644 645 cell_1rw
* cell instance $23334 r0 *1 74.025,169.26
X$23334 275 638 276 644 645 cell_1rw
* cell instance $23335 m0 *1 74.025,171.99
X$23335 275 640 276 644 645 cell_1rw
* cell instance $23336 r0 *1 74.025,171.99
X$23336 275 641 276 644 645 cell_1rw
* cell instance $23337 m0 *1 74.025,174.72
X$23337 275 642 276 644 645 cell_1rw
* cell instance $23338 r0 *1 74.025,174.72
X$23338 275 643 276 644 645 cell_1rw
* cell instance $23339 r0 *1 74.73,87.36
X$23339 277 322 278 644 645 cell_1rw
* cell instance $23340 m0 *1 74.73,90.09
X$23340 277 581 278 644 645 cell_1rw
* cell instance $23341 r0 *1 74.73,90.09
X$23341 277 580 278 644 645 cell_1rw
* cell instance $23342 m0 *1 74.73,92.82
X$23342 277 583 278 644 645 cell_1rw
* cell instance $23343 m0 *1 74.73,95.55
X$23343 277 584 278 644 645 cell_1rw
* cell instance $23344 r0 *1 74.73,92.82
X$23344 277 582 278 644 645 cell_1rw
* cell instance $23345 m0 *1 74.73,98.28
X$23345 277 586 278 644 645 cell_1rw
* cell instance $23346 r0 *1 74.73,95.55
X$23346 277 585 278 644 645 cell_1rw
* cell instance $23347 r0 *1 74.73,98.28
X$23347 277 587 278 644 645 cell_1rw
* cell instance $23348 m0 *1 74.73,101.01
X$23348 277 588 278 644 645 cell_1rw
* cell instance $23349 r0 *1 74.73,101.01
X$23349 277 589 278 644 645 cell_1rw
* cell instance $23350 m0 *1 74.73,103.74
X$23350 277 590 278 644 645 cell_1rw
* cell instance $23351 r0 *1 74.73,103.74
X$23351 277 591 278 644 645 cell_1rw
* cell instance $23352 m0 *1 74.73,106.47
X$23352 277 593 278 644 645 cell_1rw
* cell instance $23353 r0 *1 74.73,106.47
X$23353 277 592 278 644 645 cell_1rw
* cell instance $23354 m0 *1 74.73,109.2
X$23354 277 594 278 644 645 cell_1rw
* cell instance $23355 r0 *1 74.73,109.2
X$23355 277 595 278 644 645 cell_1rw
* cell instance $23356 m0 *1 74.73,111.93
X$23356 277 597 278 644 645 cell_1rw
* cell instance $23357 r0 *1 74.73,111.93
X$23357 277 596 278 644 645 cell_1rw
* cell instance $23358 m0 *1 74.73,114.66
X$23358 277 598 278 644 645 cell_1rw
* cell instance $23359 r0 *1 74.73,114.66
X$23359 277 599 278 644 645 cell_1rw
* cell instance $23360 m0 *1 74.73,117.39
X$23360 277 600 278 644 645 cell_1rw
* cell instance $23361 r0 *1 74.73,117.39
X$23361 277 601 278 644 645 cell_1rw
* cell instance $23362 m0 *1 74.73,120.12
X$23362 277 602 278 644 645 cell_1rw
* cell instance $23363 r0 *1 74.73,120.12
X$23363 277 603 278 644 645 cell_1rw
* cell instance $23364 m0 *1 74.73,122.85
X$23364 277 604 278 644 645 cell_1rw
* cell instance $23365 m0 *1 74.73,125.58
X$23365 277 606 278 644 645 cell_1rw
* cell instance $23366 r0 *1 74.73,122.85
X$23366 277 605 278 644 645 cell_1rw
* cell instance $23367 r0 *1 74.73,125.58
X$23367 277 607 278 644 645 cell_1rw
* cell instance $23368 m0 *1 74.73,128.31
X$23368 277 609 278 644 645 cell_1rw
* cell instance $23369 r0 *1 74.73,128.31
X$23369 277 608 278 644 645 cell_1rw
* cell instance $23370 m0 *1 74.73,131.04
X$23370 277 610 278 644 645 cell_1rw
* cell instance $23371 r0 *1 74.73,131.04
X$23371 277 611 278 644 645 cell_1rw
* cell instance $23372 m0 *1 74.73,133.77
X$23372 277 612 278 644 645 cell_1rw
* cell instance $23373 r0 *1 74.73,133.77
X$23373 277 613 278 644 645 cell_1rw
* cell instance $23374 m0 *1 74.73,136.5
X$23374 277 615 278 644 645 cell_1rw
* cell instance $23375 r0 *1 74.73,136.5
X$23375 277 614 278 644 645 cell_1rw
* cell instance $23376 m0 *1 74.73,139.23
X$23376 277 617 278 644 645 cell_1rw
* cell instance $23377 m0 *1 74.73,141.96
X$23377 277 618 278 644 645 cell_1rw
* cell instance $23378 r0 *1 74.73,139.23
X$23378 277 616 278 644 645 cell_1rw
* cell instance $23379 r0 *1 74.73,141.96
X$23379 277 619 278 644 645 cell_1rw
* cell instance $23380 m0 *1 74.73,144.69
X$23380 277 620 278 644 645 cell_1rw
* cell instance $23381 r0 *1 74.73,144.69
X$23381 277 621 278 644 645 cell_1rw
* cell instance $23382 m0 *1 74.73,147.42
X$23382 277 622 278 644 645 cell_1rw
* cell instance $23383 r0 *1 74.73,147.42
X$23383 277 623 278 644 645 cell_1rw
* cell instance $23384 m0 *1 74.73,150.15
X$23384 277 624 278 644 645 cell_1rw
* cell instance $23385 r0 *1 74.73,150.15
X$23385 277 625 278 644 645 cell_1rw
* cell instance $23386 m0 *1 74.73,152.88
X$23386 277 626 278 644 645 cell_1rw
* cell instance $23387 r0 *1 74.73,152.88
X$23387 277 627 278 644 645 cell_1rw
* cell instance $23388 m0 *1 74.73,155.61
X$23388 277 628 278 644 645 cell_1rw
* cell instance $23389 r0 *1 74.73,155.61
X$23389 277 629 278 644 645 cell_1rw
* cell instance $23390 m0 *1 74.73,158.34
X$23390 277 630 278 644 645 cell_1rw
* cell instance $23391 m0 *1 74.73,161.07
X$23391 277 632 278 644 645 cell_1rw
* cell instance $23392 r0 *1 74.73,158.34
X$23392 277 631 278 644 645 cell_1rw
* cell instance $23393 r0 *1 74.73,161.07
X$23393 277 633 278 644 645 cell_1rw
* cell instance $23394 m0 *1 74.73,163.8
X$23394 277 634 278 644 645 cell_1rw
* cell instance $23395 r0 *1 74.73,163.8
X$23395 277 635 278 644 645 cell_1rw
* cell instance $23396 m0 *1 74.73,166.53
X$23396 277 637 278 644 645 cell_1rw
* cell instance $23397 m0 *1 74.73,169.26
X$23397 277 639 278 644 645 cell_1rw
* cell instance $23398 r0 *1 74.73,166.53
X$23398 277 636 278 644 645 cell_1rw
* cell instance $23399 r0 *1 74.73,169.26
X$23399 277 638 278 644 645 cell_1rw
* cell instance $23400 m0 *1 74.73,171.99
X$23400 277 640 278 644 645 cell_1rw
* cell instance $23401 r0 *1 74.73,171.99
X$23401 277 641 278 644 645 cell_1rw
* cell instance $23402 m0 *1 74.73,174.72
X$23402 277 642 278 644 645 cell_1rw
* cell instance $23403 r0 *1 74.73,174.72
X$23403 277 643 278 644 645 cell_1rw
* cell instance $23404 r0 *1 75.435,87.36
X$23404 279 322 280 644 645 cell_1rw
* cell instance $23405 m0 *1 75.435,90.09
X$23405 279 581 280 644 645 cell_1rw
* cell instance $23406 m0 *1 75.435,92.82
X$23406 279 583 280 644 645 cell_1rw
* cell instance $23407 r0 *1 75.435,90.09
X$23407 279 580 280 644 645 cell_1rw
* cell instance $23408 m0 *1 75.435,95.55
X$23408 279 584 280 644 645 cell_1rw
* cell instance $23409 r0 *1 75.435,92.82
X$23409 279 582 280 644 645 cell_1rw
* cell instance $23410 m0 *1 75.435,98.28
X$23410 279 586 280 644 645 cell_1rw
* cell instance $23411 r0 *1 75.435,95.55
X$23411 279 585 280 644 645 cell_1rw
* cell instance $23412 r0 *1 75.435,98.28
X$23412 279 587 280 644 645 cell_1rw
* cell instance $23413 m0 *1 75.435,101.01
X$23413 279 588 280 644 645 cell_1rw
* cell instance $23414 r0 *1 75.435,101.01
X$23414 279 589 280 644 645 cell_1rw
* cell instance $23415 m0 *1 75.435,103.74
X$23415 279 590 280 644 645 cell_1rw
* cell instance $23416 m0 *1 75.435,106.47
X$23416 279 593 280 644 645 cell_1rw
* cell instance $23417 r0 *1 75.435,103.74
X$23417 279 591 280 644 645 cell_1rw
* cell instance $23418 r0 *1 75.435,106.47
X$23418 279 592 280 644 645 cell_1rw
* cell instance $23419 m0 *1 75.435,109.2
X$23419 279 594 280 644 645 cell_1rw
* cell instance $23420 r0 *1 75.435,109.2
X$23420 279 595 280 644 645 cell_1rw
* cell instance $23421 m0 *1 75.435,111.93
X$23421 279 597 280 644 645 cell_1rw
* cell instance $23422 r0 *1 75.435,111.93
X$23422 279 596 280 644 645 cell_1rw
* cell instance $23423 m0 *1 75.435,114.66
X$23423 279 598 280 644 645 cell_1rw
* cell instance $23424 r0 *1 75.435,114.66
X$23424 279 599 280 644 645 cell_1rw
* cell instance $23425 m0 *1 75.435,117.39
X$23425 279 600 280 644 645 cell_1rw
* cell instance $23426 r0 *1 75.435,117.39
X$23426 279 601 280 644 645 cell_1rw
* cell instance $23427 m0 *1 75.435,120.12
X$23427 279 602 280 644 645 cell_1rw
* cell instance $23428 r0 *1 75.435,120.12
X$23428 279 603 280 644 645 cell_1rw
* cell instance $23429 m0 *1 75.435,122.85
X$23429 279 604 280 644 645 cell_1rw
* cell instance $23430 r0 *1 75.435,122.85
X$23430 279 605 280 644 645 cell_1rw
* cell instance $23431 m0 *1 75.435,125.58
X$23431 279 606 280 644 645 cell_1rw
* cell instance $23432 m0 *1 75.435,128.31
X$23432 279 609 280 644 645 cell_1rw
* cell instance $23433 r0 *1 75.435,125.58
X$23433 279 607 280 644 645 cell_1rw
* cell instance $23434 r0 *1 75.435,128.31
X$23434 279 608 280 644 645 cell_1rw
* cell instance $23435 m0 *1 75.435,131.04
X$23435 279 610 280 644 645 cell_1rw
* cell instance $23436 r0 *1 75.435,131.04
X$23436 279 611 280 644 645 cell_1rw
* cell instance $23437 m0 *1 75.435,133.77
X$23437 279 612 280 644 645 cell_1rw
* cell instance $23438 r0 *1 75.435,133.77
X$23438 279 613 280 644 645 cell_1rw
* cell instance $23439 m0 *1 75.435,136.5
X$23439 279 615 280 644 645 cell_1rw
* cell instance $23440 r0 *1 75.435,136.5
X$23440 279 614 280 644 645 cell_1rw
* cell instance $23441 m0 *1 75.435,139.23
X$23441 279 617 280 644 645 cell_1rw
* cell instance $23442 m0 *1 75.435,141.96
X$23442 279 618 280 644 645 cell_1rw
* cell instance $23443 r0 *1 75.435,139.23
X$23443 279 616 280 644 645 cell_1rw
* cell instance $23444 r0 *1 75.435,141.96
X$23444 279 619 280 644 645 cell_1rw
* cell instance $23445 m0 *1 75.435,144.69
X$23445 279 620 280 644 645 cell_1rw
* cell instance $23446 m0 *1 75.435,147.42
X$23446 279 622 280 644 645 cell_1rw
* cell instance $23447 r0 *1 75.435,144.69
X$23447 279 621 280 644 645 cell_1rw
* cell instance $23448 r0 *1 75.435,147.42
X$23448 279 623 280 644 645 cell_1rw
* cell instance $23449 m0 *1 75.435,150.15
X$23449 279 624 280 644 645 cell_1rw
* cell instance $23450 r0 *1 75.435,150.15
X$23450 279 625 280 644 645 cell_1rw
* cell instance $23451 m0 *1 75.435,152.88
X$23451 279 626 280 644 645 cell_1rw
* cell instance $23452 r0 *1 75.435,152.88
X$23452 279 627 280 644 645 cell_1rw
* cell instance $23453 m0 *1 75.435,155.61
X$23453 279 628 280 644 645 cell_1rw
* cell instance $23454 r0 *1 75.435,155.61
X$23454 279 629 280 644 645 cell_1rw
* cell instance $23455 m0 *1 75.435,158.34
X$23455 279 630 280 644 645 cell_1rw
* cell instance $23456 r0 *1 75.435,158.34
X$23456 279 631 280 644 645 cell_1rw
* cell instance $23457 m0 *1 75.435,161.07
X$23457 279 632 280 644 645 cell_1rw
* cell instance $23458 r0 *1 75.435,161.07
X$23458 279 633 280 644 645 cell_1rw
* cell instance $23459 m0 *1 75.435,163.8
X$23459 279 634 280 644 645 cell_1rw
* cell instance $23460 r0 *1 75.435,163.8
X$23460 279 635 280 644 645 cell_1rw
* cell instance $23461 m0 *1 75.435,166.53
X$23461 279 637 280 644 645 cell_1rw
* cell instance $23462 r0 *1 75.435,166.53
X$23462 279 636 280 644 645 cell_1rw
* cell instance $23463 m0 *1 75.435,169.26
X$23463 279 639 280 644 645 cell_1rw
* cell instance $23464 m0 *1 75.435,171.99
X$23464 279 640 280 644 645 cell_1rw
* cell instance $23465 r0 *1 75.435,169.26
X$23465 279 638 280 644 645 cell_1rw
* cell instance $23466 r0 *1 75.435,171.99
X$23466 279 641 280 644 645 cell_1rw
* cell instance $23467 m0 *1 75.435,174.72
X$23467 279 642 280 644 645 cell_1rw
* cell instance $23468 r0 *1 75.435,174.72
X$23468 279 643 280 644 645 cell_1rw
* cell instance $23469 r0 *1 76.14,87.36
X$23469 281 322 282 644 645 cell_1rw
* cell instance $23470 m0 *1 76.14,90.09
X$23470 281 581 282 644 645 cell_1rw
* cell instance $23471 r0 *1 76.14,90.09
X$23471 281 580 282 644 645 cell_1rw
* cell instance $23472 m0 *1 76.14,92.82
X$23472 281 583 282 644 645 cell_1rw
* cell instance $23473 r0 *1 76.14,92.82
X$23473 281 582 282 644 645 cell_1rw
* cell instance $23474 m0 *1 76.14,95.55
X$23474 281 584 282 644 645 cell_1rw
* cell instance $23475 r0 *1 76.14,95.55
X$23475 281 585 282 644 645 cell_1rw
* cell instance $23476 m0 *1 76.14,98.28
X$23476 281 586 282 644 645 cell_1rw
* cell instance $23477 r0 *1 76.14,98.28
X$23477 281 587 282 644 645 cell_1rw
* cell instance $23478 m0 *1 76.14,101.01
X$23478 281 588 282 644 645 cell_1rw
* cell instance $23479 r0 *1 76.14,101.01
X$23479 281 589 282 644 645 cell_1rw
* cell instance $23480 m0 *1 76.14,103.74
X$23480 281 590 282 644 645 cell_1rw
* cell instance $23481 m0 *1 76.14,106.47
X$23481 281 593 282 644 645 cell_1rw
* cell instance $23482 r0 *1 76.14,103.74
X$23482 281 591 282 644 645 cell_1rw
* cell instance $23483 r0 *1 76.14,106.47
X$23483 281 592 282 644 645 cell_1rw
* cell instance $23484 m0 *1 76.14,109.2
X$23484 281 594 282 644 645 cell_1rw
* cell instance $23485 m0 *1 76.14,111.93
X$23485 281 597 282 644 645 cell_1rw
* cell instance $23486 r0 *1 76.14,109.2
X$23486 281 595 282 644 645 cell_1rw
* cell instance $23487 r0 *1 76.14,111.93
X$23487 281 596 282 644 645 cell_1rw
* cell instance $23488 m0 *1 76.14,114.66
X$23488 281 598 282 644 645 cell_1rw
* cell instance $23489 r0 *1 76.14,114.66
X$23489 281 599 282 644 645 cell_1rw
* cell instance $23490 m0 *1 76.14,117.39
X$23490 281 600 282 644 645 cell_1rw
* cell instance $23491 m0 *1 76.14,120.12
X$23491 281 602 282 644 645 cell_1rw
* cell instance $23492 r0 *1 76.14,117.39
X$23492 281 601 282 644 645 cell_1rw
* cell instance $23493 r0 *1 76.14,120.12
X$23493 281 603 282 644 645 cell_1rw
* cell instance $23494 m0 *1 76.14,122.85
X$23494 281 604 282 644 645 cell_1rw
* cell instance $23495 r0 *1 76.14,122.85
X$23495 281 605 282 644 645 cell_1rw
* cell instance $23496 m0 *1 76.14,125.58
X$23496 281 606 282 644 645 cell_1rw
* cell instance $23497 r0 *1 76.14,125.58
X$23497 281 607 282 644 645 cell_1rw
* cell instance $23498 m0 *1 76.14,128.31
X$23498 281 609 282 644 645 cell_1rw
* cell instance $23499 r0 *1 76.14,128.31
X$23499 281 608 282 644 645 cell_1rw
* cell instance $23500 m0 *1 76.14,131.04
X$23500 281 610 282 644 645 cell_1rw
* cell instance $23501 r0 *1 76.14,131.04
X$23501 281 611 282 644 645 cell_1rw
* cell instance $23502 m0 *1 76.14,133.77
X$23502 281 612 282 644 645 cell_1rw
* cell instance $23503 r0 *1 76.14,133.77
X$23503 281 613 282 644 645 cell_1rw
* cell instance $23504 m0 *1 76.14,136.5
X$23504 281 615 282 644 645 cell_1rw
* cell instance $23505 r0 *1 76.14,136.5
X$23505 281 614 282 644 645 cell_1rw
* cell instance $23506 m0 *1 76.14,139.23
X$23506 281 617 282 644 645 cell_1rw
* cell instance $23507 m0 *1 76.14,141.96
X$23507 281 618 282 644 645 cell_1rw
* cell instance $23508 r0 *1 76.14,139.23
X$23508 281 616 282 644 645 cell_1rw
* cell instance $23509 r0 *1 76.14,141.96
X$23509 281 619 282 644 645 cell_1rw
* cell instance $23510 m0 *1 76.14,144.69
X$23510 281 620 282 644 645 cell_1rw
* cell instance $23511 r0 *1 76.14,144.69
X$23511 281 621 282 644 645 cell_1rw
* cell instance $23512 m0 *1 76.14,147.42
X$23512 281 622 282 644 645 cell_1rw
* cell instance $23513 r0 *1 76.14,147.42
X$23513 281 623 282 644 645 cell_1rw
* cell instance $23514 m0 *1 76.14,150.15
X$23514 281 624 282 644 645 cell_1rw
* cell instance $23515 r0 *1 76.14,150.15
X$23515 281 625 282 644 645 cell_1rw
* cell instance $23516 m0 *1 76.14,152.88
X$23516 281 626 282 644 645 cell_1rw
* cell instance $23517 r0 *1 76.14,152.88
X$23517 281 627 282 644 645 cell_1rw
* cell instance $23518 m0 *1 76.14,155.61
X$23518 281 628 282 644 645 cell_1rw
* cell instance $23519 r0 *1 76.14,155.61
X$23519 281 629 282 644 645 cell_1rw
* cell instance $23520 m0 *1 76.14,158.34
X$23520 281 630 282 644 645 cell_1rw
* cell instance $23521 r0 *1 76.14,158.34
X$23521 281 631 282 644 645 cell_1rw
* cell instance $23522 m0 *1 76.14,161.07
X$23522 281 632 282 644 645 cell_1rw
* cell instance $23523 r0 *1 76.14,161.07
X$23523 281 633 282 644 645 cell_1rw
* cell instance $23524 m0 *1 76.14,163.8
X$23524 281 634 282 644 645 cell_1rw
* cell instance $23525 m0 *1 76.14,166.53
X$23525 281 637 282 644 645 cell_1rw
* cell instance $23526 r0 *1 76.14,163.8
X$23526 281 635 282 644 645 cell_1rw
* cell instance $23527 r0 *1 76.14,166.53
X$23527 281 636 282 644 645 cell_1rw
* cell instance $23528 m0 *1 76.14,169.26
X$23528 281 639 282 644 645 cell_1rw
* cell instance $23529 r0 *1 76.14,169.26
X$23529 281 638 282 644 645 cell_1rw
* cell instance $23530 m0 *1 76.14,171.99
X$23530 281 640 282 644 645 cell_1rw
* cell instance $23531 r0 *1 76.14,171.99
X$23531 281 641 282 644 645 cell_1rw
* cell instance $23532 m0 *1 76.14,174.72
X$23532 281 642 282 644 645 cell_1rw
* cell instance $23533 r0 *1 76.14,174.72
X$23533 281 643 282 644 645 cell_1rw
* cell instance $23534 m0 *1 76.845,90.09
X$23534 283 581 284 644 645 cell_1rw
* cell instance $23535 r0 *1 76.845,87.36
X$23535 283 322 284 644 645 cell_1rw
* cell instance $23536 r0 *1 76.845,90.09
X$23536 283 580 284 644 645 cell_1rw
* cell instance $23537 m0 *1 76.845,92.82
X$23537 283 583 284 644 645 cell_1rw
* cell instance $23538 m0 *1 76.845,95.55
X$23538 283 584 284 644 645 cell_1rw
* cell instance $23539 r0 *1 76.845,92.82
X$23539 283 582 284 644 645 cell_1rw
* cell instance $23540 r0 *1 76.845,95.55
X$23540 283 585 284 644 645 cell_1rw
* cell instance $23541 m0 *1 76.845,98.28
X$23541 283 586 284 644 645 cell_1rw
* cell instance $23542 r0 *1 76.845,98.28
X$23542 283 587 284 644 645 cell_1rw
* cell instance $23543 m0 *1 76.845,101.01
X$23543 283 588 284 644 645 cell_1rw
* cell instance $23544 r0 *1 76.845,101.01
X$23544 283 589 284 644 645 cell_1rw
* cell instance $23545 m0 *1 76.845,103.74
X$23545 283 590 284 644 645 cell_1rw
* cell instance $23546 r0 *1 76.845,103.74
X$23546 283 591 284 644 645 cell_1rw
* cell instance $23547 m0 *1 76.845,106.47
X$23547 283 593 284 644 645 cell_1rw
* cell instance $23548 m0 *1 76.845,109.2
X$23548 283 594 284 644 645 cell_1rw
* cell instance $23549 r0 *1 76.845,106.47
X$23549 283 592 284 644 645 cell_1rw
* cell instance $23550 m0 *1 76.845,111.93
X$23550 283 597 284 644 645 cell_1rw
* cell instance $23551 r0 *1 76.845,109.2
X$23551 283 595 284 644 645 cell_1rw
* cell instance $23552 r0 *1 76.845,111.93
X$23552 283 596 284 644 645 cell_1rw
* cell instance $23553 m0 *1 76.845,114.66
X$23553 283 598 284 644 645 cell_1rw
* cell instance $23554 m0 *1 76.845,117.39
X$23554 283 600 284 644 645 cell_1rw
* cell instance $23555 r0 *1 76.845,114.66
X$23555 283 599 284 644 645 cell_1rw
* cell instance $23556 r0 *1 76.845,117.39
X$23556 283 601 284 644 645 cell_1rw
* cell instance $23557 m0 *1 76.845,120.12
X$23557 283 602 284 644 645 cell_1rw
* cell instance $23558 r0 *1 76.845,120.12
X$23558 283 603 284 644 645 cell_1rw
* cell instance $23559 m0 *1 76.845,122.85
X$23559 283 604 284 644 645 cell_1rw
* cell instance $23560 r0 *1 76.845,122.85
X$23560 283 605 284 644 645 cell_1rw
* cell instance $23561 m0 *1 76.845,125.58
X$23561 283 606 284 644 645 cell_1rw
* cell instance $23562 r0 *1 76.845,125.58
X$23562 283 607 284 644 645 cell_1rw
* cell instance $23563 m0 *1 76.845,128.31
X$23563 283 609 284 644 645 cell_1rw
* cell instance $23564 r0 *1 76.845,128.31
X$23564 283 608 284 644 645 cell_1rw
* cell instance $23565 m0 *1 76.845,131.04
X$23565 283 610 284 644 645 cell_1rw
* cell instance $23566 r0 *1 76.845,131.04
X$23566 283 611 284 644 645 cell_1rw
* cell instance $23567 m0 *1 76.845,133.77
X$23567 283 612 284 644 645 cell_1rw
* cell instance $23568 m0 *1 76.845,136.5
X$23568 283 615 284 644 645 cell_1rw
* cell instance $23569 r0 *1 76.845,133.77
X$23569 283 613 284 644 645 cell_1rw
* cell instance $23570 r0 *1 76.845,136.5
X$23570 283 614 284 644 645 cell_1rw
* cell instance $23571 m0 *1 76.845,139.23
X$23571 283 617 284 644 645 cell_1rw
* cell instance $23572 r0 *1 76.845,139.23
X$23572 283 616 284 644 645 cell_1rw
* cell instance $23573 m0 *1 76.845,141.96
X$23573 283 618 284 644 645 cell_1rw
* cell instance $23574 r0 *1 76.845,141.96
X$23574 283 619 284 644 645 cell_1rw
* cell instance $23575 m0 *1 76.845,144.69
X$23575 283 620 284 644 645 cell_1rw
* cell instance $23576 r0 *1 76.845,144.69
X$23576 283 621 284 644 645 cell_1rw
* cell instance $23577 m0 *1 76.845,147.42
X$23577 283 622 284 644 645 cell_1rw
* cell instance $23578 m0 *1 76.845,150.15
X$23578 283 624 284 644 645 cell_1rw
* cell instance $23579 r0 *1 76.845,147.42
X$23579 283 623 284 644 645 cell_1rw
* cell instance $23580 r0 *1 76.845,150.15
X$23580 283 625 284 644 645 cell_1rw
* cell instance $23581 m0 *1 76.845,152.88
X$23581 283 626 284 644 645 cell_1rw
* cell instance $23582 r0 *1 76.845,152.88
X$23582 283 627 284 644 645 cell_1rw
* cell instance $23583 m0 *1 76.845,155.61
X$23583 283 628 284 644 645 cell_1rw
* cell instance $23584 r0 *1 76.845,155.61
X$23584 283 629 284 644 645 cell_1rw
* cell instance $23585 m0 *1 76.845,158.34
X$23585 283 630 284 644 645 cell_1rw
* cell instance $23586 r0 *1 76.845,158.34
X$23586 283 631 284 644 645 cell_1rw
* cell instance $23587 m0 *1 76.845,161.07
X$23587 283 632 284 644 645 cell_1rw
* cell instance $23588 r0 *1 76.845,161.07
X$23588 283 633 284 644 645 cell_1rw
* cell instance $23589 m0 *1 76.845,163.8
X$23589 283 634 284 644 645 cell_1rw
* cell instance $23590 m0 *1 76.845,166.53
X$23590 283 637 284 644 645 cell_1rw
* cell instance $23591 r0 *1 76.845,163.8
X$23591 283 635 284 644 645 cell_1rw
* cell instance $23592 r0 *1 76.845,166.53
X$23592 283 636 284 644 645 cell_1rw
* cell instance $23593 m0 *1 76.845,169.26
X$23593 283 639 284 644 645 cell_1rw
* cell instance $23594 r0 *1 76.845,169.26
X$23594 283 638 284 644 645 cell_1rw
* cell instance $23595 m0 *1 76.845,171.99
X$23595 283 640 284 644 645 cell_1rw
* cell instance $23596 r0 *1 76.845,171.99
X$23596 283 641 284 644 645 cell_1rw
* cell instance $23597 m0 *1 76.845,174.72
X$23597 283 642 284 644 645 cell_1rw
* cell instance $23598 r0 *1 76.845,174.72
X$23598 283 643 284 644 645 cell_1rw
* cell instance $23599 r0 *1 77.55,87.36
X$23599 285 322 286 644 645 cell_1rw
* cell instance $23600 m0 *1 77.55,90.09
X$23600 285 581 286 644 645 cell_1rw
* cell instance $23601 r0 *1 77.55,90.09
X$23601 285 580 286 644 645 cell_1rw
* cell instance $23602 m0 *1 77.55,92.82
X$23602 285 583 286 644 645 cell_1rw
* cell instance $23603 r0 *1 77.55,92.82
X$23603 285 582 286 644 645 cell_1rw
* cell instance $23604 m0 *1 77.55,95.55
X$23604 285 584 286 644 645 cell_1rw
* cell instance $23605 r0 *1 77.55,95.55
X$23605 285 585 286 644 645 cell_1rw
* cell instance $23606 m0 *1 77.55,98.28
X$23606 285 586 286 644 645 cell_1rw
* cell instance $23607 r0 *1 77.55,98.28
X$23607 285 587 286 644 645 cell_1rw
* cell instance $23608 m0 *1 77.55,101.01
X$23608 285 588 286 644 645 cell_1rw
* cell instance $23609 r0 *1 77.55,101.01
X$23609 285 589 286 644 645 cell_1rw
* cell instance $23610 m0 *1 77.55,103.74
X$23610 285 590 286 644 645 cell_1rw
* cell instance $23611 r0 *1 77.55,103.74
X$23611 285 591 286 644 645 cell_1rw
* cell instance $23612 m0 *1 77.55,106.47
X$23612 285 593 286 644 645 cell_1rw
* cell instance $23613 r0 *1 77.55,106.47
X$23613 285 592 286 644 645 cell_1rw
* cell instance $23614 m0 *1 77.55,109.2
X$23614 285 594 286 644 645 cell_1rw
* cell instance $23615 r0 *1 77.55,109.2
X$23615 285 595 286 644 645 cell_1rw
* cell instance $23616 m0 *1 77.55,111.93
X$23616 285 597 286 644 645 cell_1rw
* cell instance $23617 r0 *1 77.55,111.93
X$23617 285 596 286 644 645 cell_1rw
* cell instance $23618 m0 *1 77.55,114.66
X$23618 285 598 286 644 645 cell_1rw
* cell instance $23619 r0 *1 77.55,114.66
X$23619 285 599 286 644 645 cell_1rw
* cell instance $23620 m0 *1 77.55,117.39
X$23620 285 600 286 644 645 cell_1rw
* cell instance $23621 r0 *1 77.55,117.39
X$23621 285 601 286 644 645 cell_1rw
* cell instance $23622 m0 *1 77.55,120.12
X$23622 285 602 286 644 645 cell_1rw
* cell instance $23623 r0 *1 77.55,120.12
X$23623 285 603 286 644 645 cell_1rw
* cell instance $23624 m0 *1 77.55,122.85
X$23624 285 604 286 644 645 cell_1rw
* cell instance $23625 r0 *1 77.55,122.85
X$23625 285 605 286 644 645 cell_1rw
* cell instance $23626 m0 *1 77.55,125.58
X$23626 285 606 286 644 645 cell_1rw
* cell instance $23627 r0 *1 77.55,125.58
X$23627 285 607 286 644 645 cell_1rw
* cell instance $23628 m0 *1 77.55,128.31
X$23628 285 609 286 644 645 cell_1rw
* cell instance $23629 r0 *1 77.55,128.31
X$23629 285 608 286 644 645 cell_1rw
* cell instance $23630 m0 *1 77.55,131.04
X$23630 285 610 286 644 645 cell_1rw
* cell instance $23631 r0 *1 77.55,131.04
X$23631 285 611 286 644 645 cell_1rw
* cell instance $23632 m0 *1 77.55,133.77
X$23632 285 612 286 644 645 cell_1rw
* cell instance $23633 r0 *1 77.55,133.77
X$23633 285 613 286 644 645 cell_1rw
* cell instance $23634 m0 *1 77.55,136.5
X$23634 285 615 286 644 645 cell_1rw
* cell instance $23635 r0 *1 77.55,136.5
X$23635 285 614 286 644 645 cell_1rw
* cell instance $23636 m0 *1 77.55,139.23
X$23636 285 617 286 644 645 cell_1rw
* cell instance $23637 r0 *1 77.55,139.23
X$23637 285 616 286 644 645 cell_1rw
* cell instance $23638 m0 *1 77.55,141.96
X$23638 285 618 286 644 645 cell_1rw
* cell instance $23639 r0 *1 77.55,141.96
X$23639 285 619 286 644 645 cell_1rw
* cell instance $23640 m0 *1 77.55,144.69
X$23640 285 620 286 644 645 cell_1rw
* cell instance $23641 m0 *1 77.55,147.42
X$23641 285 622 286 644 645 cell_1rw
* cell instance $23642 r0 *1 77.55,144.69
X$23642 285 621 286 644 645 cell_1rw
* cell instance $23643 r0 *1 77.55,147.42
X$23643 285 623 286 644 645 cell_1rw
* cell instance $23644 m0 *1 77.55,150.15
X$23644 285 624 286 644 645 cell_1rw
* cell instance $23645 r0 *1 77.55,150.15
X$23645 285 625 286 644 645 cell_1rw
* cell instance $23646 m0 *1 77.55,152.88
X$23646 285 626 286 644 645 cell_1rw
* cell instance $23647 r0 *1 77.55,152.88
X$23647 285 627 286 644 645 cell_1rw
* cell instance $23648 m0 *1 77.55,155.61
X$23648 285 628 286 644 645 cell_1rw
* cell instance $23649 r0 *1 77.55,155.61
X$23649 285 629 286 644 645 cell_1rw
* cell instance $23650 m0 *1 77.55,158.34
X$23650 285 630 286 644 645 cell_1rw
* cell instance $23651 r0 *1 77.55,158.34
X$23651 285 631 286 644 645 cell_1rw
* cell instance $23652 m0 *1 77.55,161.07
X$23652 285 632 286 644 645 cell_1rw
* cell instance $23653 r0 *1 77.55,161.07
X$23653 285 633 286 644 645 cell_1rw
* cell instance $23654 m0 *1 77.55,163.8
X$23654 285 634 286 644 645 cell_1rw
* cell instance $23655 r0 *1 77.55,163.8
X$23655 285 635 286 644 645 cell_1rw
* cell instance $23656 m0 *1 77.55,166.53
X$23656 285 637 286 644 645 cell_1rw
* cell instance $23657 r0 *1 77.55,166.53
X$23657 285 636 286 644 645 cell_1rw
* cell instance $23658 m0 *1 77.55,169.26
X$23658 285 639 286 644 645 cell_1rw
* cell instance $23659 r0 *1 77.55,169.26
X$23659 285 638 286 644 645 cell_1rw
* cell instance $23660 m0 *1 77.55,171.99
X$23660 285 640 286 644 645 cell_1rw
* cell instance $23661 m0 *1 77.55,174.72
X$23661 285 642 286 644 645 cell_1rw
* cell instance $23662 r0 *1 77.55,171.99
X$23662 285 641 286 644 645 cell_1rw
* cell instance $23663 r0 *1 77.55,174.72
X$23663 285 643 286 644 645 cell_1rw
* cell instance $23664 m0 *1 78.255,90.09
X$23664 287 581 288 644 645 cell_1rw
* cell instance $23665 r0 *1 78.255,87.36
X$23665 287 322 288 644 645 cell_1rw
* cell instance $23666 r0 *1 78.255,90.09
X$23666 287 580 288 644 645 cell_1rw
* cell instance $23667 m0 *1 78.255,92.82
X$23667 287 583 288 644 645 cell_1rw
* cell instance $23668 r0 *1 78.255,92.82
X$23668 287 582 288 644 645 cell_1rw
* cell instance $23669 m0 *1 78.255,95.55
X$23669 287 584 288 644 645 cell_1rw
* cell instance $23670 r0 *1 78.255,95.55
X$23670 287 585 288 644 645 cell_1rw
* cell instance $23671 m0 *1 78.255,98.28
X$23671 287 586 288 644 645 cell_1rw
* cell instance $23672 m0 *1 78.255,101.01
X$23672 287 588 288 644 645 cell_1rw
* cell instance $23673 r0 *1 78.255,98.28
X$23673 287 587 288 644 645 cell_1rw
* cell instance $23674 r0 *1 78.255,101.01
X$23674 287 589 288 644 645 cell_1rw
* cell instance $23675 m0 *1 78.255,103.74
X$23675 287 590 288 644 645 cell_1rw
* cell instance $23676 m0 *1 78.255,106.47
X$23676 287 593 288 644 645 cell_1rw
* cell instance $23677 r0 *1 78.255,103.74
X$23677 287 591 288 644 645 cell_1rw
* cell instance $23678 r0 *1 78.255,106.47
X$23678 287 592 288 644 645 cell_1rw
* cell instance $23679 m0 *1 78.255,109.2
X$23679 287 594 288 644 645 cell_1rw
* cell instance $23680 r0 *1 78.255,109.2
X$23680 287 595 288 644 645 cell_1rw
* cell instance $23681 m0 *1 78.255,111.93
X$23681 287 597 288 644 645 cell_1rw
* cell instance $23682 r0 *1 78.255,111.93
X$23682 287 596 288 644 645 cell_1rw
* cell instance $23683 m0 *1 78.255,114.66
X$23683 287 598 288 644 645 cell_1rw
* cell instance $23684 m0 *1 78.255,117.39
X$23684 287 600 288 644 645 cell_1rw
* cell instance $23685 r0 *1 78.255,114.66
X$23685 287 599 288 644 645 cell_1rw
* cell instance $23686 r0 *1 78.255,117.39
X$23686 287 601 288 644 645 cell_1rw
* cell instance $23687 m0 *1 78.255,120.12
X$23687 287 602 288 644 645 cell_1rw
* cell instance $23688 m0 *1 78.255,122.85
X$23688 287 604 288 644 645 cell_1rw
* cell instance $23689 r0 *1 78.255,120.12
X$23689 287 603 288 644 645 cell_1rw
* cell instance $23690 r0 *1 78.255,122.85
X$23690 287 605 288 644 645 cell_1rw
* cell instance $23691 m0 *1 78.255,125.58
X$23691 287 606 288 644 645 cell_1rw
* cell instance $23692 r0 *1 78.255,125.58
X$23692 287 607 288 644 645 cell_1rw
* cell instance $23693 m0 *1 78.255,128.31
X$23693 287 609 288 644 645 cell_1rw
* cell instance $23694 r0 *1 78.255,128.31
X$23694 287 608 288 644 645 cell_1rw
* cell instance $23695 m0 *1 78.255,131.04
X$23695 287 610 288 644 645 cell_1rw
* cell instance $23696 m0 *1 78.255,133.77
X$23696 287 612 288 644 645 cell_1rw
* cell instance $23697 r0 *1 78.255,131.04
X$23697 287 611 288 644 645 cell_1rw
* cell instance $23698 r0 *1 78.255,133.77
X$23698 287 613 288 644 645 cell_1rw
* cell instance $23699 m0 *1 78.255,136.5
X$23699 287 615 288 644 645 cell_1rw
* cell instance $23700 r0 *1 78.255,136.5
X$23700 287 614 288 644 645 cell_1rw
* cell instance $23701 m0 *1 78.255,139.23
X$23701 287 617 288 644 645 cell_1rw
* cell instance $23702 r0 *1 78.255,139.23
X$23702 287 616 288 644 645 cell_1rw
* cell instance $23703 m0 *1 78.255,141.96
X$23703 287 618 288 644 645 cell_1rw
* cell instance $23704 r0 *1 78.255,141.96
X$23704 287 619 288 644 645 cell_1rw
* cell instance $23705 m0 *1 78.255,144.69
X$23705 287 620 288 644 645 cell_1rw
* cell instance $23706 r0 *1 78.255,144.69
X$23706 287 621 288 644 645 cell_1rw
* cell instance $23707 m0 *1 78.255,147.42
X$23707 287 622 288 644 645 cell_1rw
* cell instance $23708 m0 *1 78.255,150.15
X$23708 287 624 288 644 645 cell_1rw
* cell instance $23709 r0 *1 78.255,147.42
X$23709 287 623 288 644 645 cell_1rw
* cell instance $23710 r0 *1 78.255,150.15
X$23710 287 625 288 644 645 cell_1rw
* cell instance $23711 m0 *1 78.255,152.88
X$23711 287 626 288 644 645 cell_1rw
* cell instance $23712 r0 *1 78.255,152.88
X$23712 287 627 288 644 645 cell_1rw
* cell instance $23713 m0 *1 78.255,155.61
X$23713 287 628 288 644 645 cell_1rw
* cell instance $23714 r0 *1 78.255,155.61
X$23714 287 629 288 644 645 cell_1rw
* cell instance $23715 m0 *1 78.255,158.34
X$23715 287 630 288 644 645 cell_1rw
* cell instance $23716 m0 *1 78.255,161.07
X$23716 287 632 288 644 645 cell_1rw
* cell instance $23717 r0 *1 78.255,158.34
X$23717 287 631 288 644 645 cell_1rw
* cell instance $23718 r0 *1 78.255,161.07
X$23718 287 633 288 644 645 cell_1rw
* cell instance $23719 m0 *1 78.255,163.8
X$23719 287 634 288 644 645 cell_1rw
* cell instance $23720 r0 *1 78.255,163.8
X$23720 287 635 288 644 645 cell_1rw
* cell instance $23721 m0 *1 78.255,166.53
X$23721 287 637 288 644 645 cell_1rw
* cell instance $23722 r0 *1 78.255,166.53
X$23722 287 636 288 644 645 cell_1rw
* cell instance $23723 m0 *1 78.255,169.26
X$23723 287 639 288 644 645 cell_1rw
* cell instance $23724 r0 *1 78.255,169.26
X$23724 287 638 288 644 645 cell_1rw
* cell instance $23725 m0 *1 78.255,171.99
X$23725 287 640 288 644 645 cell_1rw
* cell instance $23726 r0 *1 78.255,171.99
X$23726 287 641 288 644 645 cell_1rw
* cell instance $23727 m0 *1 78.255,174.72
X$23727 287 642 288 644 645 cell_1rw
* cell instance $23728 r0 *1 78.255,174.72
X$23728 287 643 288 644 645 cell_1rw
* cell instance $23729 r0 *1 78.96,87.36
X$23729 289 322 290 644 645 cell_1rw
* cell instance $23730 m0 *1 78.96,90.09
X$23730 289 581 290 644 645 cell_1rw
* cell instance $23731 r0 *1 78.96,90.09
X$23731 289 580 290 644 645 cell_1rw
* cell instance $23732 m0 *1 78.96,92.82
X$23732 289 583 290 644 645 cell_1rw
* cell instance $23733 m0 *1 78.96,95.55
X$23733 289 584 290 644 645 cell_1rw
* cell instance $23734 r0 *1 78.96,92.82
X$23734 289 582 290 644 645 cell_1rw
* cell instance $23735 r0 *1 78.96,95.55
X$23735 289 585 290 644 645 cell_1rw
* cell instance $23736 m0 *1 78.96,98.28
X$23736 289 586 290 644 645 cell_1rw
* cell instance $23737 r0 *1 78.96,98.28
X$23737 289 587 290 644 645 cell_1rw
* cell instance $23738 m0 *1 78.96,101.01
X$23738 289 588 290 644 645 cell_1rw
* cell instance $23739 m0 *1 78.96,103.74
X$23739 289 590 290 644 645 cell_1rw
* cell instance $23740 r0 *1 78.96,101.01
X$23740 289 589 290 644 645 cell_1rw
* cell instance $23741 r0 *1 78.96,103.74
X$23741 289 591 290 644 645 cell_1rw
* cell instance $23742 m0 *1 78.96,106.47
X$23742 289 593 290 644 645 cell_1rw
* cell instance $23743 r0 *1 78.96,106.47
X$23743 289 592 290 644 645 cell_1rw
* cell instance $23744 m0 *1 78.96,109.2
X$23744 289 594 290 644 645 cell_1rw
* cell instance $23745 r0 *1 78.96,109.2
X$23745 289 595 290 644 645 cell_1rw
* cell instance $23746 m0 *1 78.96,111.93
X$23746 289 597 290 644 645 cell_1rw
* cell instance $23747 r0 *1 78.96,111.93
X$23747 289 596 290 644 645 cell_1rw
* cell instance $23748 m0 *1 78.96,114.66
X$23748 289 598 290 644 645 cell_1rw
* cell instance $23749 r0 *1 78.96,114.66
X$23749 289 599 290 644 645 cell_1rw
* cell instance $23750 m0 *1 78.96,117.39
X$23750 289 600 290 644 645 cell_1rw
* cell instance $23751 r0 *1 78.96,117.39
X$23751 289 601 290 644 645 cell_1rw
* cell instance $23752 m0 *1 78.96,120.12
X$23752 289 602 290 644 645 cell_1rw
* cell instance $23753 r0 *1 78.96,120.12
X$23753 289 603 290 644 645 cell_1rw
* cell instance $23754 m0 *1 78.96,122.85
X$23754 289 604 290 644 645 cell_1rw
* cell instance $23755 r0 *1 78.96,122.85
X$23755 289 605 290 644 645 cell_1rw
* cell instance $23756 m0 *1 78.96,125.58
X$23756 289 606 290 644 645 cell_1rw
* cell instance $23757 r0 *1 78.96,125.58
X$23757 289 607 290 644 645 cell_1rw
* cell instance $23758 m0 *1 78.96,128.31
X$23758 289 609 290 644 645 cell_1rw
* cell instance $23759 r0 *1 78.96,128.31
X$23759 289 608 290 644 645 cell_1rw
* cell instance $23760 m0 *1 78.96,131.04
X$23760 289 610 290 644 645 cell_1rw
* cell instance $23761 r0 *1 78.96,131.04
X$23761 289 611 290 644 645 cell_1rw
* cell instance $23762 m0 *1 78.96,133.77
X$23762 289 612 290 644 645 cell_1rw
* cell instance $23763 r0 *1 78.96,133.77
X$23763 289 613 290 644 645 cell_1rw
* cell instance $23764 m0 *1 78.96,136.5
X$23764 289 615 290 644 645 cell_1rw
* cell instance $23765 r0 *1 78.96,136.5
X$23765 289 614 290 644 645 cell_1rw
* cell instance $23766 m0 *1 78.96,139.23
X$23766 289 617 290 644 645 cell_1rw
* cell instance $23767 r0 *1 78.96,139.23
X$23767 289 616 290 644 645 cell_1rw
* cell instance $23768 m0 *1 78.96,141.96
X$23768 289 618 290 644 645 cell_1rw
* cell instance $23769 r0 *1 78.96,141.96
X$23769 289 619 290 644 645 cell_1rw
* cell instance $23770 m0 *1 78.96,144.69
X$23770 289 620 290 644 645 cell_1rw
* cell instance $23771 r0 *1 78.96,144.69
X$23771 289 621 290 644 645 cell_1rw
* cell instance $23772 m0 *1 78.96,147.42
X$23772 289 622 290 644 645 cell_1rw
* cell instance $23773 r0 *1 78.96,147.42
X$23773 289 623 290 644 645 cell_1rw
* cell instance $23774 m0 *1 78.96,150.15
X$23774 289 624 290 644 645 cell_1rw
* cell instance $23775 r0 *1 78.96,150.15
X$23775 289 625 290 644 645 cell_1rw
* cell instance $23776 m0 *1 78.96,152.88
X$23776 289 626 290 644 645 cell_1rw
* cell instance $23777 r0 *1 78.96,152.88
X$23777 289 627 290 644 645 cell_1rw
* cell instance $23778 m0 *1 78.96,155.61
X$23778 289 628 290 644 645 cell_1rw
* cell instance $23779 m0 *1 78.96,158.34
X$23779 289 630 290 644 645 cell_1rw
* cell instance $23780 r0 *1 78.96,155.61
X$23780 289 629 290 644 645 cell_1rw
* cell instance $23781 r0 *1 78.96,158.34
X$23781 289 631 290 644 645 cell_1rw
* cell instance $23782 m0 *1 78.96,161.07
X$23782 289 632 290 644 645 cell_1rw
* cell instance $23783 m0 *1 78.96,163.8
X$23783 289 634 290 644 645 cell_1rw
* cell instance $23784 r0 *1 78.96,161.07
X$23784 289 633 290 644 645 cell_1rw
* cell instance $23785 r0 *1 78.96,163.8
X$23785 289 635 290 644 645 cell_1rw
* cell instance $23786 m0 *1 78.96,166.53
X$23786 289 637 290 644 645 cell_1rw
* cell instance $23787 r0 *1 78.96,166.53
X$23787 289 636 290 644 645 cell_1rw
* cell instance $23788 m0 *1 78.96,169.26
X$23788 289 639 290 644 645 cell_1rw
* cell instance $23789 m0 *1 78.96,171.99
X$23789 289 640 290 644 645 cell_1rw
* cell instance $23790 r0 *1 78.96,169.26
X$23790 289 638 290 644 645 cell_1rw
* cell instance $23791 m0 *1 78.96,174.72
X$23791 289 642 290 644 645 cell_1rw
* cell instance $23792 r0 *1 78.96,171.99
X$23792 289 641 290 644 645 cell_1rw
* cell instance $23793 r0 *1 78.96,174.72
X$23793 289 643 290 644 645 cell_1rw
* cell instance $23794 r0 *1 79.665,87.36
X$23794 291 322 292 644 645 cell_1rw
* cell instance $23795 m0 *1 79.665,90.09
X$23795 291 581 292 644 645 cell_1rw
* cell instance $23796 r0 *1 79.665,90.09
X$23796 291 580 292 644 645 cell_1rw
* cell instance $23797 m0 *1 79.665,92.82
X$23797 291 583 292 644 645 cell_1rw
* cell instance $23798 r0 *1 79.665,92.82
X$23798 291 582 292 644 645 cell_1rw
* cell instance $23799 m0 *1 79.665,95.55
X$23799 291 584 292 644 645 cell_1rw
* cell instance $23800 r0 *1 79.665,95.55
X$23800 291 585 292 644 645 cell_1rw
* cell instance $23801 m0 *1 79.665,98.28
X$23801 291 586 292 644 645 cell_1rw
* cell instance $23802 m0 *1 79.665,101.01
X$23802 291 588 292 644 645 cell_1rw
* cell instance $23803 r0 *1 79.665,98.28
X$23803 291 587 292 644 645 cell_1rw
* cell instance $23804 r0 *1 79.665,101.01
X$23804 291 589 292 644 645 cell_1rw
* cell instance $23805 m0 *1 79.665,103.74
X$23805 291 590 292 644 645 cell_1rw
* cell instance $23806 m0 *1 79.665,106.47
X$23806 291 593 292 644 645 cell_1rw
* cell instance $23807 r0 *1 79.665,103.74
X$23807 291 591 292 644 645 cell_1rw
* cell instance $23808 r0 *1 79.665,106.47
X$23808 291 592 292 644 645 cell_1rw
* cell instance $23809 m0 *1 79.665,109.2
X$23809 291 594 292 644 645 cell_1rw
* cell instance $23810 r0 *1 79.665,109.2
X$23810 291 595 292 644 645 cell_1rw
* cell instance $23811 m0 *1 79.665,111.93
X$23811 291 597 292 644 645 cell_1rw
* cell instance $23812 r0 *1 79.665,111.93
X$23812 291 596 292 644 645 cell_1rw
* cell instance $23813 m0 *1 79.665,114.66
X$23813 291 598 292 644 645 cell_1rw
* cell instance $23814 r0 *1 79.665,114.66
X$23814 291 599 292 644 645 cell_1rw
* cell instance $23815 m0 *1 79.665,117.39
X$23815 291 600 292 644 645 cell_1rw
* cell instance $23816 r0 *1 79.665,117.39
X$23816 291 601 292 644 645 cell_1rw
* cell instance $23817 m0 *1 79.665,120.12
X$23817 291 602 292 644 645 cell_1rw
* cell instance $23818 r0 *1 79.665,120.12
X$23818 291 603 292 644 645 cell_1rw
* cell instance $23819 m0 *1 79.665,122.85
X$23819 291 604 292 644 645 cell_1rw
* cell instance $23820 r0 *1 79.665,122.85
X$23820 291 605 292 644 645 cell_1rw
* cell instance $23821 m0 *1 79.665,125.58
X$23821 291 606 292 644 645 cell_1rw
* cell instance $23822 r0 *1 79.665,125.58
X$23822 291 607 292 644 645 cell_1rw
* cell instance $23823 m0 *1 79.665,128.31
X$23823 291 609 292 644 645 cell_1rw
* cell instance $23824 r0 *1 79.665,128.31
X$23824 291 608 292 644 645 cell_1rw
* cell instance $23825 m0 *1 79.665,131.04
X$23825 291 610 292 644 645 cell_1rw
* cell instance $23826 r0 *1 79.665,131.04
X$23826 291 611 292 644 645 cell_1rw
* cell instance $23827 m0 *1 79.665,133.77
X$23827 291 612 292 644 645 cell_1rw
* cell instance $23828 r0 *1 79.665,133.77
X$23828 291 613 292 644 645 cell_1rw
* cell instance $23829 m0 *1 79.665,136.5
X$23829 291 615 292 644 645 cell_1rw
* cell instance $23830 m0 *1 79.665,139.23
X$23830 291 617 292 644 645 cell_1rw
* cell instance $23831 r0 *1 79.665,136.5
X$23831 291 614 292 644 645 cell_1rw
* cell instance $23832 m0 *1 79.665,141.96
X$23832 291 618 292 644 645 cell_1rw
* cell instance $23833 r0 *1 79.665,139.23
X$23833 291 616 292 644 645 cell_1rw
* cell instance $23834 r0 *1 79.665,141.96
X$23834 291 619 292 644 645 cell_1rw
* cell instance $23835 m0 *1 79.665,144.69
X$23835 291 620 292 644 645 cell_1rw
* cell instance $23836 r0 *1 79.665,144.69
X$23836 291 621 292 644 645 cell_1rw
* cell instance $23837 m0 *1 79.665,147.42
X$23837 291 622 292 644 645 cell_1rw
* cell instance $23838 r0 *1 79.665,147.42
X$23838 291 623 292 644 645 cell_1rw
* cell instance $23839 m0 *1 79.665,150.15
X$23839 291 624 292 644 645 cell_1rw
* cell instance $23840 r0 *1 79.665,150.15
X$23840 291 625 292 644 645 cell_1rw
* cell instance $23841 m0 *1 79.665,152.88
X$23841 291 626 292 644 645 cell_1rw
* cell instance $23842 r0 *1 79.665,152.88
X$23842 291 627 292 644 645 cell_1rw
* cell instance $23843 m0 *1 79.665,155.61
X$23843 291 628 292 644 645 cell_1rw
* cell instance $23844 r0 *1 79.665,155.61
X$23844 291 629 292 644 645 cell_1rw
* cell instance $23845 m0 *1 79.665,158.34
X$23845 291 630 292 644 645 cell_1rw
* cell instance $23846 r0 *1 79.665,158.34
X$23846 291 631 292 644 645 cell_1rw
* cell instance $23847 m0 *1 79.665,161.07
X$23847 291 632 292 644 645 cell_1rw
* cell instance $23848 r0 *1 79.665,161.07
X$23848 291 633 292 644 645 cell_1rw
* cell instance $23849 m0 *1 79.665,163.8
X$23849 291 634 292 644 645 cell_1rw
* cell instance $23850 r0 *1 79.665,163.8
X$23850 291 635 292 644 645 cell_1rw
* cell instance $23851 m0 *1 79.665,166.53
X$23851 291 637 292 644 645 cell_1rw
* cell instance $23852 r0 *1 79.665,166.53
X$23852 291 636 292 644 645 cell_1rw
* cell instance $23853 m0 *1 79.665,169.26
X$23853 291 639 292 644 645 cell_1rw
* cell instance $23854 r0 *1 79.665,169.26
X$23854 291 638 292 644 645 cell_1rw
* cell instance $23855 m0 *1 79.665,171.99
X$23855 291 640 292 644 645 cell_1rw
* cell instance $23856 m0 *1 79.665,174.72
X$23856 291 642 292 644 645 cell_1rw
* cell instance $23857 r0 *1 79.665,171.99
X$23857 291 641 292 644 645 cell_1rw
* cell instance $23858 r0 *1 79.665,174.72
X$23858 291 643 292 644 645 cell_1rw
* cell instance $23859 m0 *1 80.37,90.09
X$23859 293 581 294 644 645 cell_1rw
* cell instance $23860 r0 *1 80.37,87.36
X$23860 293 322 294 644 645 cell_1rw
* cell instance $23861 r0 *1 80.37,90.09
X$23861 293 580 294 644 645 cell_1rw
* cell instance $23862 m0 *1 80.37,92.82
X$23862 293 583 294 644 645 cell_1rw
* cell instance $23863 r0 *1 80.37,92.82
X$23863 293 582 294 644 645 cell_1rw
* cell instance $23864 m0 *1 80.37,95.55
X$23864 293 584 294 644 645 cell_1rw
* cell instance $23865 m0 *1 80.37,98.28
X$23865 293 586 294 644 645 cell_1rw
* cell instance $23866 r0 *1 80.37,95.55
X$23866 293 585 294 644 645 cell_1rw
* cell instance $23867 r0 *1 80.37,98.28
X$23867 293 587 294 644 645 cell_1rw
* cell instance $23868 m0 *1 80.37,101.01
X$23868 293 588 294 644 645 cell_1rw
* cell instance $23869 r0 *1 80.37,101.01
X$23869 293 589 294 644 645 cell_1rw
* cell instance $23870 m0 *1 80.37,103.74
X$23870 293 590 294 644 645 cell_1rw
* cell instance $23871 r0 *1 80.37,103.74
X$23871 293 591 294 644 645 cell_1rw
* cell instance $23872 m0 *1 80.37,106.47
X$23872 293 593 294 644 645 cell_1rw
* cell instance $23873 r0 *1 80.37,106.47
X$23873 293 592 294 644 645 cell_1rw
* cell instance $23874 m0 *1 80.37,109.2
X$23874 293 594 294 644 645 cell_1rw
* cell instance $23875 r0 *1 80.37,109.2
X$23875 293 595 294 644 645 cell_1rw
* cell instance $23876 m0 *1 80.37,111.93
X$23876 293 597 294 644 645 cell_1rw
* cell instance $23877 m0 *1 80.37,114.66
X$23877 293 598 294 644 645 cell_1rw
* cell instance $23878 r0 *1 80.37,111.93
X$23878 293 596 294 644 645 cell_1rw
* cell instance $23879 r0 *1 80.37,114.66
X$23879 293 599 294 644 645 cell_1rw
* cell instance $23880 m0 *1 80.37,117.39
X$23880 293 600 294 644 645 cell_1rw
* cell instance $23881 m0 *1 80.37,120.12
X$23881 293 602 294 644 645 cell_1rw
* cell instance $23882 r0 *1 80.37,117.39
X$23882 293 601 294 644 645 cell_1rw
* cell instance $23883 m0 *1 80.37,122.85
X$23883 293 604 294 644 645 cell_1rw
* cell instance $23884 r0 *1 80.37,120.12
X$23884 293 603 294 644 645 cell_1rw
* cell instance $23885 r0 *1 80.37,122.85
X$23885 293 605 294 644 645 cell_1rw
* cell instance $23886 m0 *1 80.37,125.58
X$23886 293 606 294 644 645 cell_1rw
* cell instance $23887 r0 *1 80.37,125.58
X$23887 293 607 294 644 645 cell_1rw
* cell instance $23888 m0 *1 80.37,128.31
X$23888 293 609 294 644 645 cell_1rw
* cell instance $23889 r0 *1 80.37,128.31
X$23889 293 608 294 644 645 cell_1rw
* cell instance $23890 m0 *1 80.37,131.04
X$23890 293 610 294 644 645 cell_1rw
* cell instance $23891 r0 *1 80.37,131.04
X$23891 293 611 294 644 645 cell_1rw
* cell instance $23892 m0 *1 80.37,133.77
X$23892 293 612 294 644 645 cell_1rw
* cell instance $23893 r0 *1 80.37,133.77
X$23893 293 613 294 644 645 cell_1rw
* cell instance $23894 m0 *1 80.37,136.5
X$23894 293 615 294 644 645 cell_1rw
* cell instance $23895 r0 *1 80.37,136.5
X$23895 293 614 294 644 645 cell_1rw
* cell instance $23896 m0 *1 80.37,139.23
X$23896 293 617 294 644 645 cell_1rw
* cell instance $23897 r0 *1 80.37,139.23
X$23897 293 616 294 644 645 cell_1rw
* cell instance $23898 m0 *1 80.37,141.96
X$23898 293 618 294 644 645 cell_1rw
* cell instance $23899 m0 *1 80.37,144.69
X$23899 293 620 294 644 645 cell_1rw
* cell instance $23900 r0 *1 80.37,141.96
X$23900 293 619 294 644 645 cell_1rw
* cell instance $23901 r0 *1 80.37,144.69
X$23901 293 621 294 644 645 cell_1rw
* cell instance $23902 m0 *1 80.37,147.42
X$23902 293 622 294 644 645 cell_1rw
* cell instance $23903 r0 *1 80.37,147.42
X$23903 293 623 294 644 645 cell_1rw
* cell instance $23904 m0 *1 80.37,150.15
X$23904 293 624 294 644 645 cell_1rw
* cell instance $23905 r0 *1 80.37,150.15
X$23905 293 625 294 644 645 cell_1rw
* cell instance $23906 m0 *1 80.37,152.88
X$23906 293 626 294 644 645 cell_1rw
* cell instance $23907 r0 *1 80.37,152.88
X$23907 293 627 294 644 645 cell_1rw
* cell instance $23908 m0 *1 80.37,155.61
X$23908 293 628 294 644 645 cell_1rw
* cell instance $23909 r0 *1 80.37,155.61
X$23909 293 629 294 644 645 cell_1rw
* cell instance $23910 m0 *1 80.37,158.34
X$23910 293 630 294 644 645 cell_1rw
* cell instance $23911 r0 *1 80.37,158.34
X$23911 293 631 294 644 645 cell_1rw
* cell instance $23912 m0 *1 80.37,161.07
X$23912 293 632 294 644 645 cell_1rw
* cell instance $23913 r0 *1 80.37,161.07
X$23913 293 633 294 644 645 cell_1rw
* cell instance $23914 m0 *1 80.37,163.8
X$23914 293 634 294 644 645 cell_1rw
* cell instance $23915 m0 *1 80.37,166.53
X$23915 293 637 294 644 645 cell_1rw
* cell instance $23916 r0 *1 80.37,163.8
X$23916 293 635 294 644 645 cell_1rw
* cell instance $23917 m0 *1 80.37,169.26
X$23917 293 639 294 644 645 cell_1rw
* cell instance $23918 r0 *1 80.37,166.53
X$23918 293 636 294 644 645 cell_1rw
* cell instance $23919 r0 *1 80.37,169.26
X$23919 293 638 294 644 645 cell_1rw
* cell instance $23920 m0 *1 80.37,171.99
X$23920 293 640 294 644 645 cell_1rw
* cell instance $23921 r0 *1 80.37,171.99
X$23921 293 641 294 644 645 cell_1rw
* cell instance $23922 m0 *1 80.37,174.72
X$23922 293 642 294 644 645 cell_1rw
* cell instance $23923 r0 *1 80.37,174.72
X$23923 293 643 294 644 645 cell_1rw
* cell instance $23924 r0 *1 81.075,87.36
X$23924 295 322 296 644 645 cell_1rw
* cell instance $23925 m0 *1 81.075,90.09
X$23925 295 581 296 644 645 cell_1rw
* cell instance $23926 r0 *1 81.075,90.09
X$23926 295 580 296 644 645 cell_1rw
* cell instance $23927 m0 *1 81.075,92.82
X$23927 295 583 296 644 645 cell_1rw
* cell instance $23928 r0 *1 81.075,92.82
X$23928 295 582 296 644 645 cell_1rw
* cell instance $23929 m0 *1 81.075,95.55
X$23929 295 584 296 644 645 cell_1rw
* cell instance $23930 m0 *1 81.075,98.28
X$23930 295 586 296 644 645 cell_1rw
* cell instance $23931 r0 *1 81.075,95.55
X$23931 295 585 296 644 645 cell_1rw
* cell instance $23932 r0 *1 81.075,98.28
X$23932 295 587 296 644 645 cell_1rw
* cell instance $23933 m0 *1 81.075,101.01
X$23933 295 588 296 644 645 cell_1rw
* cell instance $23934 m0 *1 81.075,103.74
X$23934 295 590 296 644 645 cell_1rw
* cell instance $23935 r0 *1 81.075,101.01
X$23935 295 589 296 644 645 cell_1rw
* cell instance $23936 r0 *1 81.075,103.74
X$23936 295 591 296 644 645 cell_1rw
* cell instance $23937 m0 *1 81.075,106.47
X$23937 295 593 296 644 645 cell_1rw
* cell instance $23938 r0 *1 81.075,106.47
X$23938 295 592 296 644 645 cell_1rw
* cell instance $23939 m0 *1 81.075,109.2
X$23939 295 594 296 644 645 cell_1rw
* cell instance $23940 m0 *1 81.075,111.93
X$23940 295 597 296 644 645 cell_1rw
* cell instance $23941 r0 *1 81.075,109.2
X$23941 295 595 296 644 645 cell_1rw
* cell instance $23942 r0 *1 81.075,111.93
X$23942 295 596 296 644 645 cell_1rw
* cell instance $23943 m0 *1 81.075,114.66
X$23943 295 598 296 644 645 cell_1rw
* cell instance $23944 r0 *1 81.075,114.66
X$23944 295 599 296 644 645 cell_1rw
* cell instance $23945 m0 *1 81.075,117.39
X$23945 295 600 296 644 645 cell_1rw
* cell instance $23946 m0 *1 81.075,120.12
X$23946 295 602 296 644 645 cell_1rw
* cell instance $23947 r0 *1 81.075,117.39
X$23947 295 601 296 644 645 cell_1rw
* cell instance $23948 r0 *1 81.075,120.12
X$23948 295 603 296 644 645 cell_1rw
* cell instance $23949 m0 *1 81.075,122.85
X$23949 295 604 296 644 645 cell_1rw
* cell instance $23950 r0 *1 81.075,122.85
X$23950 295 605 296 644 645 cell_1rw
* cell instance $23951 m0 *1 81.075,125.58
X$23951 295 606 296 644 645 cell_1rw
* cell instance $23952 r0 *1 81.075,125.58
X$23952 295 607 296 644 645 cell_1rw
* cell instance $23953 m0 *1 81.075,128.31
X$23953 295 609 296 644 645 cell_1rw
* cell instance $23954 m0 *1 81.075,131.04
X$23954 295 610 296 644 645 cell_1rw
* cell instance $23955 r0 *1 81.075,128.31
X$23955 295 608 296 644 645 cell_1rw
* cell instance $23956 r0 *1 81.075,131.04
X$23956 295 611 296 644 645 cell_1rw
* cell instance $23957 m0 *1 81.075,133.77
X$23957 295 612 296 644 645 cell_1rw
* cell instance $23958 r0 *1 81.075,133.77
X$23958 295 613 296 644 645 cell_1rw
* cell instance $23959 m0 *1 81.075,136.5
X$23959 295 615 296 644 645 cell_1rw
* cell instance $23960 r0 *1 81.075,136.5
X$23960 295 614 296 644 645 cell_1rw
* cell instance $23961 m0 *1 81.075,139.23
X$23961 295 617 296 644 645 cell_1rw
* cell instance $23962 r0 *1 81.075,139.23
X$23962 295 616 296 644 645 cell_1rw
* cell instance $23963 m0 *1 81.075,141.96
X$23963 295 618 296 644 645 cell_1rw
* cell instance $23964 r0 *1 81.075,141.96
X$23964 295 619 296 644 645 cell_1rw
* cell instance $23965 m0 *1 81.075,144.69
X$23965 295 620 296 644 645 cell_1rw
* cell instance $23966 r0 *1 81.075,144.69
X$23966 295 621 296 644 645 cell_1rw
* cell instance $23967 m0 *1 81.075,147.42
X$23967 295 622 296 644 645 cell_1rw
* cell instance $23968 r0 *1 81.075,147.42
X$23968 295 623 296 644 645 cell_1rw
* cell instance $23969 m0 *1 81.075,150.15
X$23969 295 624 296 644 645 cell_1rw
* cell instance $23970 r0 *1 81.075,150.15
X$23970 295 625 296 644 645 cell_1rw
* cell instance $23971 m0 *1 81.075,152.88
X$23971 295 626 296 644 645 cell_1rw
* cell instance $23972 r0 *1 81.075,152.88
X$23972 295 627 296 644 645 cell_1rw
* cell instance $23973 m0 *1 81.075,155.61
X$23973 295 628 296 644 645 cell_1rw
* cell instance $23974 r0 *1 81.075,155.61
X$23974 295 629 296 644 645 cell_1rw
* cell instance $23975 m0 *1 81.075,158.34
X$23975 295 630 296 644 645 cell_1rw
* cell instance $23976 m0 *1 81.075,161.07
X$23976 295 632 296 644 645 cell_1rw
* cell instance $23977 r0 *1 81.075,158.34
X$23977 295 631 296 644 645 cell_1rw
* cell instance $23978 r0 *1 81.075,161.07
X$23978 295 633 296 644 645 cell_1rw
* cell instance $23979 m0 *1 81.075,163.8
X$23979 295 634 296 644 645 cell_1rw
* cell instance $23980 r0 *1 81.075,163.8
X$23980 295 635 296 644 645 cell_1rw
* cell instance $23981 m0 *1 81.075,166.53
X$23981 295 637 296 644 645 cell_1rw
* cell instance $23982 r0 *1 81.075,166.53
X$23982 295 636 296 644 645 cell_1rw
* cell instance $23983 m0 *1 81.075,169.26
X$23983 295 639 296 644 645 cell_1rw
* cell instance $23984 m0 *1 81.075,171.99
X$23984 295 640 296 644 645 cell_1rw
* cell instance $23985 r0 *1 81.075,169.26
X$23985 295 638 296 644 645 cell_1rw
* cell instance $23986 r0 *1 81.075,171.99
X$23986 295 641 296 644 645 cell_1rw
* cell instance $23987 m0 *1 81.075,174.72
X$23987 295 642 296 644 645 cell_1rw
* cell instance $23988 r0 *1 81.075,174.72
X$23988 295 643 296 644 645 cell_1rw
* cell instance $23989 r0 *1 81.78,87.36
X$23989 297 322 298 644 645 cell_1rw
* cell instance $23990 m0 *1 81.78,90.09
X$23990 297 581 298 644 645 cell_1rw
* cell instance $23991 r0 *1 81.78,90.09
X$23991 297 580 298 644 645 cell_1rw
* cell instance $23992 m0 *1 81.78,92.82
X$23992 297 583 298 644 645 cell_1rw
* cell instance $23993 r0 *1 81.78,92.82
X$23993 297 582 298 644 645 cell_1rw
* cell instance $23994 m0 *1 81.78,95.55
X$23994 297 584 298 644 645 cell_1rw
* cell instance $23995 r0 *1 81.78,95.55
X$23995 297 585 298 644 645 cell_1rw
* cell instance $23996 m0 *1 81.78,98.28
X$23996 297 586 298 644 645 cell_1rw
* cell instance $23997 r0 *1 81.78,98.28
X$23997 297 587 298 644 645 cell_1rw
* cell instance $23998 m0 *1 81.78,101.01
X$23998 297 588 298 644 645 cell_1rw
* cell instance $23999 r0 *1 81.78,101.01
X$23999 297 589 298 644 645 cell_1rw
* cell instance $24000 m0 *1 81.78,103.74
X$24000 297 590 298 644 645 cell_1rw
* cell instance $24001 r0 *1 81.78,103.74
X$24001 297 591 298 644 645 cell_1rw
* cell instance $24002 m0 *1 81.78,106.47
X$24002 297 593 298 644 645 cell_1rw
* cell instance $24003 m0 *1 81.78,109.2
X$24003 297 594 298 644 645 cell_1rw
* cell instance $24004 r0 *1 81.78,106.47
X$24004 297 592 298 644 645 cell_1rw
* cell instance $24005 r0 *1 81.78,109.2
X$24005 297 595 298 644 645 cell_1rw
* cell instance $24006 m0 *1 81.78,111.93
X$24006 297 597 298 644 645 cell_1rw
* cell instance $24007 m0 *1 81.78,114.66
X$24007 297 598 298 644 645 cell_1rw
* cell instance $24008 r0 *1 81.78,111.93
X$24008 297 596 298 644 645 cell_1rw
* cell instance $24009 r0 *1 81.78,114.66
X$24009 297 599 298 644 645 cell_1rw
* cell instance $24010 m0 *1 81.78,117.39
X$24010 297 600 298 644 645 cell_1rw
* cell instance $24011 r0 *1 81.78,117.39
X$24011 297 601 298 644 645 cell_1rw
* cell instance $24012 m0 *1 81.78,120.12
X$24012 297 602 298 644 645 cell_1rw
* cell instance $24013 r0 *1 81.78,120.12
X$24013 297 603 298 644 645 cell_1rw
* cell instance $24014 m0 *1 81.78,122.85
X$24014 297 604 298 644 645 cell_1rw
* cell instance $24015 r0 *1 81.78,122.85
X$24015 297 605 298 644 645 cell_1rw
* cell instance $24016 m0 *1 81.78,125.58
X$24016 297 606 298 644 645 cell_1rw
* cell instance $24017 r0 *1 81.78,125.58
X$24017 297 607 298 644 645 cell_1rw
* cell instance $24018 m0 *1 81.78,128.31
X$24018 297 609 298 644 645 cell_1rw
* cell instance $24019 r0 *1 81.78,128.31
X$24019 297 608 298 644 645 cell_1rw
* cell instance $24020 m0 *1 81.78,131.04
X$24020 297 610 298 644 645 cell_1rw
* cell instance $24021 r0 *1 81.78,131.04
X$24021 297 611 298 644 645 cell_1rw
* cell instance $24022 m0 *1 81.78,133.77
X$24022 297 612 298 644 645 cell_1rw
* cell instance $24023 m0 *1 81.78,136.5
X$24023 297 615 298 644 645 cell_1rw
* cell instance $24024 r0 *1 81.78,133.77
X$24024 297 613 298 644 645 cell_1rw
* cell instance $24025 r0 *1 81.78,136.5
X$24025 297 614 298 644 645 cell_1rw
* cell instance $24026 m0 *1 81.78,139.23
X$24026 297 617 298 644 645 cell_1rw
* cell instance $24027 m0 *1 81.78,141.96
X$24027 297 618 298 644 645 cell_1rw
* cell instance $24028 r0 *1 81.78,139.23
X$24028 297 616 298 644 645 cell_1rw
* cell instance $24029 r0 *1 81.78,141.96
X$24029 297 619 298 644 645 cell_1rw
* cell instance $24030 m0 *1 81.78,144.69
X$24030 297 620 298 644 645 cell_1rw
* cell instance $24031 r0 *1 81.78,144.69
X$24031 297 621 298 644 645 cell_1rw
* cell instance $24032 m0 *1 81.78,147.42
X$24032 297 622 298 644 645 cell_1rw
* cell instance $24033 m0 *1 81.78,150.15
X$24033 297 624 298 644 645 cell_1rw
* cell instance $24034 r0 *1 81.78,147.42
X$24034 297 623 298 644 645 cell_1rw
* cell instance $24035 r0 *1 81.78,150.15
X$24035 297 625 298 644 645 cell_1rw
* cell instance $24036 m0 *1 81.78,152.88
X$24036 297 626 298 644 645 cell_1rw
* cell instance $24037 r0 *1 81.78,152.88
X$24037 297 627 298 644 645 cell_1rw
* cell instance $24038 m0 *1 81.78,155.61
X$24038 297 628 298 644 645 cell_1rw
* cell instance $24039 m0 *1 81.78,158.34
X$24039 297 630 298 644 645 cell_1rw
* cell instance $24040 r0 *1 81.78,155.61
X$24040 297 629 298 644 645 cell_1rw
* cell instance $24041 r0 *1 81.78,158.34
X$24041 297 631 298 644 645 cell_1rw
* cell instance $24042 m0 *1 81.78,161.07
X$24042 297 632 298 644 645 cell_1rw
* cell instance $24043 r0 *1 81.78,161.07
X$24043 297 633 298 644 645 cell_1rw
* cell instance $24044 m0 *1 81.78,163.8
X$24044 297 634 298 644 645 cell_1rw
* cell instance $24045 r0 *1 81.78,163.8
X$24045 297 635 298 644 645 cell_1rw
* cell instance $24046 m0 *1 81.78,166.53
X$24046 297 637 298 644 645 cell_1rw
* cell instance $24047 r0 *1 81.78,166.53
X$24047 297 636 298 644 645 cell_1rw
* cell instance $24048 m0 *1 81.78,169.26
X$24048 297 639 298 644 645 cell_1rw
* cell instance $24049 r0 *1 81.78,169.26
X$24049 297 638 298 644 645 cell_1rw
* cell instance $24050 m0 *1 81.78,171.99
X$24050 297 640 298 644 645 cell_1rw
* cell instance $24051 r0 *1 81.78,171.99
X$24051 297 641 298 644 645 cell_1rw
* cell instance $24052 m0 *1 81.78,174.72
X$24052 297 642 298 644 645 cell_1rw
* cell instance $24053 r0 *1 81.78,174.72
X$24053 297 643 298 644 645 cell_1rw
* cell instance $24054 r0 *1 82.485,87.36
X$24054 299 322 300 644 645 cell_1rw
* cell instance $24055 m0 *1 82.485,90.09
X$24055 299 581 300 644 645 cell_1rw
* cell instance $24056 r0 *1 82.485,90.09
X$24056 299 580 300 644 645 cell_1rw
* cell instance $24057 m0 *1 82.485,92.82
X$24057 299 583 300 644 645 cell_1rw
* cell instance $24058 m0 *1 82.485,95.55
X$24058 299 584 300 644 645 cell_1rw
* cell instance $24059 r0 *1 82.485,92.82
X$24059 299 582 300 644 645 cell_1rw
* cell instance $24060 r0 *1 82.485,95.55
X$24060 299 585 300 644 645 cell_1rw
* cell instance $24061 m0 *1 82.485,98.28
X$24061 299 586 300 644 645 cell_1rw
* cell instance $24062 r0 *1 82.485,98.28
X$24062 299 587 300 644 645 cell_1rw
* cell instance $24063 m0 *1 82.485,101.01
X$24063 299 588 300 644 645 cell_1rw
* cell instance $24064 m0 *1 82.485,103.74
X$24064 299 590 300 644 645 cell_1rw
* cell instance $24065 r0 *1 82.485,101.01
X$24065 299 589 300 644 645 cell_1rw
* cell instance $24066 r0 *1 82.485,103.74
X$24066 299 591 300 644 645 cell_1rw
* cell instance $24067 m0 *1 82.485,106.47
X$24067 299 593 300 644 645 cell_1rw
* cell instance $24068 r0 *1 82.485,106.47
X$24068 299 592 300 644 645 cell_1rw
* cell instance $24069 m0 *1 82.485,109.2
X$24069 299 594 300 644 645 cell_1rw
* cell instance $24070 r0 *1 82.485,109.2
X$24070 299 595 300 644 645 cell_1rw
* cell instance $24071 m0 *1 82.485,111.93
X$24071 299 597 300 644 645 cell_1rw
* cell instance $24072 r0 *1 82.485,111.93
X$24072 299 596 300 644 645 cell_1rw
* cell instance $24073 m0 *1 82.485,114.66
X$24073 299 598 300 644 645 cell_1rw
* cell instance $24074 r0 *1 82.485,114.66
X$24074 299 599 300 644 645 cell_1rw
* cell instance $24075 m0 *1 82.485,117.39
X$24075 299 600 300 644 645 cell_1rw
* cell instance $24076 r0 *1 82.485,117.39
X$24076 299 601 300 644 645 cell_1rw
* cell instance $24077 m0 *1 82.485,120.12
X$24077 299 602 300 644 645 cell_1rw
* cell instance $24078 r0 *1 82.485,120.12
X$24078 299 603 300 644 645 cell_1rw
* cell instance $24079 m0 *1 82.485,122.85
X$24079 299 604 300 644 645 cell_1rw
* cell instance $24080 r0 *1 82.485,122.85
X$24080 299 605 300 644 645 cell_1rw
* cell instance $24081 m0 *1 82.485,125.58
X$24081 299 606 300 644 645 cell_1rw
* cell instance $24082 r0 *1 82.485,125.58
X$24082 299 607 300 644 645 cell_1rw
* cell instance $24083 m0 *1 82.485,128.31
X$24083 299 609 300 644 645 cell_1rw
* cell instance $24084 r0 *1 82.485,128.31
X$24084 299 608 300 644 645 cell_1rw
* cell instance $24085 m0 *1 82.485,131.04
X$24085 299 610 300 644 645 cell_1rw
* cell instance $24086 r0 *1 82.485,131.04
X$24086 299 611 300 644 645 cell_1rw
* cell instance $24087 m0 *1 82.485,133.77
X$24087 299 612 300 644 645 cell_1rw
* cell instance $24088 r0 *1 82.485,133.77
X$24088 299 613 300 644 645 cell_1rw
* cell instance $24089 m0 *1 82.485,136.5
X$24089 299 615 300 644 645 cell_1rw
* cell instance $24090 r0 *1 82.485,136.5
X$24090 299 614 300 644 645 cell_1rw
* cell instance $24091 m0 *1 82.485,139.23
X$24091 299 617 300 644 645 cell_1rw
* cell instance $24092 r0 *1 82.485,139.23
X$24092 299 616 300 644 645 cell_1rw
* cell instance $24093 m0 *1 82.485,141.96
X$24093 299 618 300 644 645 cell_1rw
* cell instance $24094 r0 *1 82.485,141.96
X$24094 299 619 300 644 645 cell_1rw
* cell instance $24095 m0 *1 82.485,144.69
X$24095 299 620 300 644 645 cell_1rw
* cell instance $24096 r0 *1 82.485,144.69
X$24096 299 621 300 644 645 cell_1rw
* cell instance $24097 m0 *1 82.485,147.42
X$24097 299 622 300 644 645 cell_1rw
* cell instance $24098 r0 *1 82.485,147.42
X$24098 299 623 300 644 645 cell_1rw
* cell instance $24099 m0 *1 82.485,150.15
X$24099 299 624 300 644 645 cell_1rw
* cell instance $24100 r0 *1 82.485,150.15
X$24100 299 625 300 644 645 cell_1rw
* cell instance $24101 m0 *1 82.485,152.88
X$24101 299 626 300 644 645 cell_1rw
* cell instance $24102 r0 *1 82.485,152.88
X$24102 299 627 300 644 645 cell_1rw
* cell instance $24103 m0 *1 82.485,155.61
X$24103 299 628 300 644 645 cell_1rw
* cell instance $24104 r0 *1 82.485,155.61
X$24104 299 629 300 644 645 cell_1rw
* cell instance $24105 m0 *1 82.485,158.34
X$24105 299 630 300 644 645 cell_1rw
* cell instance $24106 r0 *1 82.485,158.34
X$24106 299 631 300 644 645 cell_1rw
* cell instance $24107 m0 *1 82.485,161.07
X$24107 299 632 300 644 645 cell_1rw
* cell instance $24108 r0 *1 82.485,161.07
X$24108 299 633 300 644 645 cell_1rw
* cell instance $24109 m0 *1 82.485,163.8
X$24109 299 634 300 644 645 cell_1rw
* cell instance $24110 r0 *1 82.485,163.8
X$24110 299 635 300 644 645 cell_1rw
* cell instance $24111 m0 *1 82.485,166.53
X$24111 299 637 300 644 645 cell_1rw
* cell instance $24112 r0 *1 82.485,166.53
X$24112 299 636 300 644 645 cell_1rw
* cell instance $24113 m0 *1 82.485,169.26
X$24113 299 639 300 644 645 cell_1rw
* cell instance $24114 r0 *1 82.485,169.26
X$24114 299 638 300 644 645 cell_1rw
* cell instance $24115 m0 *1 82.485,171.99
X$24115 299 640 300 644 645 cell_1rw
* cell instance $24116 r0 *1 82.485,171.99
X$24116 299 641 300 644 645 cell_1rw
* cell instance $24117 m0 *1 82.485,174.72
X$24117 299 642 300 644 645 cell_1rw
* cell instance $24118 r0 *1 82.485,174.72
X$24118 299 643 300 644 645 cell_1rw
* cell instance $24119 r0 *1 83.19,87.36
X$24119 301 322 302 644 645 cell_1rw
* cell instance $24120 m0 *1 83.19,90.09
X$24120 301 581 302 644 645 cell_1rw
* cell instance $24121 r0 *1 83.19,90.09
X$24121 301 580 302 644 645 cell_1rw
* cell instance $24122 m0 *1 83.19,92.82
X$24122 301 583 302 644 645 cell_1rw
* cell instance $24123 r0 *1 83.19,92.82
X$24123 301 582 302 644 645 cell_1rw
* cell instance $24124 m0 *1 83.19,95.55
X$24124 301 584 302 644 645 cell_1rw
* cell instance $24125 r0 *1 83.19,95.55
X$24125 301 585 302 644 645 cell_1rw
* cell instance $24126 m0 *1 83.19,98.28
X$24126 301 586 302 644 645 cell_1rw
* cell instance $24127 r0 *1 83.19,98.28
X$24127 301 587 302 644 645 cell_1rw
* cell instance $24128 m0 *1 83.19,101.01
X$24128 301 588 302 644 645 cell_1rw
* cell instance $24129 r0 *1 83.19,101.01
X$24129 301 589 302 644 645 cell_1rw
* cell instance $24130 m0 *1 83.19,103.74
X$24130 301 590 302 644 645 cell_1rw
* cell instance $24131 m0 *1 83.19,106.47
X$24131 301 593 302 644 645 cell_1rw
* cell instance $24132 r0 *1 83.19,103.74
X$24132 301 591 302 644 645 cell_1rw
* cell instance $24133 r0 *1 83.19,106.47
X$24133 301 592 302 644 645 cell_1rw
* cell instance $24134 m0 *1 83.19,109.2
X$24134 301 594 302 644 645 cell_1rw
* cell instance $24135 m0 *1 83.19,111.93
X$24135 301 597 302 644 645 cell_1rw
* cell instance $24136 r0 *1 83.19,109.2
X$24136 301 595 302 644 645 cell_1rw
* cell instance $24137 r0 *1 83.19,111.93
X$24137 301 596 302 644 645 cell_1rw
* cell instance $24138 m0 *1 83.19,114.66
X$24138 301 598 302 644 645 cell_1rw
* cell instance $24139 m0 *1 83.19,117.39
X$24139 301 600 302 644 645 cell_1rw
* cell instance $24140 r0 *1 83.19,114.66
X$24140 301 599 302 644 645 cell_1rw
* cell instance $24141 m0 *1 83.19,120.12
X$24141 301 602 302 644 645 cell_1rw
* cell instance $24142 r0 *1 83.19,117.39
X$24142 301 601 302 644 645 cell_1rw
* cell instance $24143 r0 *1 83.19,120.12
X$24143 301 603 302 644 645 cell_1rw
* cell instance $24144 m0 *1 83.19,122.85
X$24144 301 604 302 644 645 cell_1rw
* cell instance $24145 m0 *1 83.19,125.58
X$24145 301 606 302 644 645 cell_1rw
* cell instance $24146 r0 *1 83.19,122.85
X$24146 301 605 302 644 645 cell_1rw
* cell instance $24147 r0 *1 83.19,125.58
X$24147 301 607 302 644 645 cell_1rw
* cell instance $24148 m0 *1 83.19,128.31
X$24148 301 609 302 644 645 cell_1rw
* cell instance $24149 r0 *1 83.19,128.31
X$24149 301 608 302 644 645 cell_1rw
* cell instance $24150 m0 *1 83.19,131.04
X$24150 301 610 302 644 645 cell_1rw
* cell instance $24151 r0 *1 83.19,131.04
X$24151 301 611 302 644 645 cell_1rw
* cell instance $24152 m0 *1 83.19,133.77
X$24152 301 612 302 644 645 cell_1rw
* cell instance $24153 r0 *1 83.19,133.77
X$24153 301 613 302 644 645 cell_1rw
* cell instance $24154 m0 *1 83.19,136.5
X$24154 301 615 302 644 645 cell_1rw
* cell instance $24155 r0 *1 83.19,136.5
X$24155 301 614 302 644 645 cell_1rw
* cell instance $24156 m0 *1 83.19,139.23
X$24156 301 617 302 644 645 cell_1rw
* cell instance $24157 m0 *1 83.19,141.96
X$24157 301 618 302 644 645 cell_1rw
* cell instance $24158 r0 *1 83.19,139.23
X$24158 301 616 302 644 645 cell_1rw
* cell instance $24159 r0 *1 83.19,141.96
X$24159 301 619 302 644 645 cell_1rw
* cell instance $24160 m0 *1 83.19,144.69
X$24160 301 620 302 644 645 cell_1rw
* cell instance $24161 r0 *1 83.19,144.69
X$24161 301 621 302 644 645 cell_1rw
* cell instance $24162 m0 *1 83.19,147.42
X$24162 301 622 302 644 645 cell_1rw
* cell instance $24163 r0 *1 83.19,147.42
X$24163 301 623 302 644 645 cell_1rw
* cell instance $24164 m0 *1 83.19,150.15
X$24164 301 624 302 644 645 cell_1rw
* cell instance $24165 r0 *1 83.19,150.15
X$24165 301 625 302 644 645 cell_1rw
* cell instance $24166 m0 *1 83.19,152.88
X$24166 301 626 302 644 645 cell_1rw
* cell instance $24167 r0 *1 83.19,152.88
X$24167 301 627 302 644 645 cell_1rw
* cell instance $24168 m0 *1 83.19,155.61
X$24168 301 628 302 644 645 cell_1rw
* cell instance $24169 r0 *1 83.19,155.61
X$24169 301 629 302 644 645 cell_1rw
* cell instance $24170 m0 *1 83.19,158.34
X$24170 301 630 302 644 645 cell_1rw
* cell instance $24171 r0 *1 83.19,158.34
X$24171 301 631 302 644 645 cell_1rw
* cell instance $24172 m0 *1 83.19,161.07
X$24172 301 632 302 644 645 cell_1rw
* cell instance $24173 r0 *1 83.19,161.07
X$24173 301 633 302 644 645 cell_1rw
* cell instance $24174 m0 *1 83.19,163.8
X$24174 301 634 302 644 645 cell_1rw
* cell instance $24175 m0 *1 83.19,166.53
X$24175 301 637 302 644 645 cell_1rw
* cell instance $24176 r0 *1 83.19,163.8
X$24176 301 635 302 644 645 cell_1rw
* cell instance $24177 r0 *1 83.19,166.53
X$24177 301 636 302 644 645 cell_1rw
* cell instance $24178 m0 *1 83.19,169.26
X$24178 301 639 302 644 645 cell_1rw
* cell instance $24179 m0 *1 83.19,171.99
X$24179 301 640 302 644 645 cell_1rw
* cell instance $24180 r0 *1 83.19,169.26
X$24180 301 638 302 644 645 cell_1rw
* cell instance $24181 r0 *1 83.19,171.99
X$24181 301 641 302 644 645 cell_1rw
* cell instance $24182 m0 *1 83.19,174.72
X$24182 301 642 302 644 645 cell_1rw
* cell instance $24183 r0 *1 83.19,174.72
X$24183 301 643 302 644 645 cell_1rw
* cell instance $24184 r0 *1 83.895,87.36
X$24184 303 322 304 644 645 cell_1rw
* cell instance $24185 m0 *1 83.895,90.09
X$24185 303 581 304 644 645 cell_1rw
* cell instance $24186 r0 *1 83.895,90.09
X$24186 303 580 304 644 645 cell_1rw
* cell instance $24187 m0 *1 83.895,92.82
X$24187 303 583 304 644 645 cell_1rw
* cell instance $24188 r0 *1 83.895,92.82
X$24188 303 582 304 644 645 cell_1rw
* cell instance $24189 m0 *1 83.895,95.55
X$24189 303 584 304 644 645 cell_1rw
* cell instance $24190 r0 *1 83.895,95.55
X$24190 303 585 304 644 645 cell_1rw
* cell instance $24191 m0 *1 83.895,98.28
X$24191 303 586 304 644 645 cell_1rw
* cell instance $24192 r0 *1 83.895,98.28
X$24192 303 587 304 644 645 cell_1rw
* cell instance $24193 m0 *1 83.895,101.01
X$24193 303 588 304 644 645 cell_1rw
* cell instance $24194 r0 *1 83.895,101.01
X$24194 303 589 304 644 645 cell_1rw
* cell instance $24195 m0 *1 83.895,103.74
X$24195 303 590 304 644 645 cell_1rw
* cell instance $24196 r0 *1 83.895,103.74
X$24196 303 591 304 644 645 cell_1rw
* cell instance $24197 m0 *1 83.895,106.47
X$24197 303 593 304 644 645 cell_1rw
* cell instance $24198 r0 *1 83.895,106.47
X$24198 303 592 304 644 645 cell_1rw
* cell instance $24199 m0 *1 83.895,109.2
X$24199 303 594 304 644 645 cell_1rw
* cell instance $24200 m0 *1 83.895,111.93
X$24200 303 597 304 644 645 cell_1rw
* cell instance $24201 r0 *1 83.895,109.2
X$24201 303 595 304 644 645 cell_1rw
* cell instance $24202 m0 *1 83.895,114.66
X$24202 303 598 304 644 645 cell_1rw
* cell instance $24203 r0 *1 83.895,111.93
X$24203 303 596 304 644 645 cell_1rw
* cell instance $24204 r0 *1 83.895,114.66
X$24204 303 599 304 644 645 cell_1rw
* cell instance $24205 m0 *1 83.895,117.39
X$24205 303 600 304 644 645 cell_1rw
* cell instance $24206 r0 *1 83.895,117.39
X$24206 303 601 304 644 645 cell_1rw
* cell instance $24207 m0 *1 83.895,120.12
X$24207 303 602 304 644 645 cell_1rw
* cell instance $24208 r0 *1 83.895,120.12
X$24208 303 603 304 644 645 cell_1rw
* cell instance $24209 m0 *1 83.895,122.85
X$24209 303 604 304 644 645 cell_1rw
* cell instance $24210 m0 *1 83.895,125.58
X$24210 303 606 304 644 645 cell_1rw
* cell instance $24211 r0 *1 83.895,122.85
X$24211 303 605 304 644 645 cell_1rw
* cell instance $24212 r0 *1 83.895,125.58
X$24212 303 607 304 644 645 cell_1rw
* cell instance $24213 m0 *1 83.895,128.31
X$24213 303 609 304 644 645 cell_1rw
* cell instance $24214 r0 *1 83.895,128.31
X$24214 303 608 304 644 645 cell_1rw
* cell instance $24215 m0 *1 83.895,131.04
X$24215 303 610 304 644 645 cell_1rw
* cell instance $24216 r0 *1 83.895,131.04
X$24216 303 611 304 644 645 cell_1rw
* cell instance $24217 m0 *1 83.895,133.77
X$24217 303 612 304 644 645 cell_1rw
* cell instance $24218 r0 *1 83.895,133.77
X$24218 303 613 304 644 645 cell_1rw
* cell instance $24219 m0 *1 83.895,136.5
X$24219 303 615 304 644 645 cell_1rw
* cell instance $24220 m0 *1 83.895,139.23
X$24220 303 617 304 644 645 cell_1rw
* cell instance $24221 r0 *1 83.895,136.5
X$24221 303 614 304 644 645 cell_1rw
* cell instance $24222 r0 *1 83.895,139.23
X$24222 303 616 304 644 645 cell_1rw
* cell instance $24223 m0 *1 83.895,141.96
X$24223 303 618 304 644 645 cell_1rw
* cell instance $24224 r0 *1 83.895,141.96
X$24224 303 619 304 644 645 cell_1rw
* cell instance $24225 m0 *1 83.895,144.69
X$24225 303 620 304 644 645 cell_1rw
* cell instance $24226 r0 *1 83.895,144.69
X$24226 303 621 304 644 645 cell_1rw
* cell instance $24227 m0 *1 83.895,147.42
X$24227 303 622 304 644 645 cell_1rw
* cell instance $24228 r0 *1 83.895,147.42
X$24228 303 623 304 644 645 cell_1rw
* cell instance $24229 m0 *1 83.895,150.15
X$24229 303 624 304 644 645 cell_1rw
* cell instance $24230 r0 *1 83.895,150.15
X$24230 303 625 304 644 645 cell_1rw
* cell instance $24231 m0 *1 83.895,152.88
X$24231 303 626 304 644 645 cell_1rw
* cell instance $24232 r0 *1 83.895,152.88
X$24232 303 627 304 644 645 cell_1rw
* cell instance $24233 m0 *1 83.895,155.61
X$24233 303 628 304 644 645 cell_1rw
* cell instance $24234 r0 *1 83.895,155.61
X$24234 303 629 304 644 645 cell_1rw
* cell instance $24235 m0 *1 83.895,158.34
X$24235 303 630 304 644 645 cell_1rw
* cell instance $24236 r0 *1 83.895,158.34
X$24236 303 631 304 644 645 cell_1rw
* cell instance $24237 m0 *1 83.895,161.07
X$24237 303 632 304 644 645 cell_1rw
* cell instance $24238 r0 *1 83.895,161.07
X$24238 303 633 304 644 645 cell_1rw
* cell instance $24239 m0 *1 83.895,163.8
X$24239 303 634 304 644 645 cell_1rw
* cell instance $24240 r0 *1 83.895,163.8
X$24240 303 635 304 644 645 cell_1rw
* cell instance $24241 m0 *1 83.895,166.53
X$24241 303 637 304 644 645 cell_1rw
* cell instance $24242 r0 *1 83.895,166.53
X$24242 303 636 304 644 645 cell_1rw
* cell instance $24243 m0 *1 83.895,169.26
X$24243 303 639 304 644 645 cell_1rw
* cell instance $24244 m0 *1 83.895,171.99
X$24244 303 640 304 644 645 cell_1rw
* cell instance $24245 r0 *1 83.895,169.26
X$24245 303 638 304 644 645 cell_1rw
* cell instance $24246 r0 *1 83.895,171.99
X$24246 303 641 304 644 645 cell_1rw
* cell instance $24247 m0 *1 83.895,174.72
X$24247 303 642 304 644 645 cell_1rw
* cell instance $24248 r0 *1 83.895,174.72
X$24248 303 643 304 644 645 cell_1rw
* cell instance $24249 r0 *1 84.6,87.36
X$24249 305 322 306 644 645 cell_1rw
* cell instance $24250 m0 *1 84.6,90.09
X$24250 305 581 306 644 645 cell_1rw
* cell instance $24251 r0 *1 84.6,90.09
X$24251 305 580 306 644 645 cell_1rw
* cell instance $24252 m0 *1 84.6,92.82
X$24252 305 583 306 644 645 cell_1rw
* cell instance $24253 r0 *1 84.6,92.82
X$24253 305 582 306 644 645 cell_1rw
* cell instance $24254 m0 *1 84.6,95.55
X$24254 305 584 306 644 645 cell_1rw
* cell instance $24255 r0 *1 84.6,95.55
X$24255 305 585 306 644 645 cell_1rw
* cell instance $24256 m0 *1 84.6,98.28
X$24256 305 586 306 644 645 cell_1rw
* cell instance $24257 r0 *1 84.6,98.28
X$24257 305 587 306 644 645 cell_1rw
* cell instance $24258 m0 *1 84.6,101.01
X$24258 305 588 306 644 645 cell_1rw
* cell instance $24259 r0 *1 84.6,101.01
X$24259 305 589 306 644 645 cell_1rw
* cell instance $24260 m0 *1 84.6,103.74
X$24260 305 590 306 644 645 cell_1rw
* cell instance $24261 m0 *1 84.6,106.47
X$24261 305 593 306 644 645 cell_1rw
* cell instance $24262 r0 *1 84.6,103.74
X$24262 305 591 306 644 645 cell_1rw
* cell instance $24263 r0 *1 84.6,106.47
X$24263 305 592 306 644 645 cell_1rw
* cell instance $24264 m0 *1 84.6,109.2
X$24264 305 594 306 644 645 cell_1rw
* cell instance $24265 m0 *1 84.6,111.93
X$24265 305 597 306 644 645 cell_1rw
* cell instance $24266 r0 *1 84.6,109.2
X$24266 305 595 306 644 645 cell_1rw
* cell instance $24267 r0 *1 84.6,111.93
X$24267 305 596 306 644 645 cell_1rw
* cell instance $24268 m0 *1 84.6,114.66
X$24268 305 598 306 644 645 cell_1rw
* cell instance $24269 r0 *1 84.6,114.66
X$24269 305 599 306 644 645 cell_1rw
* cell instance $24270 m0 *1 84.6,117.39
X$24270 305 600 306 644 645 cell_1rw
* cell instance $24271 r0 *1 84.6,117.39
X$24271 305 601 306 644 645 cell_1rw
* cell instance $24272 m0 *1 84.6,120.12
X$24272 305 602 306 644 645 cell_1rw
* cell instance $24273 r0 *1 84.6,120.12
X$24273 305 603 306 644 645 cell_1rw
* cell instance $24274 m0 *1 84.6,122.85
X$24274 305 604 306 644 645 cell_1rw
* cell instance $24275 r0 *1 84.6,122.85
X$24275 305 605 306 644 645 cell_1rw
* cell instance $24276 m0 *1 84.6,125.58
X$24276 305 606 306 644 645 cell_1rw
* cell instance $24277 r0 *1 84.6,125.58
X$24277 305 607 306 644 645 cell_1rw
* cell instance $24278 m0 *1 84.6,128.31
X$24278 305 609 306 644 645 cell_1rw
* cell instance $24279 m0 *1 84.6,131.04
X$24279 305 610 306 644 645 cell_1rw
* cell instance $24280 r0 *1 84.6,128.31
X$24280 305 608 306 644 645 cell_1rw
* cell instance $24281 r0 *1 84.6,131.04
X$24281 305 611 306 644 645 cell_1rw
* cell instance $24282 m0 *1 84.6,133.77
X$24282 305 612 306 644 645 cell_1rw
* cell instance $24283 r0 *1 84.6,133.77
X$24283 305 613 306 644 645 cell_1rw
* cell instance $24284 m0 *1 84.6,136.5
X$24284 305 615 306 644 645 cell_1rw
* cell instance $24285 r0 *1 84.6,136.5
X$24285 305 614 306 644 645 cell_1rw
* cell instance $24286 m0 *1 84.6,139.23
X$24286 305 617 306 644 645 cell_1rw
* cell instance $24287 m0 *1 84.6,141.96
X$24287 305 618 306 644 645 cell_1rw
* cell instance $24288 r0 *1 84.6,139.23
X$24288 305 616 306 644 645 cell_1rw
* cell instance $24289 r0 *1 84.6,141.96
X$24289 305 619 306 644 645 cell_1rw
* cell instance $24290 m0 *1 84.6,144.69
X$24290 305 620 306 644 645 cell_1rw
* cell instance $24291 m0 *1 84.6,147.42
X$24291 305 622 306 644 645 cell_1rw
* cell instance $24292 r0 *1 84.6,144.69
X$24292 305 621 306 644 645 cell_1rw
* cell instance $24293 r0 *1 84.6,147.42
X$24293 305 623 306 644 645 cell_1rw
* cell instance $24294 m0 *1 84.6,150.15
X$24294 305 624 306 644 645 cell_1rw
* cell instance $24295 m0 *1 84.6,152.88
X$24295 305 626 306 644 645 cell_1rw
* cell instance $24296 r0 *1 84.6,150.15
X$24296 305 625 306 644 645 cell_1rw
* cell instance $24297 m0 *1 84.6,155.61
X$24297 305 628 306 644 645 cell_1rw
* cell instance $24298 r0 *1 84.6,152.88
X$24298 305 627 306 644 645 cell_1rw
* cell instance $24299 r0 *1 84.6,155.61
X$24299 305 629 306 644 645 cell_1rw
* cell instance $24300 m0 *1 84.6,158.34
X$24300 305 630 306 644 645 cell_1rw
* cell instance $24301 r0 *1 84.6,158.34
X$24301 305 631 306 644 645 cell_1rw
* cell instance $24302 m0 *1 84.6,161.07
X$24302 305 632 306 644 645 cell_1rw
* cell instance $24303 r0 *1 84.6,161.07
X$24303 305 633 306 644 645 cell_1rw
* cell instance $24304 m0 *1 84.6,163.8
X$24304 305 634 306 644 645 cell_1rw
* cell instance $24305 m0 *1 84.6,166.53
X$24305 305 637 306 644 645 cell_1rw
* cell instance $24306 r0 *1 84.6,163.8
X$24306 305 635 306 644 645 cell_1rw
* cell instance $24307 m0 *1 84.6,169.26
X$24307 305 639 306 644 645 cell_1rw
* cell instance $24308 r0 *1 84.6,166.53
X$24308 305 636 306 644 645 cell_1rw
* cell instance $24309 r0 *1 84.6,169.26
X$24309 305 638 306 644 645 cell_1rw
* cell instance $24310 m0 *1 84.6,171.99
X$24310 305 640 306 644 645 cell_1rw
* cell instance $24311 r0 *1 84.6,171.99
X$24311 305 641 306 644 645 cell_1rw
* cell instance $24312 m0 *1 84.6,174.72
X$24312 305 642 306 644 645 cell_1rw
* cell instance $24313 r0 *1 84.6,174.72
X$24313 305 643 306 644 645 cell_1rw
* cell instance $24314 r0 *1 85.305,87.36
X$24314 307 322 308 644 645 cell_1rw
* cell instance $24315 m0 *1 85.305,90.09
X$24315 307 581 308 644 645 cell_1rw
* cell instance $24316 r0 *1 85.305,90.09
X$24316 307 580 308 644 645 cell_1rw
* cell instance $24317 m0 *1 85.305,92.82
X$24317 307 583 308 644 645 cell_1rw
* cell instance $24318 r0 *1 85.305,92.82
X$24318 307 582 308 644 645 cell_1rw
* cell instance $24319 m0 *1 85.305,95.55
X$24319 307 584 308 644 645 cell_1rw
* cell instance $24320 r0 *1 85.305,95.55
X$24320 307 585 308 644 645 cell_1rw
* cell instance $24321 m0 *1 85.305,98.28
X$24321 307 586 308 644 645 cell_1rw
* cell instance $24322 m0 *1 85.305,101.01
X$24322 307 588 308 644 645 cell_1rw
* cell instance $24323 r0 *1 85.305,98.28
X$24323 307 587 308 644 645 cell_1rw
* cell instance $24324 r0 *1 85.305,101.01
X$24324 307 589 308 644 645 cell_1rw
* cell instance $24325 m0 *1 85.305,103.74
X$24325 307 590 308 644 645 cell_1rw
* cell instance $24326 r0 *1 85.305,103.74
X$24326 307 591 308 644 645 cell_1rw
* cell instance $24327 m0 *1 85.305,106.47
X$24327 307 593 308 644 645 cell_1rw
* cell instance $24328 r0 *1 85.305,106.47
X$24328 307 592 308 644 645 cell_1rw
* cell instance $24329 m0 *1 85.305,109.2
X$24329 307 594 308 644 645 cell_1rw
* cell instance $24330 r0 *1 85.305,109.2
X$24330 307 595 308 644 645 cell_1rw
* cell instance $24331 m0 *1 85.305,111.93
X$24331 307 597 308 644 645 cell_1rw
* cell instance $24332 r0 *1 85.305,111.93
X$24332 307 596 308 644 645 cell_1rw
* cell instance $24333 m0 *1 85.305,114.66
X$24333 307 598 308 644 645 cell_1rw
* cell instance $24334 r0 *1 85.305,114.66
X$24334 307 599 308 644 645 cell_1rw
* cell instance $24335 m0 *1 85.305,117.39
X$24335 307 600 308 644 645 cell_1rw
* cell instance $24336 m0 *1 85.305,120.12
X$24336 307 602 308 644 645 cell_1rw
* cell instance $24337 r0 *1 85.305,117.39
X$24337 307 601 308 644 645 cell_1rw
* cell instance $24338 r0 *1 85.305,120.12
X$24338 307 603 308 644 645 cell_1rw
* cell instance $24339 m0 *1 85.305,122.85
X$24339 307 604 308 644 645 cell_1rw
* cell instance $24340 r0 *1 85.305,122.85
X$24340 307 605 308 644 645 cell_1rw
* cell instance $24341 m0 *1 85.305,125.58
X$24341 307 606 308 644 645 cell_1rw
* cell instance $24342 m0 *1 85.305,128.31
X$24342 307 609 308 644 645 cell_1rw
* cell instance $24343 r0 *1 85.305,125.58
X$24343 307 607 308 644 645 cell_1rw
* cell instance $24344 r0 *1 85.305,128.31
X$24344 307 608 308 644 645 cell_1rw
* cell instance $24345 m0 *1 85.305,131.04
X$24345 307 610 308 644 645 cell_1rw
* cell instance $24346 m0 *1 85.305,133.77
X$24346 307 612 308 644 645 cell_1rw
* cell instance $24347 r0 *1 85.305,131.04
X$24347 307 611 308 644 645 cell_1rw
* cell instance $24348 r0 *1 85.305,133.77
X$24348 307 613 308 644 645 cell_1rw
* cell instance $24349 m0 *1 85.305,136.5
X$24349 307 615 308 644 645 cell_1rw
* cell instance $24350 r0 *1 85.305,136.5
X$24350 307 614 308 644 645 cell_1rw
* cell instance $24351 m0 *1 85.305,139.23
X$24351 307 617 308 644 645 cell_1rw
* cell instance $24352 r0 *1 85.305,139.23
X$24352 307 616 308 644 645 cell_1rw
* cell instance $24353 m0 *1 85.305,141.96
X$24353 307 618 308 644 645 cell_1rw
* cell instance $24354 m0 *1 85.305,144.69
X$24354 307 620 308 644 645 cell_1rw
* cell instance $24355 r0 *1 85.305,141.96
X$24355 307 619 308 644 645 cell_1rw
* cell instance $24356 r0 *1 85.305,144.69
X$24356 307 621 308 644 645 cell_1rw
* cell instance $24357 m0 *1 85.305,147.42
X$24357 307 622 308 644 645 cell_1rw
* cell instance $24358 r0 *1 85.305,147.42
X$24358 307 623 308 644 645 cell_1rw
* cell instance $24359 m0 *1 85.305,150.15
X$24359 307 624 308 644 645 cell_1rw
* cell instance $24360 r0 *1 85.305,150.15
X$24360 307 625 308 644 645 cell_1rw
* cell instance $24361 m0 *1 85.305,152.88
X$24361 307 626 308 644 645 cell_1rw
* cell instance $24362 r0 *1 85.305,152.88
X$24362 307 627 308 644 645 cell_1rw
* cell instance $24363 m0 *1 85.305,155.61
X$24363 307 628 308 644 645 cell_1rw
* cell instance $24364 r0 *1 85.305,155.61
X$24364 307 629 308 644 645 cell_1rw
* cell instance $24365 m0 *1 85.305,158.34
X$24365 307 630 308 644 645 cell_1rw
* cell instance $24366 m0 *1 85.305,161.07
X$24366 307 632 308 644 645 cell_1rw
* cell instance $24367 r0 *1 85.305,158.34
X$24367 307 631 308 644 645 cell_1rw
* cell instance $24368 r0 *1 85.305,161.07
X$24368 307 633 308 644 645 cell_1rw
* cell instance $24369 m0 *1 85.305,163.8
X$24369 307 634 308 644 645 cell_1rw
* cell instance $24370 r0 *1 85.305,163.8
X$24370 307 635 308 644 645 cell_1rw
* cell instance $24371 m0 *1 85.305,166.53
X$24371 307 637 308 644 645 cell_1rw
* cell instance $24372 m0 *1 85.305,169.26
X$24372 307 639 308 644 645 cell_1rw
* cell instance $24373 r0 *1 85.305,166.53
X$24373 307 636 308 644 645 cell_1rw
* cell instance $24374 r0 *1 85.305,169.26
X$24374 307 638 308 644 645 cell_1rw
* cell instance $24375 m0 *1 85.305,171.99
X$24375 307 640 308 644 645 cell_1rw
* cell instance $24376 m0 *1 85.305,174.72
X$24376 307 642 308 644 645 cell_1rw
* cell instance $24377 r0 *1 85.305,171.99
X$24377 307 641 308 644 645 cell_1rw
* cell instance $24378 r0 *1 85.305,174.72
X$24378 307 643 308 644 645 cell_1rw
* cell instance $24379 r0 *1 86.01,87.36
X$24379 309 322 310 644 645 cell_1rw
* cell instance $24380 m0 *1 86.01,90.09
X$24380 309 581 310 644 645 cell_1rw
* cell instance $24381 m0 *1 86.01,92.82
X$24381 309 583 310 644 645 cell_1rw
* cell instance $24382 r0 *1 86.01,90.09
X$24382 309 580 310 644 645 cell_1rw
* cell instance $24383 m0 *1 86.01,95.55
X$24383 309 584 310 644 645 cell_1rw
* cell instance $24384 r0 *1 86.01,92.82
X$24384 309 582 310 644 645 cell_1rw
* cell instance $24385 r0 *1 86.01,95.55
X$24385 309 585 310 644 645 cell_1rw
* cell instance $24386 m0 *1 86.01,98.28
X$24386 309 586 310 644 645 cell_1rw
* cell instance $24387 r0 *1 86.01,98.28
X$24387 309 587 310 644 645 cell_1rw
* cell instance $24388 m0 *1 86.01,101.01
X$24388 309 588 310 644 645 cell_1rw
* cell instance $24389 r0 *1 86.01,101.01
X$24389 309 589 310 644 645 cell_1rw
* cell instance $24390 m0 *1 86.01,103.74
X$24390 309 590 310 644 645 cell_1rw
* cell instance $24391 r0 *1 86.01,103.74
X$24391 309 591 310 644 645 cell_1rw
* cell instance $24392 m0 *1 86.01,106.47
X$24392 309 593 310 644 645 cell_1rw
* cell instance $24393 r0 *1 86.01,106.47
X$24393 309 592 310 644 645 cell_1rw
* cell instance $24394 m0 *1 86.01,109.2
X$24394 309 594 310 644 645 cell_1rw
* cell instance $24395 m0 *1 86.01,111.93
X$24395 309 597 310 644 645 cell_1rw
* cell instance $24396 r0 *1 86.01,109.2
X$24396 309 595 310 644 645 cell_1rw
* cell instance $24397 m0 *1 86.01,114.66
X$24397 309 598 310 644 645 cell_1rw
* cell instance $24398 r0 *1 86.01,111.93
X$24398 309 596 310 644 645 cell_1rw
* cell instance $24399 r0 *1 86.01,114.66
X$24399 309 599 310 644 645 cell_1rw
* cell instance $24400 m0 *1 86.01,117.39
X$24400 309 600 310 644 645 cell_1rw
* cell instance $24401 r0 *1 86.01,117.39
X$24401 309 601 310 644 645 cell_1rw
* cell instance $24402 m0 *1 86.01,120.12
X$24402 309 602 310 644 645 cell_1rw
* cell instance $24403 r0 *1 86.01,120.12
X$24403 309 603 310 644 645 cell_1rw
* cell instance $24404 m0 *1 86.01,122.85
X$24404 309 604 310 644 645 cell_1rw
* cell instance $24405 r0 *1 86.01,122.85
X$24405 309 605 310 644 645 cell_1rw
* cell instance $24406 m0 *1 86.01,125.58
X$24406 309 606 310 644 645 cell_1rw
* cell instance $24407 r0 *1 86.01,125.58
X$24407 309 607 310 644 645 cell_1rw
* cell instance $24408 m0 *1 86.01,128.31
X$24408 309 609 310 644 645 cell_1rw
* cell instance $24409 r0 *1 86.01,128.31
X$24409 309 608 310 644 645 cell_1rw
* cell instance $24410 m0 *1 86.01,131.04
X$24410 309 610 310 644 645 cell_1rw
* cell instance $24411 r0 *1 86.01,131.04
X$24411 309 611 310 644 645 cell_1rw
* cell instance $24412 m0 *1 86.01,133.77
X$24412 309 612 310 644 645 cell_1rw
* cell instance $24413 r0 *1 86.01,133.77
X$24413 309 613 310 644 645 cell_1rw
* cell instance $24414 m0 *1 86.01,136.5
X$24414 309 615 310 644 645 cell_1rw
* cell instance $24415 r0 *1 86.01,136.5
X$24415 309 614 310 644 645 cell_1rw
* cell instance $24416 m0 *1 86.01,139.23
X$24416 309 617 310 644 645 cell_1rw
* cell instance $24417 r0 *1 86.01,139.23
X$24417 309 616 310 644 645 cell_1rw
* cell instance $24418 m0 *1 86.01,141.96
X$24418 309 618 310 644 645 cell_1rw
* cell instance $24419 m0 *1 86.01,144.69
X$24419 309 620 310 644 645 cell_1rw
* cell instance $24420 r0 *1 86.01,141.96
X$24420 309 619 310 644 645 cell_1rw
* cell instance $24421 r0 *1 86.01,144.69
X$24421 309 621 310 644 645 cell_1rw
* cell instance $24422 m0 *1 86.01,147.42
X$24422 309 622 310 644 645 cell_1rw
* cell instance $24423 r0 *1 86.01,147.42
X$24423 309 623 310 644 645 cell_1rw
* cell instance $24424 m0 *1 86.01,150.15
X$24424 309 624 310 644 645 cell_1rw
* cell instance $24425 r0 *1 86.01,150.15
X$24425 309 625 310 644 645 cell_1rw
* cell instance $24426 m0 *1 86.01,152.88
X$24426 309 626 310 644 645 cell_1rw
* cell instance $24427 r0 *1 86.01,152.88
X$24427 309 627 310 644 645 cell_1rw
* cell instance $24428 m0 *1 86.01,155.61
X$24428 309 628 310 644 645 cell_1rw
* cell instance $24429 r0 *1 86.01,155.61
X$24429 309 629 310 644 645 cell_1rw
* cell instance $24430 m0 *1 86.01,158.34
X$24430 309 630 310 644 645 cell_1rw
* cell instance $24431 r0 *1 86.01,158.34
X$24431 309 631 310 644 645 cell_1rw
* cell instance $24432 m0 *1 86.01,161.07
X$24432 309 632 310 644 645 cell_1rw
* cell instance $24433 r0 *1 86.01,161.07
X$24433 309 633 310 644 645 cell_1rw
* cell instance $24434 m0 *1 86.01,163.8
X$24434 309 634 310 644 645 cell_1rw
* cell instance $24435 r0 *1 86.01,163.8
X$24435 309 635 310 644 645 cell_1rw
* cell instance $24436 m0 *1 86.01,166.53
X$24436 309 637 310 644 645 cell_1rw
* cell instance $24437 r0 *1 86.01,166.53
X$24437 309 636 310 644 645 cell_1rw
* cell instance $24438 m0 *1 86.01,169.26
X$24438 309 639 310 644 645 cell_1rw
* cell instance $24439 r0 *1 86.01,169.26
X$24439 309 638 310 644 645 cell_1rw
* cell instance $24440 m0 *1 86.01,171.99
X$24440 309 640 310 644 645 cell_1rw
* cell instance $24441 r0 *1 86.01,171.99
X$24441 309 641 310 644 645 cell_1rw
* cell instance $24442 m0 *1 86.01,174.72
X$24442 309 642 310 644 645 cell_1rw
* cell instance $24443 r0 *1 86.01,174.72
X$24443 309 643 310 644 645 cell_1rw
* cell instance $24444 r0 *1 86.715,87.36
X$24444 311 322 312 644 645 cell_1rw
* cell instance $24445 m0 *1 86.715,90.09
X$24445 311 581 312 644 645 cell_1rw
* cell instance $24446 r0 *1 86.715,90.09
X$24446 311 580 312 644 645 cell_1rw
* cell instance $24447 m0 *1 86.715,92.82
X$24447 311 583 312 644 645 cell_1rw
* cell instance $24448 r0 *1 86.715,92.82
X$24448 311 582 312 644 645 cell_1rw
* cell instance $24449 m0 *1 86.715,95.55
X$24449 311 584 312 644 645 cell_1rw
* cell instance $24450 m0 *1 86.715,98.28
X$24450 311 586 312 644 645 cell_1rw
* cell instance $24451 r0 *1 86.715,95.55
X$24451 311 585 312 644 645 cell_1rw
* cell instance $24452 r0 *1 86.715,98.28
X$24452 311 587 312 644 645 cell_1rw
* cell instance $24453 m0 *1 86.715,101.01
X$24453 311 588 312 644 645 cell_1rw
* cell instance $24454 m0 *1 86.715,103.74
X$24454 311 590 312 644 645 cell_1rw
* cell instance $24455 r0 *1 86.715,101.01
X$24455 311 589 312 644 645 cell_1rw
* cell instance $24456 r0 *1 86.715,103.74
X$24456 311 591 312 644 645 cell_1rw
* cell instance $24457 m0 *1 86.715,106.47
X$24457 311 593 312 644 645 cell_1rw
* cell instance $24458 r0 *1 86.715,106.47
X$24458 311 592 312 644 645 cell_1rw
* cell instance $24459 m0 *1 86.715,109.2
X$24459 311 594 312 644 645 cell_1rw
* cell instance $24460 r0 *1 86.715,109.2
X$24460 311 595 312 644 645 cell_1rw
* cell instance $24461 m0 *1 86.715,111.93
X$24461 311 597 312 644 645 cell_1rw
* cell instance $24462 r0 *1 86.715,111.93
X$24462 311 596 312 644 645 cell_1rw
* cell instance $24463 m0 *1 86.715,114.66
X$24463 311 598 312 644 645 cell_1rw
* cell instance $24464 r0 *1 86.715,114.66
X$24464 311 599 312 644 645 cell_1rw
* cell instance $24465 m0 *1 86.715,117.39
X$24465 311 600 312 644 645 cell_1rw
* cell instance $24466 r0 *1 86.715,117.39
X$24466 311 601 312 644 645 cell_1rw
* cell instance $24467 m0 *1 86.715,120.12
X$24467 311 602 312 644 645 cell_1rw
* cell instance $24468 r0 *1 86.715,120.12
X$24468 311 603 312 644 645 cell_1rw
* cell instance $24469 m0 *1 86.715,122.85
X$24469 311 604 312 644 645 cell_1rw
* cell instance $24470 r0 *1 86.715,122.85
X$24470 311 605 312 644 645 cell_1rw
* cell instance $24471 m0 *1 86.715,125.58
X$24471 311 606 312 644 645 cell_1rw
* cell instance $24472 r0 *1 86.715,125.58
X$24472 311 607 312 644 645 cell_1rw
* cell instance $24473 m0 *1 86.715,128.31
X$24473 311 609 312 644 645 cell_1rw
* cell instance $24474 r0 *1 86.715,128.31
X$24474 311 608 312 644 645 cell_1rw
* cell instance $24475 m0 *1 86.715,131.04
X$24475 311 610 312 644 645 cell_1rw
* cell instance $24476 r0 *1 86.715,131.04
X$24476 311 611 312 644 645 cell_1rw
* cell instance $24477 m0 *1 86.715,133.77
X$24477 311 612 312 644 645 cell_1rw
* cell instance $24478 r0 *1 86.715,133.77
X$24478 311 613 312 644 645 cell_1rw
* cell instance $24479 m0 *1 86.715,136.5
X$24479 311 615 312 644 645 cell_1rw
* cell instance $24480 r0 *1 86.715,136.5
X$24480 311 614 312 644 645 cell_1rw
* cell instance $24481 m0 *1 86.715,139.23
X$24481 311 617 312 644 645 cell_1rw
* cell instance $24482 r0 *1 86.715,139.23
X$24482 311 616 312 644 645 cell_1rw
* cell instance $24483 m0 *1 86.715,141.96
X$24483 311 618 312 644 645 cell_1rw
* cell instance $24484 m0 *1 86.715,144.69
X$24484 311 620 312 644 645 cell_1rw
* cell instance $24485 r0 *1 86.715,141.96
X$24485 311 619 312 644 645 cell_1rw
* cell instance $24486 r0 *1 86.715,144.69
X$24486 311 621 312 644 645 cell_1rw
* cell instance $24487 m0 *1 86.715,147.42
X$24487 311 622 312 644 645 cell_1rw
* cell instance $24488 r0 *1 86.715,147.42
X$24488 311 623 312 644 645 cell_1rw
* cell instance $24489 m0 *1 86.715,150.15
X$24489 311 624 312 644 645 cell_1rw
* cell instance $24490 r0 *1 86.715,150.15
X$24490 311 625 312 644 645 cell_1rw
* cell instance $24491 m0 *1 86.715,152.88
X$24491 311 626 312 644 645 cell_1rw
* cell instance $24492 r0 *1 86.715,152.88
X$24492 311 627 312 644 645 cell_1rw
* cell instance $24493 m0 *1 86.715,155.61
X$24493 311 628 312 644 645 cell_1rw
* cell instance $24494 r0 *1 86.715,155.61
X$24494 311 629 312 644 645 cell_1rw
* cell instance $24495 m0 *1 86.715,158.34
X$24495 311 630 312 644 645 cell_1rw
* cell instance $24496 r0 *1 86.715,158.34
X$24496 311 631 312 644 645 cell_1rw
* cell instance $24497 m0 *1 86.715,161.07
X$24497 311 632 312 644 645 cell_1rw
* cell instance $24498 r0 *1 86.715,161.07
X$24498 311 633 312 644 645 cell_1rw
* cell instance $24499 m0 *1 86.715,163.8
X$24499 311 634 312 644 645 cell_1rw
* cell instance $24500 r0 *1 86.715,163.8
X$24500 311 635 312 644 645 cell_1rw
* cell instance $24501 m0 *1 86.715,166.53
X$24501 311 637 312 644 645 cell_1rw
* cell instance $24502 m0 *1 86.715,169.26
X$24502 311 639 312 644 645 cell_1rw
* cell instance $24503 r0 *1 86.715,166.53
X$24503 311 636 312 644 645 cell_1rw
* cell instance $24504 m0 *1 86.715,171.99
X$24504 311 640 312 644 645 cell_1rw
* cell instance $24505 r0 *1 86.715,169.26
X$24505 311 638 312 644 645 cell_1rw
* cell instance $24506 r0 *1 86.715,171.99
X$24506 311 641 312 644 645 cell_1rw
* cell instance $24507 m0 *1 86.715,174.72
X$24507 311 642 312 644 645 cell_1rw
* cell instance $24508 r0 *1 86.715,174.72
X$24508 311 643 312 644 645 cell_1rw
* cell instance $24509 r0 *1 87.42,87.36
X$24509 313 322 314 644 645 cell_1rw
* cell instance $24510 m0 *1 87.42,90.09
X$24510 313 581 314 644 645 cell_1rw
* cell instance $24511 r0 *1 87.42,90.09
X$24511 313 580 314 644 645 cell_1rw
* cell instance $24512 m0 *1 87.42,92.82
X$24512 313 583 314 644 645 cell_1rw
* cell instance $24513 r0 *1 87.42,92.82
X$24513 313 582 314 644 645 cell_1rw
* cell instance $24514 m0 *1 87.42,95.55
X$24514 313 584 314 644 645 cell_1rw
* cell instance $24515 r0 *1 87.42,95.55
X$24515 313 585 314 644 645 cell_1rw
* cell instance $24516 m0 *1 87.42,98.28
X$24516 313 586 314 644 645 cell_1rw
* cell instance $24517 r0 *1 87.42,98.28
X$24517 313 587 314 644 645 cell_1rw
* cell instance $24518 m0 *1 87.42,101.01
X$24518 313 588 314 644 645 cell_1rw
* cell instance $24519 r0 *1 87.42,101.01
X$24519 313 589 314 644 645 cell_1rw
* cell instance $24520 m0 *1 87.42,103.74
X$24520 313 590 314 644 645 cell_1rw
* cell instance $24521 r0 *1 87.42,103.74
X$24521 313 591 314 644 645 cell_1rw
* cell instance $24522 m0 *1 87.42,106.47
X$24522 313 593 314 644 645 cell_1rw
* cell instance $24523 r0 *1 87.42,106.47
X$24523 313 592 314 644 645 cell_1rw
* cell instance $24524 m0 *1 87.42,109.2
X$24524 313 594 314 644 645 cell_1rw
* cell instance $24525 r0 *1 87.42,109.2
X$24525 313 595 314 644 645 cell_1rw
* cell instance $24526 m0 *1 87.42,111.93
X$24526 313 597 314 644 645 cell_1rw
* cell instance $24527 r0 *1 87.42,111.93
X$24527 313 596 314 644 645 cell_1rw
* cell instance $24528 m0 *1 87.42,114.66
X$24528 313 598 314 644 645 cell_1rw
* cell instance $24529 r0 *1 87.42,114.66
X$24529 313 599 314 644 645 cell_1rw
* cell instance $24530 m0 *1 87.42,117.39
X$24530 313 600 314 644 645 cell_1rw
* cell instance $24531 m0 *1 87.42,120.12
X$24531 313 602 314 644 645 cell_1rw
* cell instance $24532 r0 *1 87.42,117.39
X$24532 313 601 314 644 645 cell_1rw
* cell instance $24533 r0 *1 87.42,120.12
X$24533 313 603 314 644 645 cell_1rw
* cell instance $24534 m0 *1 87.42,122.85
X$24534 313 604 314 644 645 cell_1rw
* cell instance $24535 r0 *1 87.42,122.85
X$24535 313 605 314 644 645 cell_1rw
* cell instance $24536 m0 *1 87.42,125.58
X$24536 313 606 314 644 645 cell_1rw
* cell instance $24537 r0 *1 87.42,125.58
X$24537 313 607 314 644 645 cell_1rw
* cell instance $24538 m0 *1 87.42,128.31
X$24538 313 609 314 644 645 cell_1rw
* cell instance $24539 r0 *1 87.42,128.31
X$24539 313 608 314 644 645 cell_1rw
* cell instance $24540 m0 *1 87.42,131.04
X$24540 313 610 314 644 645 cell_1rw
* cell instance $24541 r0 *1 87.42,131.04
X$24541 313 611 314 644 645 cell_1rw
* cell instance $24542 m0 *1 87.42,133.77
X$24542 313 612 314 644 645 cell_1rw
* cell instance $24543 r0 *1 87.42,133.77
X$24543 313 613 314 644 645 cell_1rw
* cell instance $24544 m0 *1 87.42,136.5
X$24544 313 615 314 644 645 cell_1rw
* cell instance $24545 r0 *1 87.42,136.5
X$24545 313 614 314 644 645 cell_1rw
* cell instance $24546 m0 *1 87.42,139.23
X$24546 313 617 314 644 645 cell_1rw
* cell instance $24547 r0 *1 87.42,139.23
X$24547 313 616 314 644 645 cell_1rw
* cell instance $24548 m0 *1 87.42,141.96
X$24548 313 618 314 644 645 cell_1rw
* cell instance $24549 r0 *1 87.42,141.96
X$24549 313 619 314 644 645 cell_1rw
* cell instance $24550 m0 *1 87.42,144.69
X$24550 313 620 314 644 645 cell_1rw
* cell instance $24551 r0 *1 87.42,144.69
X$24551 313 621 314 644 645 cell_1rw
* cell instance $24552 m0 *1 87.42,147.42
X$24552 313 622 314 644 645 cell_1rw
* cell instance $24553 m0 *1 87.42,150.15
X$24553 313 624 314 644 645 cell_1rw
* cell instance $24554 r0 *1 87.42,147.42
X$24554 313 623 314 644 645 cell_1rw
* cell instance $24555 r0 *1 87.42,150.15
X$24555 313 625 314 644 645 cell_1rw
* cell instance $24556 m0 *1 87.42,152.88
X$24556 313 626 314 644 645 cell_1rw
* cell instance $24557 r0 *1 87.42,152.88
X$24557 313 627 314 644 645 cell_1rw
* cell instance $24558 m0 *1 87.42,155.61
X$24558 313 628 314 644 645 cell_1rw
* cell instance $24559 r0 *1 87.42,155.61
X$24559 313 629 314 644 645 cell_1rw
* cell instance $24560 m0 *1 87.42,158.34
X$24560 313 630 314 644 645 cell_1rw
* cell instance $24561 r0 *1 87.42,158.34
X$24561 313 631 314 644 645 cell_1rw
* cell instance $24562 m0 *1 87.42,161.07
X$24562 313 632 314 644 645 cell_1rw
* cell instance $24563 r0 *1 87.42,161.07
X$24563 313 633 314 644 645 cell_1rw
* cell instance $24564 m0 *1 87.42,163.8
X$24564 313 634 314 644 645 cell_1rw
* cell instance $24565 r0 *1 87.42,163.8
X$24565 313 635 314 644 645 cell_1rw
* cell instance $24566 m0 *1 87.42,166.53
X$24566 313 637 314 644 645 cell_1rw
* cell instance $24567 m0 *1 87.42,169.26
X$24567 313 639 314 644 645 cell_1rw
* cell instance $24568 r0 *1 87.42,166.53
X$24568 313 636 314 644 645 cell_1rw
* cell instance $24569 r0 *1 87.42,169.26
X$24569 313 638 314 644 645 cell_1rw
* cell instance $24570 m0 *1 87.42,171.99
X$24570 313 640 314 644 645 cell_1rw
* cell instance $24571 r0 *1 87.42,171.99
X$24571 313 641 314 644 645 cell_1rw
* cell instance $24572 m0 *1 87.42,174.72
X$24572 313 642 314 644 645 cell_1rw
* cell instance $24573 r0 *1 87.42,174.72
X$24573 313 643 314 644 645 cell_1rw
* cell instance $24574 m0 *1 88.125,90.09
X$24574 315 581 316 644 645 cell_1rw
* cell instance $24575 r0 *1 88.125,87.36
X$24575 315 322 316 644 645 cell_1rw
* cell instance $24576 r0 *1 88.125,90.09
X$24576 315 580 316 644 645 cell_1rw
* cell instance $24577 m0 *1 88.125,92.82
X$24577 315 583 316 644 645 cell_1rw
* cell instance $24578 r0 *1 88.125,92.82
X$24578 315 582 316 644 645 cell_1rw
* cell instance $24579 m0 *1 88.125,95.55
X$24579 315 584 316 644 645 cell_1rw
* cell instance $24580 m0 *1 88.125,98.28
X$24580 315 586 316 644 645 cell_1rw
* cell instance $24581 r0 *1 88.125,95.55
X$24581 315 585 316 644 645 cell_1rw
* cell instance $24582 r0 *1 88.125,98.28
X$24582 315 587 316 644 645 cell_1rw
* cell instance $24583 m0 *1 88.125,101.01
X$24583 315 588 316 644 645 cell_1rw
* cell instance $24584 r0 *1 88.125,101.01
X$24584 315 589 316 644 645 cell_1rw
* cell instance $24585 m0 *1 88.125,103.74
X$24585 315 590 316 644 645 cell_1rw
* cell instance $24586 r0 *1 88.125,103.74
X$24586 315 591 316 644 645 cell_1rw
* cell instance $24587 m0 *1 88.125,106.47
X$24587 315 593 316 644 645 cell_1rw
* cell instance $24588 r0 *1 88.125,106.47
X$24588 315 592 316 644 645 cell_1rw
* cell instance $24589 m0 *1 88.125,109.2
X$24589 315 594 316 644 645 cell_1rw
* cell instance $24590 r0 *1 88.125,109.2
X$24590 315 595 316 644 645 cell_1rw
* cell instance $24591 m0 *1 88.125,111.93
X$24591 315 597 316 644 645 cell_1rw
* cell instance $24592 r0 *1 88.125,111.93
X$24592 315 596 316 644 645 cell_1rw
* cell instance $24593 m0 *1 88.125,114.66
X$24593 315 598 316 644 645 cell_1rw
* cell instance $24594 r0 *1 88.125,114.66
X$24594 315 599 316 644 645 cell_1rw
* cell instance $24595 m0 *1 88.125,117.39
X$24595 315 600 316 644 645 cell_1rw
* cell instance $24596 r0 *1 88.125,117.39
X$24596 315 601 316 644 645 cell_1rw
* cell instance $24597 m0 *1 88.125,120.12
X$24597 315 602 316 644 645 cell_1rw
* cell instance $24598 m0 *1 88.125,122.85
X$24598 315 604 316 644 645 cell_1rw
* cell instance $24599 r0 *1 88.125,120.12
X$24599 315 603 316 644 645 cell_1rw
* cell instance $24600 r0 *1 88.125,122.85
X$24600 315 605 316 644 645 cell_1rw
* cell instance $24601 m0 *1 88.125,125.58
X$24601 315 606 316 644 645 cell_1rw
* cell instance $24602 m0 *1 88.125,128.31
X$24602 315 609 316 644 645 cell_1rw
* cell instance $24603 r0 *1 88.125,125.58
X$24603 315 607 316 644 645 cell_1rw
* cell instance $24604 m0 *1 88.125,131.04
X$24604 315 610 316 644 645 cell_1rw
* cell instance $24605 r0 *1 88.125,128.31
X$24605 315 608 316 644 645 cell_1rw
* cell instance $24606 r0 *1 88.125,131.04
X$24606 315 611 316 644 645 cell_1rw
* cell instance $24607 m0 *1 88.125,133.77
X$24607 315 612 316 644 645 cell_1rw
* cell instance $24608 m0 *1 88.125,136.5
X$24608 315 615 316 644 645 cell_1rw
* cell instance $24609 r0 *1 88.125,133.77
X$24609 315 613 316 644 645 cell_1rw
* cell instance $24610 r0 *1 88.125,136.5
X$24610 315 614 316 644 645 cell_1rw
* cell instance $24611 m0 *1 88.125,139.23
X$24611 315 617 316 644 645 cell_1rw
* cell instance $24612 r0 *1 88.125,139.23
X$24612 315 616 316 644 645 cell_1rw
* cell instance $24613 m0 *1 88.125,141.96
X$24613 315 618 316 644 645 cell_1rw
* cell instance $24614 r0 *1 88.125,141.96
X$24614 315 619 316 644 645 cell_1rw
* cell instance $24615 m0 *1 88.125,144.69
X$24615 315 620 316 644 645 cell_1rw
* cell instance $24616 r0 *1 88.125,144.69
X$24616 315 621 316 644 645 cell_1rw
* cell instance $24617 m0 *1 88.125,147.42
X$24617 315 622 316 644 645 cell_1rw
* cell instance $24618 m0 *1 88.125,150.15
X$24618 315 624 316 644 645 cell_1rw
* cell instance $24619 r0 *1 88.125,147.42
X$24619 315 623 316 644 645 cell_1rw
* cell instance $24620 r0 *1 88.125,150.15
X$24620 315 625 316 644 645 cell_1rw
* cell instance $24621 m0 *1 88.125,152.88
X$24621 315 626 316 644 645 cell_1rw
* cell instance $24622 r0 *1 88.125,152.88
X$24622 315 627 316 644 645 cell_1rw
* cell instance $24623 m0 *1 88.125,155.61
X$24623 315 628 316 644 645 cell_1rw
* cell instance $24624 m0 *1 88.125,158.34
X$24624 315 630 316 644 645 cell_1rw
* cell instance $24625 r0 *1 88.125,155.61
X$24625 315 629 316 644 645 cell_1rw
* cell instance $24626 m0 *1 88.125,161.07
X$24626 315 632 316 644 645 cell_1rw
* cell instance $24627 r0 *1 88.125,158.34
X$24627 315 631 316 644 645 cell_1rw
* cell instance $24628 r0 *1 88.125,161.07
X$24628 315 633 316 644 645 cell_1rw
* cell instance $24629 m0 *1 88.125,163.8
X$24629 315 634 316 644 645 cell_1rw
* cell instance $24630 r0 *1 88.125,163.8
X$24630 315 635 316 644 645 cell_1rw
* cell instance $24631 m0 *1 88.125,166.53
X$24631 315 637 316 644 645 cell_1rw
* cell instance $24632 r0 *1 88.125,166.53
X$24632 315 636 316 644 645 cell_1rw
* cell instance $24633 m0 *1 88.125,169.26
X$24633 315 639 316 644 645 cell_1rw
* cell instance $24634 r0 *1 88.125,169.26
X$24634 315 638 316 644 645 cell_1rw
* cell instance $24635 m0 *1 88.125,171.99
X$24635 315 640 316 644 645 cell_1rw
* cell instance $24636 m0 *1 88.125,174.72
X$24636 315 642 316 644 645 cell_1rw
* cell instance $24637 r0 *1 88.125,171.99
X$24637 315 641 316 644 645 cell_1rw
* cell instance $24638 r0 *1 88.125,174.72
X$24638 315 643 316 644 645 cell_1rw
* cell instance $24639 r0 *1 88.83,87.36
X$24639 317 322 318 644 645 cell_1rw
* cell instance $24640 m0 *1 88.83,90.09
X$24640 317 581 318 644 645 cell_1rw
* cell instance $24641 r0 *1 88.83,90.09
X$24641 317 580 318 644 645 cell_1rw
* cell instance $24642 m0 *1 88.83,92.82
X$24642 317 583 318 644 645 cell_1rw
* cell instance $24643 r0 *1 88.83,92.82
X$24643 317 582 318 644 645 cell_1rw
* cell instance $24644 m0 *1 88.83,95.55
X$24644 317 584 318 644 645 cell_1rw
* cell instance $24645 r0 *1 88.83,95.55
X$24645 317 585 318 644 645 cell_1rw
* cell instance $24646 m0 *1 88.83,98.28
X$24646 317 586 318 644 645 cell_1rw
* cell instance $24647 m0 *1 88.83,101.01
X$24647 317 588 318 644 645 cell_1rw
* cell instance $24648 r0 *1 88.83,98.28
X$24648 317 587 318 644 645 cell_1rw
* cell instance $24649 m0 *1 88.83,103.74
X$24649 317 590 318 644 645 cell_1rw
* cell instance $24650 r0 *1 88.83,101.01
X$24650 317 589 318 644 645 cell_1rw
* cell instance $24651 r0 *1 88.83,103.74
X$24651 317 591 318 644 645 cell_1rw
* cell instance $24652 m0 *1 88.83,106.47
X$24652 317 593 318 644 645 cell_1rw
* cell instance $24653 r0 *1 88.83,106.47
X$24653 317 592 318 644 645 cell_1rw
* cell instance $24654 m0 *1 88.83,109.2
X$24654 317 594 318 644 645 cell_1rw
* cell instance $24655 r0 *1 88.83,109.2
X$24655 317 595 318 644 645 cell_1rw
* cell instance $24656 m0 *1 88.83,111.93
X$24656 317 597 318 644 645 cell_1rw
* cell instance $24657 r0 *1 88.83,111.93
X$24657 317 596 318 644 645 cell_1rw
* cell instance $24658 m0 *1 88.83,114.66
X$24658 317 598 318 644 645 cell_1rw
* cell instance $24659 r0 *1 88.83,114.66
X$24659 317 599 318 644 645 cell_1rw
* cell instance $24660 m0 *1 88.83,117.39
X$24660 317 600 318 644 645 cell_1rw
* cell instance $24661 r0 *1 88.83,117.39
X$24661 317 601 318 644 645 cell_1rw
* cell instance $24662 m0 *1 88.83,120.12
X$24662 317 602 318 644 645 cell_1rw
* cell instance $24663 r0 *1 88.83,120.12
X$24663 317 603 318 644 645 cell_1rw
* cell instance $24664 m0 *1 88.83,122.85
X$24664 317 604 318 644 645 cell_1rw
* cell instance $24665 r0 *1 88.83,122.85
X$24665 317 605 318 644 645 cell_1rw
* cell instance $24666 m0 *1 88.83,125.58
X$24666 317 606 318 644 645 cell_1rw
* cell instance $24667 r0 *1 88.83,125.58
X$24667 317 607 318 644 645 cell_1rw
* cell instance $24668 m0 *1 88.83,128.31
X$24668 317 609 318 644 645 cell_1rw
* cell instance $24669 m0 *1 88.83,131.04
X$24669 317 610 318 644 645 cell_1rw
* cell instance $24670 r0 *1 88.83,128.31
X$24670 317 608 318 644 645 cell_1rw
* cell instance $24671 r0 *1 88.83,131.04
X$24671 317 611 318 644 645 cell_1rw
* cell instance $24672 m0 *1 88.83,133.77
X$24672 317 612 318 644 645 cell_1rw
* cell instance $24673 r0 *1 88.83,133.77
X$24673 317 613 318 644 645 cell_1rw
* cell instance $24674 m0 *1 88.83,136.5
X$24674 317 615 318 644 645 cell_1rw
* cell instance $24675 r0 *1 88.83,136.5
X$24675 317 614 318 644 645 cell_1rw
* cell instance $24676 m0 *1 88.83,139.23
X$24676 317 617 318 644 645 cell_1rw
* cell instance $24677 r0 *1 88.83,139.23
X$24677 317 616 318 644 645 cell_1rw
* cell instance $24678 m0 *1 88.83,141.96
X$24678 317 618 318 644 645 cell_1rw
* cell instance $24679 m0 *1 88.83,144.69
X$24679 317 620 318 644 645 cell_1rw
* cell instance $24680 r0 *1 88.83,141.96
X$24680 317 619 318 644 645 cell_1rw
* cell instance $24681 r0 *1 88.83,144.69
X$24681 317 621 318 644 645 cell_1rw
* cell instance $24682 m0 *1 88.83,147.42
X$24682 317 622 318 644 645 cell_1rw
* cell instance $24683 r0 *1 88.83,147.42
X$24683 317 623 318 644 645 cell_1rw
* cell instance $24684 m0 *1 88.83,150.15
X$24684 317 624 318 644 645 cell_1rw
* cell instance $24685 r0 *1 88.83,150.15
X$24685 317 625 318 644 645 cell_1rw
* cell instance $24686 m0 *1 88.83,152.88
X$24686 317 626 318 644 645 cell_1rw
* cell instance $24687 m0 *1 88.83,155.61
X$24687 317 628 318 644 645 cell_1rw
* cell instance $24688 r0 *1 88.83,152.88
X$24688 317 627 318 644 645 cell_1rw
* cell instance $24689 r0 *1 88.83,155.61
X$24689 317 629 318 644 645 cell_1rw
* cell instance $24690 m0 *1 88.83,158.34
X$24690 317 630 318 644 645 cell_1rw
* cell instance $24691 r0 *1 88.83,158.34
X$24691 317 631 318 644 645 cell_1rw
* cell instance $24692 m0 *1 88.83,161.07
X$24692 317 632 318 644 645 cell_1rw
* cell instance $24693 r0 *1 88.83,161.07
X$24693 317 633 318 644 645 cell_1rw
* cell instance $24694 m0 *1 88.83,163.8
X$24694 317 634 318 644 645 cell_1rw
* cell instance $24695 r0 *1 88.83,163.8
X$24695 317 635 318 644 645 cell_1rw
* cell instance $24696 m0 *1 88.83,166.53
X$24696 317 637 318 644 645 cell_1rw
* cell instance $24697 r0 *1 88.83,166.53
X$24697 317 636 318 644 645 cell_1rw
* cell instance $24698 m0 *1 88.83,169.26
X$24698 317 639 318 644 645 cell_1rw
* cell instance $24699 r0 *1 88.83,169.26
X$24699 317 638 318 644 645 cell_1rw
* cell instance $24700 m0 *1 88.83,171.99
X$24700 317 640 318 644 645 cell_1rw
* cell instance $24701 r0 *1 88.83,171.99
X$24701 317 641 318 644 645 cell_1rw
* cell instance $24702 m0 *1 88.83,174.72
X$24702 317 642 318 644 645 cell_1rw
* cell instance $24703 r0 *1 88.83,174.72
X$24703 317 643 318 644 645 cell_1rw
* cell instance $24704 r0 *1 89.535,87.36
X$24704 319 322 320 644 645 cell_1rw
* cell instance $24705 m0 *1 89.535,90.09
X$24705 319 581 320 644 645 cell_1rw
* cell instance $24706 r0 *1 89.535,90.09
X$24706 319 580 320 644 645 cell_1rw
* cell instance $24707 m0 *1 89.535,92.82
X$24707 319 583 320 644 645 cell_1rw
* cell instance $24708 r0 *1 89.535,92.82
X$24708 319 582 320 644 645 cell_1rw
* cell instance $24709 m0 *1 89.535,95.55
X$24709 319 584 320 644 645 cell_1rw
* cell instance $24710 r0 *1 89.535,95.55
X$24710 319 585 320 644 645 cell_1rw
* cell instance $24711 m0 *1 89.535,98.28
X$24711 319 586 320 644 645 cell_1rw
* cell instance $24712 r0 *1 89.535,98.28
X$24712 319 587 320 644 645 cell_1rw
* cell instance $24713 m0 *1 89.535,101.01
X$24713 319 588 320 644 645 cell_1rw
* cell instance $24714 m0 *1 89.535,103.74
X$24714 319 590 320 644 645 cell_1rw
* cell instance $24715 r0 *1 89.535,101.01
X$24715 319 589 320 644 645 cell_1rw
* cell instance $24716 r0 *1 89.535,103.74
X$24716 319 591 320 644 645 cell_1rw
* cell instance $24717 m0 *1 89.535,106.47
X$24717 319 593 320 644 645 cell_1rw
* cell instance $24718 r0 *1 89.535,106.47
X$24718 319 592 320 644 645 cell_1rw
* cell instance $24719 m0 *1 89.535,109.2
X$24719 319 594 320 644 645 cell_1rw
* cell instance $24720 r0 *1 89.535,109.2
X$24720 319 595 320 644 645 cell_1rw
* cell instance $24721 m0 *1 89.535,111.93
X$24721 319 597 320 644 645 cell_1rw
* cell instance $24722 r0 *1 89.535,111.93
X$24722 319 596 320 644 645 cell_1rw
* cell instance $24723 m0 *1 89.535,114.66
X$24723 319 598 320 644 645 cell_1rw
* cell instance $24724 r0 *1 89.535,114.66
X$24724 319 599 320 644 645 cell_1rw
* cell instance $24725 m0 *1 89.535,117.39
X$24725 319 600 320 644 645 cell_1rw
* cell instance $24726 m0 *1 89.535,120.12
X$24726 319 602 320 644 645 cell_1rw
* cell instance $24727 r0 *1 89.535,117.39
X$24727 319 601 320 644 645 cell_1rw
* cell instance $24728 r0 *1 89.535,120.12
X$24728 319 603 320 644 645 cell_1rw
* cell instance $24729 m0 *1 89.535,122.85
X$24729 319 604 320 644 645 cell_1rw
* cell instance $24730 r0 *1 89.535,122.85
X$24730 319 605 320 644 645 cell_1rw
* cell instance $24731 m0 *1 89.535,125.58
X$24731 319 606 320 644 645 cell_1rw
* cell instance $24732 m0 *1 89.535,128.31
X$24732 319 609 320 644 645 cell_1rw
* cell instance $24733 r0 *1 89.535,125.58
X$24733 319 607 320 644 645 cell_1rw
* cell instance $24734 r0 *1 89.535,128.31
X$24734 319 608 320 644 645 cell_1rw
* cell instance $24735 m0 *1 89.535,131.04
X$24735 319 610 320 644 645 cell_1rw
* cell instance $24736 r0 *1 89.535,131.04
X$24736 319 611 320 644 645 cell_1rw
* cell instance $24737 m0 *1 89.535,133.77
X$24737 319 612 320 644 645 cell_1rw
* cell instance $24738 m0 *1 89.535,136.5
X$24738 319 615 320 644 645 cell_1rw
* cell instance $24739 r0 *1 89.535,133.77
X$24739 319 613 320 644 645 cell_1rw
* cell instance $24740 r0 *1 89.535,136.5
X$24740 319 614 320 644 645 cell_1rw
* cell instance $24741 m0 *1 89.535,139.23
X$24741 319 617 320 644 645 cell_1rw
* cell instance $24742 m0 *1 89.535,141.96
X$24742 319 618 320 644 645 cell_1rw
* cell instance $24743 r0 *1 89.535,139.23
X$24743 319 616 320 644 645 cell_1rw
* cell instance $24744 r0 *1 89.535,141.96
X$24744 319 619 320 644 645 cell_1rw
* cell instance $24745 m0 *1 89.535,144.69
X$24745 319 620 320 644 645 cell_1rw
* cell instance $24746 m0 *1 89.535,147.42
X$24746 319 622 320 644 645 cell_1rw
* cell instance $24747 r0 *1 89.535,144.69
X$24747 319 621 320 644 645 cell_1rw
* cell instance $24748 r0 *1 89.535,147.42
X$24748 319 623 320 644 645 cell_1rw
* cell instance $24749 m0 *1 89.535,150.15
X$24749 319 624 320 644 645 cell_1rw
* cell instance $24750 r0 *1 89.535,150.15
X$24750 319 625 320 644 645 cell_1rw
* cell instance $24751 m0 *1 89.535,152.88
X$24751 319 626 320 644 645 cell_1rw
* cell instance $24752 r0 *1 89.535,152.88
X$24752 319 627 320 644 645 cell_1rw
* cell instance $24753 m0 *1 89.535,155.61
X$24753 319 628 320 644 645 cell_1rw
* cell instance $24754 r0 *1 89.535,155.61
X$24754 319 629 320 644 645 cell_1rw
* cell instance $24755 m0 *1 89.535,158.34
X$24755 319 630 320 644 645 cell_1rw
* cell instance $24756 r0 *1 89.535,158.34
X$24756 319 631 320 644 645 cell_1rw
* cell instance $24757 m0 *1 89.535,161.07
X$24757 319 632 320 644 645 cell_1rw
* cell instance $24758 r0 *1 89.535,161.07
X$24758 319 633 320 644 645 cell_1rw
* cell instance $24759 m0 *1 89.535,163.8
X$24759 319 634 320 644 645 cell_1rw
* cell instance $24760 r0 *1 89.535,163.8
X$24760 319 635 320 644 645 cell_1rw
* cell instance $24761 m0 *1 89.535,166.53
X$24761 319 637 320 644 645 cell_1rw
* cell instance $24762 r0 *1 89.535,166.53
X$24762 319 636 320 644 645 cell_1rw
* cell instance $24763 m0 *1 89.535,169.26
X$24763 319 639 320 644 645 cell_1rw
* cell instance $24764 r0 *1 89.535,169.26
X$24764 319 638 320 644 645 cell_1rw
* cell instance $24765 m0 *1 89.535,171.99
X$24765 319 640 320 644 645 cell_1rw
* cell instance $24766 r0 *1 89.535,171.99
X$24766 319 641 320 644 645 cell_1rw
* cell instance $24767 m0 *1 89.535,174.72
X$24767 319 642 320 644 645 cell_1rw
* cell instance $24768 r0 *1 89.535,174.72
X$24768 319 643 320 644 645 cell_1rw
* cell instance $24769 r0 *1 90.24,87.36
X$24769 321 322 323 644 645 cell_1rw
* cell instance $24770 m0 *1 90.24,90.09
X$24770 321 581 323 644 645 cell_1rw
* cell instance $24771 r0 *1 90.24,90.09
X$24771 321 580 323 644 645 cell_1rw
* cell instance $24772 m0 *1 90.24,92.82
X$24772 321 583 323 644 645 cell_1rw
* cell instance $24773 r0 *1 90.24,92.82
X$24773 321 582 323 644 645 cell_1rw
* cell instance $24774 m0 *1 90.24,95.55
X$24774 321 584 323 644 645 cell_1rw
* cell instance $24775 m0 *1 90.24,98.28
X$24775 321 586 323 644 645 cell_1rw
* cell instance $24776 r0 *1 90.24,95.55
X$24776 321 585 323 644 645 cell_1rw
* cell instance $24777 r0 *1 90.24,98.28
X$24777 321 587 323 644 645 cell_1rw
* cell instance $24778 m0 *1 90.24,101.01
X$24778 321 588 323 644 645 cell_1rw
* cell instance $24779 r0 *1 90.24,101.01
X$24779 321 589 323 644 645 cell_1rw
* cell instance $24780 m0 *1 90.24,103.74
X$24780 321 590 323 644 645 cell_1rw
* cell instance $24781 r0 *1 90.24,103.74
X$24781 321 591 323 644 645 cell_1rw
* cell instance $24782 m0 *1 90.24,106.47
X$24782 321 593 323 644 645 cell_1rw
* cell instance $24783 r0 *1 90.24,106.47
X$24783 321 592 323 644 645 cell_1rw
* cell instance $24784 m0 *1 90.24,109.2
X$24784 321 594 323 644 645 cell_1rw
* cell instance $24785 r0 *1 90.24,109.2
X$24785 321 595 323 644 645 cell_1rw
* cell instance $24786 m0 *1 90.24,111.93
X$24786 321 597 323 644 645 cell_1rw
* cell instance $24787 r0 *1 90.24,111.93
X$24787 321 596 323 644 645 cell_1rw
* cell instance $24788 m0 *1 90.24,114.66
X$24788 321 598 323 644 645 cell_1rw
* cell instance $24789 m0 *1 90.24,117.39
X$24789 321 600 323 644 645 cell_1rw
* cell instance $24790 r0 *1 90.24,114.66
X$24790 321 599 323 644 645 cell_1rw
* cell instance $24791 m0 *1 90.24,120.12
X$24791 321 602 323 644 645 cell_1rw
* cell instance $24792 r0 *1 90.24,117.39
X$24792 321 601 323 644 645 cell_1rw
* cell instance $24793 r0 *1 90.24,120.12
X$24793 321 603 323 644 645 cell_1rw
* cell instance $24794 m0 *1 90.24,122.85
X$24794 321 604 323 644 645 cell_1rw
* cell instance $24795 m0 *1 90.24,125.58
X$24795 321 606 323 644 645 cell_1rw
* cell instance $24796 r0 *1 90.24,122.85
X$24796 321 605 323 644 645 cell_1rw
* cell instance $24797 r0 *1 90.24,125.58
X$24797 321 607 323 644 645 cell_1rw
* cell instance $24798 m0 *1 90.24,128.31
X$24798 321 609 323 644 645 cell_1rw
* cell instance $24799 m0 *1 90.24,131.04
X$24799 321 610 323 644 645 cell_1rw
* cell instance $24800 r0 *1 90.24,128.31
X$24800 321 608 323 644 645 cell_1rw
* cell instance $24801 r0 *1 90.24,131.04
X$24801 321 611 323 644 645 cell_1rw
* cell instance $24802 m0 *1 90.24,133.77
X$24802 321 612 323 644 645 cell_1rw
* cell instance $24803 r0 *1 90.24,133.77
X$24803 321 613 323 644 645 cell_1rw
* cell instance $24804 m0 *1 90.24,136.5
X$24804 321 615 323 644 645 cell_1rw
* cell instance $24805 r0 *1 90.24,136.5
X$24805 321 614 323 644 645 cell_1rw
* cell instance $24806 m0 *1 90.24,139.23
X$24806 321 617 323 644 645 cell_1rw
* cell instance $24807 r0 *1 90.24,139.23
X$24807 321 616 323 644 645 cell_1rw
* cell instance $24808 m0 *1 90.24,141.96
X$24808 321 618 323 644 645 cell_1rw
* cell instance $24809 r0 *1 90.24,141.96
X$24809 321 619 323 644 645 cell_1rw
* cell instance $24810 m0 *1 90.24,144.69
X$24810 321 620 323 644 645 cell_1rw
* cell instance $24811 r0 *1 90.24,144.69
X$24811 321 621 323 644 645 cell_1rw
* cell instance $24812 m0 *1 90.24,147.42
X$24812 321 622 323 644 645 cell_1rw
* cell instance $24813 r0 *1 90.24,147.42
X$24813 321 623 323 644 645 cell_1rw
* cell instance $24814 m0 *1 90.24,150.15
X$24814 321 624 323 644 645 cell_1rw
* cell instance $24815 r0 *1 90.24,150.15
X$24815 321 625 323 644 645 cell_1rw
* cell instance $24816 m0 *1 90.24,152.88
X$24816 321 626 323 644 645 cell_1rw
* cell instance $24817 r0 *1 90.24,152.88
X$24817 321 627 323 644 645 cell_1rw
* cell instance $24818 m0 *1 90.24,155.61
X$24818 321 628 323 644 645 cell_1rw
* cell instance $24819 r0 *1 90.24,155.61
X$24819 321 629 323 644 645 cell_1rw
* cell instance $24820 m0 *1 90.24,158.34
X$24820 321 630 323 644 645 cell_1rw
* cell instance $24821 r0 *1 90.24,158.34
X$24821 321 631 323 644 645 cell_1rw
* cell instance $24822 m0 *1 90.24,161.07
X$24822 321 632 323 644 645 cell_1rw
* cell instance $24823 m0 *1 90.24,163.8
X$24823 321 634 323 644 645 cell_1rw
* cell instance $24824 r0 *1 90.24,161.07
X$24824 321 633 323 644 645 cell_1rw
* cell instance $24825 r0 *1 90.24,163.8
X$24825 321 635 323 644 645 cell_1rw
* cell instance $24826 m0 *1 90.24,166.53
X$24826 321 637 323 644 645 cell_1rw
* cell instance $24827 r0 *1 90.24,166.53
X$24827 321 636 323 644 645 cell_1rw
* cell instance $24828 m0 *1 90.24,169.26
X$24828 321 639 323 644 645 cell_1rw
* cell instance $24829 m0 *1 90.24,171.99
X$24829 321 640 323 644 645 cell_1rw
* cell instance $24830 r0 *1 90.24,169.26
X$24830 321 638 323 644 645 cell_1rw
* cell instance $24831 r0 *1 90.24,171.99
X$24831 321 641 323 644 645 cell_1rw
* cell instance $24832 m0 *1 90.24,174.72
X$24832 321 642 323 644 645 cell_1rw
* cell instance $24833 r0 *1 90.24,174.72
X$24833 321 643 323 644 645 cell_1rw
* cell instance $24834 r0 *1 90.945,87.36
X$24834 324 322 325 644 645 cell_1rw
* cell instance $24835 r0 *1 91.65,87.36
X$24835 326 322 327 644 645 cell_1rw
* cell instance $24836 r0 *1 92.355,87.36
X$24836 328 322 329 644 645 cell_1rw
* cell instance $24837 r0 *1 93.06,87.36
X$24837 330 322 331 644 645 cell_1rw
* cell instance $24838 r0 *1 93.765,87.36
X$24838 332 322 333 644 645 cell_1rw
* cell instance $24839 r0 *1 94.47,87.36
X$24839 334 322 335 644 645 cell_1rw
* cell instance $24840 r0 *1 95.175,87.36
X$24840 336 322 337 644 645 cell_1rw
* cell instance $24841 r0 *1 95.88,87.36
X$24841 338 322 339 644 645 cell_1rw
* cell instance $24842 r0 *1 96.585,87.36
X$24842 340 322 341 644 645 cell_1rw
* cell instance $24843 r0 *1 97.29,87.36
X$24843 342 322 343 644 645 cell_1rw
* cell instance $24844 r0 *1 97.995,87.36
X$24844 344 322 345 644 645 cell_1rw
* cell instance $24845 r0 *1 98.7,87.36
X$24845 346 322 347 644 645 cell_1rw
* cell instance $24846 r0 *1 99.405,87.36
X$24846 348 322 349 644 645 cell_1rw
* cell instance $24847 r0 *1 100.11,87.36
X$24847 350 322 351 644 645 cell_1rw
* cell instance $24848 r0 *1 100.815,87.36
X$24848 352 322 353 644 645 cell_1rw
* cell instance $24849 r0 *1 101.52,87.36
X$24849 354 322 355 644 645 cell_1rw
* cell instance $24850 r0 *1 102.225,87.36
X$24850 356 322 357 644 645 cell_1rw
* cell instance $24851 r0 *1 102.93,87.36
X$24851 358 322 359 644 645 cell_1rw
* cell instance $24852 r0 *1 103.635,87.36
X$24852 360 322 361 644 645 cell_1rw
* cell instance $24853 r0 *1 104.34,87.36
X$24853 362 322 363 644 645 cell_1rw
* cell instance $24854 r0 *1 105.045,87.36
X$24854 364 322 365 644 645 cell_1rw
* cell instance $24855 r0 *1 105.75,87.36
X$24855 366 322 367 644 645 cell_1rw
* cell instance $24856 r0 *1 106.455,87.36
X$24856 368 322 369 644 645 cell_1rw
* cell instance $24857 r0 *1 107.16,87.36
X$24857 370 322 371 644 645 cell_1rw
* cell instance $24858 r0 *1 107.865,87.36
X$24858 372 322 373 644 645 cell_1rw
* cell instance $24859 r0 *1 108.57,87.36
X$24859 374 322 375 644 645 cell_1rw
* cell instance $24860 r0 *1 109.275,87.36
X$24860 376 322 377 644 645 cell_1rw
* cell instance $24861 r0 *1 109.98,87.36
X$24861 378 322 379 644 645 cell_1rw
* cell instance $24862 r0 *1 110.685,87.36
X$24862 380 322 381 644 645 cell_1rw
* cell instance $24863 r0 *1 111.39,87.36
X$24863 382 322 383 644 645 cell_1rw
* cell instance $24864 r0 *1 112.095,87.36
X$24864 384 322 385 644 645 cell_1rw
* cell instance $24865 r0 *1 112.8,87.36
X$24865 386 322 387 644 645 cell_1rw
* cell instance $24866 r0 *1 113.505,87.36
X$24866 388 322 389 644 645 cell_1rw
* cell instance $24867 r0 *1 114.21,87.36
X$24867 390 322 391 644 645 cell_1rw
* cell instance $24868 r0 *1 114.915,87.36
X$24868 392 322 393 644 645 cell_1rw
* cell instance $24869 r0 *1 115.62,87.36
X$24869 394 322 395 644 645 cell_1rw
* cell instance $24870 r0 *1 116.325,87.36
X$24870 396 322 397 644 645 cell_1rw
* cell instance $24871 r0 *1 117.03,87.36
X$24871 398 322 399 644 645 cell_1rw
* cell instance $24872 r0 *1 117.735,87.36
X$24872 400 322 401 644 645 cell_1rw
* cell instance $24873 r0 *1 118.44,87.36
X$24873 402 322 403 644 645 cell_1rw
* cell instance $24874 r0 *1 119.145,87.36
X$24874 404 322 405 644 645 cell_1rw
* cell instance $24875 r0 *1 119.85,87.36
X$24875 406 322 407 644 645 cell_1rw
* cell instance $24876 r0 *1 120.555,87.36
X$24876 408 322 409 644 645 cell_1rw
* cell instance $24877 r0 *1 121.26,87.36
X$24877 410 322 411 644 645 cell_1rw
* cell instance $24878 r0 *1 121.965,87.36
X$24878 412 322 413 644 645 cell_1rw
* cell instance $24879 r0 *1 122.67,87.36
X$24879 414 322 415 644 645 cell_1rw
* cell instance $24880 r0 *1 123.375,87.36
X$24880 416 322 417 644 645 cell_1rw
* cell instance $24881 r0 *1 124.08,87.36
X$24881 418 322 419 644 645 cell_1rw
* cell instance $24882 r0 *1 124.785,87.36
X$24882 420 322 421 644 645 cell_1rw
* cell instance $24883 r0 *1 125.49,87.36
X$24883 422 322 423 644 645 cell_1rw
* cell instance $24884 r0 *1 126.195,87.36
X$24884 424 322 425 644 645 cell_1rw
* cell instance $24885 r0 *1 126.9,87.36
X$24885 426 322 427 644 645 cell_1rw
* cell instance $24886 r0 *1 127.605,87.36
X$24886 428 322 429 644 645 cell_1rw
* cell instance $24887 r0 *1 128.31,87.36
X$24887 430 322 431 644 645 cell_1rw
* cell instance $24888 r0 *1 129.015,87.36
X$24888 432 322 433 644 645 cell_1rw
* cell instance $24889 r0 *1 129.72,87.36
X$24889 434 322 435 644 645 cell_1rw
* cell instance $24890 r0 *1 130.425,87.36
X$24890 436 322 437 644 645 cell_1rw
* cell instance $24891 r0 *1 131.13,87.36
X$24891 438 322 439 644 645 cell_1rw
* cell instance $24892 r0 *1 131.835,87.36
X$24892 440 322 441 644 645 cell_1rw
* cell instance $24893 r0 *1 132.54,87.36
X$24893 442 322 443 644 645 cell_1rw
* cell instance $24894 r0 *1 133.245,87.36
X$24894 444 322 445 644 645 cell_1rw
* cell instance $24895 r0 *1 133.95,87.36
X$24895 446 322 447 644 645 cell_1rw
* cell instance $24896 r0 *1 134.655,87.36
X$24896 448 322 449 644 645 cell_1rw
* cell instance $24897 r0 *1 135.36,87.36
X$24897 450 322 451 644 645 cell_1rw
* cell instance $24898 r0 *1 136.065,87.36
X$24898 452 322 453 644 645 cell_1rw
* cell instance $24899 r0 *1 136.77,87.36
X$24899 454 322 455 644 645 cell_1rw
* cell instance $24900 r0 *1 137.475,87.36
X$24900 456 322 457 644 645 cell_1rw
* cell instance $24901 r0 *1 138.18,87.36
X$24901 458 322 459 644 645 cell_1rw
* cell instance $24902 r0 *1 138.885,87.36
X$24902 460 322 461 644 645 cell_1rw
* cell instance $24903 r0 *1 139.59,87.36
X$24903 462 322 463 644 645 cell_1rw
* cell instance $24904 r0 *1 140.295,87.36
X$24904 464 322 465 644 645 cell_1rw
* cell instance $24905 r0 *1 141,87.36
X$24905 466 322 467 644 645 cell_1rw
* cell instance $24906 r0 *1 141.705,87.36
X$24906 468 322 469 644 645 cell_1rw
* cell instance $24907 r0 *1 142.41,87.36
X$24907 470 322 471 644 645 cell_1rw
* cell instance $24908 r0 *1 143.115,87.36
X$24908 472 322 473 644 645 cell_1rw
* cell instance $24909 r0 *1 143.82,87.36
X$24909 474 322 475 644 645 cell_1rw
* cell instance $24910 r0 *1 144.525,87.36
X$24910 476 322 477 644 645 cell_1rw
* cell instance $24911 r0 *1 145.23,87.36
X$24911 478 322 479 644 645 cell_1rw
* cell instance $24912 r0 *1 145.935,87.36
X$24912 480 322 481 644 645 cell_1rw
* cell instance $24913 r0 *1 146.64,87.36
X$24913 482 322 483 644 645 cell_1rw
* cell instance $24914 r0 *1 147.345,87.36
X$24914 484 322 485 644 645 cell_1rw
* cell instance $24915 r0 *1 148.05,87.36
X$24915 486 322 487 644 645 cell_1rw
* cell instance $24916 r0 *1 148.755,87.36
X$24916 488 322 489 644 645 cell_1rw
* cell instance $24917 r0 *1 149.46,87.36
X$24917 490 322 491 644 645 cell_1rw
* cell instance $24918 r0 *1 150.165,87.36
X$24918 492 322 493 644 645 cell_1rw
* cell instance $24919 r0 *1 150.87,87.36
X$24919 494 322 495 644 645 cell_1rw
* cell instance $24920 r0 *1 151.575,87.36
X$24920 496 322 497 644 645 cell_1rw
* cell instance $24921 r0 *1 152.28,87.36
X$24921 498 322 499 644 645 cell_1rw
* cell instance $24922 r0 *1 152.985,87.36
X$24922 500 322 501 644 645 cell_1rw
* cell instance $24923 r0 *1 153.69,87.36
X$24923 502 322 503 644 645 cell_1rw
* cell instance $24924 r0 *1 154.395,87.36
X$24924 504 322 505 644 645 cell_1rw
* cell instance $24925 r0 *1 155.1,87.36
X$24925 506 322 507 644 645 cell_1rw
* cell instance $24926 r0 *1 155.805,87.36
X$24926 508 322 509 644 645 cell_1rw
* cell instance $24927 r0 *1 156.51,87.36
X$24927 510 322 511 644 645 cell_1rw
* cell instance $24928 r0 *1 157.215,87.36
X$24928 512 322 513 644 645 cell_1rw
* cell instance $24929 r0 *1 157.92,87.36
X$24929 514 322 515 644 645 cell_1rw
* cell instance $24930 r0 *1 158.625,87.36
X$24930 516 322 517 644 645 cell_1rw
* cell instance $24931 r0 *1 159.33,87.36
X$24931 518 322 519 644 645 cell_1rw
* cell instance $24932 r0 *1 160.035,87.36
X$24932 520 322 521 644 645 cell_1rw
* cell instance $24933 r0 *1 160.74,87.36
X$24933 522 322 523 644 645 cell_1rw
* cell instance $24934 r0 *1 161.445,87.36
X$24934 524 322 525 644 645 cell_1rw
* cell instance $24935 r0 *1 162.15,87.36
X$24935 526 322 527 644 645 cell_1rw
* cell instance $24936 r0 *1 162.855,87.36
X$24936 528 322 529 644 645 cell_1rw
* cell instance $24937 r0 *1 163.56,87.36
X$24937 530 322 531 644 645 cell_1rw
* cell instance $24938 r0 *1 164.265,87.36
X$24938 532 322 533 644 645 cell_1rw
* cell instance $24939 r0 *1 164.97,87.36
X$24939 534 322 535 644 645 cell_1rw
* cell instance $24940 r0 *1 165.675,87.36
X$24940 536 322 537 644 645 cell_1rw
* cell instance $24941 r0 *1 166.38,87.36
X$24941 538 322 539 644 645 cell_1rw
* cell instance $24942 r0 *1 167.085,87.36
X$24942 540 322 541 644 645 cell_1rw
* cell instance $24943 r0 *1 167.79,87.36
X$24943 542 322 543 644 645 cell_1rw
* cell instance $24944 r0 *1 168.495,87.36
X$24944 544 322 545 644 645 cell_1rw
* cell instance $24945 r0 *1 169.2,87.36
X$24945 546 322 547 644 645 cell_1rw
* cell instance $24946 r0 *1 169.905,87.36
X$24946 548 322 549 644 645 cell_1rw
* cell instance $24947 r0 *1 170.61,87.36
X$24947 550 322 551 644 645 cell_1rw
* cell instance $24948 r0 *1 171.315,87.36
X$24948 552 322 553 644 645 cell_1rw
* cell instance $24949 r0 *1 172.02,87.36
X$24949 554 322 555 644 645 cell_1rw
* cell instance $24950 r0 *1 172.725,87.36
X$24950 556 322 557 644 645 cell_1rw
* cell instance $24951 r0 *1 173.43,87.36
X$24951 558 322 559 644 645 cell_1rw
* cell instance $24952 r0 *1 174.135,87.36
X$24952 560 322 561 644 645 cell_1rw
* cell instance $24953 r0 *1 174.84,87.36
X$24953 562 322 563 644 645 cell_1rw
* cell instance $24954 r0 *1 175.545,87.36
X$24954 564 322 565 644 645 cell_1rw
* cell instance $24955 r0 *1 176.25,87.36
X$24955 566 322 567 644 645 cell_1rw
* cell instance $24956 r0 *1 176.955,87.36
X$24956 568 322 569 644 645 cell_1rw
* cell instance $24957 r0 *1 177.66,87.36
X$24957 570 322 571 644 645 cell_1rw
* cell instance $24958 r0 *1 178.365,87.36
X$24958 572 322 573 644 645 cell_1rw
* cell instance $24959 r0 *1 179.07,87.36
X$24959 574 322 575 644 645 cell_1rw
* cell instance $24960 r0 *1 179.775,87.36
X$24960 576 322 577 644 645 cell_1rw
* cell instance $24961 r0 *1 180.48,87.36
X$24961 578 322 579 644 645 cell_1rw
* cell instance $24962 m0 *1 90.945,90.09
X$24962 324 581 325 644 645 cell_1rw
* cell instance $24963 r0 *1 90.945,90.09
X$24963 324 580 325 644 645 cell_1rw
* cell instance $24964 m0 *1 90.945,92.82
X$24964 324 583 325 644 645 cell_1rw
* cell instance $24965 m0 *1 90.945,95.55
X$24965 324 584 325 644 645 cell_1rw
* cell instance $24966 r0 *1 90.945,92.82
X$24966 324 582 325 644 645 cell_1rw
* cell instance $24967 r0 *1 90.945,95.55
X$24967 324 585 325 644 645 cell_1rw
* cell instance $24968 m0 *1 90.945,98.28
X$24968 324 586 325 644 645 cell_1rw
* cell instance $24969 r0 *1 90.945,98.28
X$24969 324 587 325 644 645 cell_1rw
* cell instance $24970 m0 *1 90.945,101.01
X$24970 324 588 325 644 645 cell_1rw
* cell instance $24971 r0 *1 90.945,101.01
X$24971 324 589 325 644 645 cell_1rw
* cell instance $24972 m0 *1 90.945,103.74
X$24972 324 590 325 644 645 cell_1rw
* cell instance $24973 r0 *1 90.945,103.74
X$24973 324 591 325 644 645 cell_1rw
* cell instance $24974 m0 *1 90.945,106.47
X$24974 324 593 325 644 645 cell_1rw
* cell instance $24975 r0 *1 90.945,106.47
X$24975 324 592 325 644 645 cell_1rw
* cell instance $24976 m0 *1 90.945,109.2
X$24976 324 594 325 644 645 cell_1rw
* cell instance $24977 r0 *1 90.945,109.2
X$24977 324 595 325 644 645 cell_1rw
* cell instance $24978 m0 *1 90.945,111.93
X$24978 324 597 325 644 645 cell_1rw
* cell instance $24979 m0 *1 90.945,114.66
X$24979 324 598 325 644 645 cell_1rw
* cell instance $24980 r0 *1 90.945,111.93
X$24980 324 596 325 644 645 cell_1rw
* cell instance $24981 r0 *1 90.945,114.66
X$24981 324 599 325 644 645 cell_1rw
* cell instance $24982 m0 *1 90.945,117.39
X$24982 324 600 325 644 645 cell_1rw
* cell instance $24983 r0 *1 90.945,117.39
X$24983 324 601 325 644 645 cell_1rw
* cell instance $24984 m0 *1 90.945,120.12
X$24984 324 602 325 644 645 cell_1rw
* cell instance $24985 m0 *1 90.945,122.85
X$24985 324 604 325 644 645 cell_1rw
* cell instance $24986 r0 *1 90.945,120.12
X$24986 324 603 325 644 645 cell_1rw
* cell instance $24987 r0 *1 90.945,122.85
X$24987 324 605 325 644 645 cell_1rw
* cell instance $24988 m0 *1 90.945,125.58
X$24988 324 606 325 644 645 cell_1rw
* cell instance $24989 r0 *1 90.945,125.58
X$24989 324 607 325 644 645 cell_1rw
* cell instance $24990 m0 *1 90.945,128.31
X$24990 324 609 325 644 645 cell_1rw
* cell instance $24991 m0 *1 90.945,131.04
X$24991 324 610 325 644 645 cell_1rw
* cell instance $24992 r0 *1 90.945,128.31
X$24992 324 608 325 644 645 cell_1rw
* cell instance $24993 r0 *1 90.945,131.04
X$24993 324 611 325 644 645 cell_1rw
* cell instance $24994 m0 *1 90.945,133.77
X$24994 324 612 325 644 645 cell_1rw
* cell instance $24995 r0 *1 90.945,133.77
X$24995 324 613 325 644 645 cell_1rw
* cell instance $24996 m0 *1 90.945,136.5
X$24996 324 615 325 644 645 cell_1rw
* cell instance $24997 r0 *1 90.945,136.5
X$24997 324 614 325 644 645 cell_1rw
* cell instance $24998 m0 *1 90.945,139.23
X$24998 324 617 325 644 645 cell_1rw
* cell instance $24999 r0 *1 90.945,139.23
X$24999 324 616 325 644 645 cell_1rw
* cell instance $25000 m0 *1 90.945,141.96
X$25000 324 618 325 644 645 cell_1rw
* cell instance $25001 r0 *1 90.945,141.96
X$25001 324 619 325 644 645 cell_1rw
* cell instance $25002 m0 *1 90.945,144.69
X$25002 324 620 325 644 645 cell_1rw
* cell instance $25003 r0 *1 90.945,144.69
X$25003 324 621 325 644 645 cell_1rw
* cell instance $25004 m0 *1 90.945,147.42
X$25004 324 622 325 644 645 cell_1rw
* cell instance $25005 r0 *1 90.945,147.42
X$25005 324 623 325 644 645 cell_1rw
* cell instance $25006 m0 *1 90.945,150.15
X$25006 324 624 325 644 645 cell_1rw
* cell instance $25007 r0 *1 90.945,150.15
X$25007 324 625 325 644 645 cell_1rw
* cell instance $25008 m0 *1 90.945,152.88
X$25008 324 626 325 644 645 cell_1rw
* cell instance $25009 r0 *1 90.945,152.88
X$25009 324 627 325 644 645 cell_1rw
* cell instance $25010 m0 *1 90.945,155.61
X$25010 324 628 325 644 645 cell_1rw
* cell instance $25011 r0 *1 90.945,155.61
X$25011 324 629 325 644 645 cell_1rw
* cell instance $25012 m0 *1 90.945,158.34
X$25012 324 630 325 644 645 cell_1rw
* cell instance $25013 r0 *1 90.945,158.34
X$25013 324 631 325 644 645 cell_1rw
* cell instance $25014 m0 *1 90.945,161.07
X$25014 324 632 325 644 645 cell_1rw
* cell instance $25015 r0 *1 90.945,161.07
X$25015 324 633 325 644 645 cell_1rw
* cell instance $25016 m0 *1 90.945,163.8
X$25016 324 634 325 644 645 cell_1rw
* cell instance $25017 r0 *1 90.945,163.8
X$25017 324 635 325 644 645 cell_1rw
* cell instance $25018 m0 *1 90.945,166.53
X$25018 324 637 325 644 645 cell_1rw
* cell instance $25019 r0 *1 90.945,166.53
X$25019 324 636 325 644 645 cell_1rw
* cell instance $25020 m0 *1 90.945,169.26
X$25020 324 639 325 644 645 cell_1rw
* cell instance $25021 r0 *1 90.945,169.26
X$25021 324 638 325 644 645 cell_1rw
* cell instance $25022 m0 *1 90.945,171.99
X$25022 324 640 325 644 645 cell_1rw
* cell instance $25023 m0 *1 90.945,174.72
X$25023 324 642 325 644 645 cell_1rw
* cell instance $25024 r0 *1 90.945,171.99
X$25024 324 641 325 644 645 cell_1rw
* cell instance $25025 r0 *1 90.945,174.72
X$25025 324 643 325 644 645 cell_1rw
* cell instance $25026 m0 *1 91.65,90.09
X$25026 326 581 327 644 645 cell_1rw
* cell instance $25027 r0 *1 91.65,90.09
X$25027 326 580 327 644 645 cell_1rw
* cell instance $25028 m0 *1 91.65,92.82
X$25028 326 583 327 644 645 cell_1rw
* cell instance $25029 r0 *1 91.65,92.82
X$25029 326 582 327 644 645 cell_1rw
* cell instance $25030 m0 *1 91.65,95.55
X$25030 326 584 327 644 645 cell_1rw
* cell instance $25031 r0 *1 91.65,95.55
X$25031 326 585 327 644 645 cell_1rw
* cell instance $25032 m0 *1 91.65,98.28
X$25032 326 586 327 644 645 cell_1rw
* cell instance $25033 r0 *1 91.65,98.28
X$25033 326 587 327 644 645 cell_1rw
* cell instance $25034 m0 *1 91.65,101.01
X$25034 326 588 327 644 645 cell_1rw
* cell instance $25035 r0 *1 91.65,101.01
X$25035 326 589 327 644 645 cell_1rw
* cell instance $25036 m0 *1 91.65,103.74
X$25036 326 590 327 644 645 cell_1rw
* cell instance $25037 m0 *1 91.65,106.47
X$25037 326 593 327 644 645 cell_1rw
* cell instance $25038 r0 *1 91.65,103.74
X$25038 326 591 327 644 645 cell_1rw
* cell instance $25039 r0 *1 91.65,106.47
X$25039 326 592 327 644 645 cell_1rw
* cell instance $25040 m0 *1 91.65,109.2
X$25040 326 594 327 644 645 cell_1rw
* cell instance $25041 r0 *1 91.65,109.2
X$25041 326 595 327 644 645 cell_1rw
* cell instance $25042 m0 *1 91.65,111.93
X$25042 326 597 327 644 645 cell_1rw
* cell instance $25043 r0 *1 91.65,111.93
X$25043 326 596 327 644 645 cell_1rw
* cell instance $25044 m0 *1 91.65,114.66
X$25044 326 598 327 644 645 cell_1rw
* cell instance $25045 r0 *1 91.65,114.66
X$25045 326 599 327 644 645 cell_1rw
* cell instance $25046 m0 *1 91.65,117.39
X$25046 326 600 327 644 645 cell_1rw
* cell instance $25047 r0 *1 91.65,117.39
X$25047 326 601 327 644 645 cell_1rw
* cell instance $25048 m0 *1 91.65,120.12
X$25048 326 602 327 644 645 cell_1rw
* cell instance $25049 r0 *1 91.65,120.12
X$25049 326 603 327 644 645 cell_1rw
* cell instance $25050 m0 *1 91.65,122.85
X$25050 326 604 327 644 645 cell_1rw
* cell instance $25051 r0 *1 91.65,122.85
X$25051 326 605 327 644 645 cell_1rw
* cell instance $25052 m0 *1 91.65,125.58
X$25052 326 606 327 644 645 cell_1rw
* cell instance $25053 r0 *1 91.65,125.58
X$25053 326 607 327 644 645 cell_1rw
* cell instance $25054 m0 *1 91.65,128.31
X$25054 326 609 327 644 645 cell_1rw
* cell instance $25055 r0 *1 91.65,128.31
X$25055 326 608 327 644 645 cell_1rw
* cell instance $25056 m0 *1 91.65,131.04
X$25056 326 610 327 644 645 cell_1rw
* cell instance $25057 r0 *1 91.65,131.04
X$25057 326 611 327 644 645 cell_1rw
* cell instance $25058 m0 *1 91.65,133.77
X$25058 326 612 327 644 645 cell_1rw
* cell instance $25059 r0 *1 91.65,133.77
X$25059 326 613 327 644 645 cell_1rw
* cell instance $25060 m0 *1 91.65,136.5
X$25060 326 615 327 644 645 cell_1rw
* cell instance $25061 r0 *1 91.65,136.5
X$25061 326 614 327 644 645 cell_1rw
* cell instance $25062 m0 *1 91.65,139.23
X$25062 326 617 327 644 645 cell_1rw
* cell instance $25063 r0 *1 91.65,139.23
X$25063 326 616 327 644 645 cell_1rw
* cell instance $25064 m0 *1 91.65,141.96
X$25064 326 618 327 644 645 cell_1rw
* cell instance $25065 r0 *1 91.65,141.96
X$25065 326 619 327 644 645 cell_1rw
* cell instance $25066 m0 *1 91.65,144.69
X$25066 326 620 327 644 645 cell_1rw
* cell instance $25067 r0 *1 91.65,144.69
X$25067 326 621 327 644 645 cell_1rw
* cell instance $25068 m0 *1 91.65,147.42
X$25068 326 622 327 644 645 cell_1rw
* cell instance $25069 r0 *1 91.65,147.42
X$25069 326 623 327 644 645 cell_1rw
* cell instance $25070 m0 *1 91.65,150.15
X$25070 326 624 327 644 645 cell_1rw
* cell instance $25071 m0 *1 91.65,152.88
X$25071 326 626 327 644 645 cell_1rw
* cell instance $25072 r0 *1 91.65,150.15
X$25072 326 625 327 644 645 cell_1rw
* cell instance $25073 r0 *1 91.65,152.88
X$25073 326 627 327 644 645 cell_1rw
* cell instance $25074 m0 *1 91.65,155.61
X$25074 326 628 327 644 645 cell_1rw
* cell instance $25075 r0 *1 91.65,155.61
X$25075 326 629 327 644 645 cell_1rw
* cell instance $25076 m0 *1 91.65,158.34
X$25076 326 630 327 644 645 cell_1rw
* cell instance $25077 r0 *1 91.65,158.34
X$25077 326 631 327 644 645 cell_1rw
* cell instance $25078 m0 *1 91.65,161.07
X$25078 326 632 327 644 645 cell_1rw
* cell instance $25079 r0 *1 91.65,161.07
X$25079 326 633 327 644 645 cell_1rw
* cell instance $25080 m0 *1 91.65,163.8
X$25080 326 634 327 644 645 cell_1rw
* cell instance $25081 r0 *1 91.65,163.8
X$25081 326 635 327 644 645 cell_1rw
* cell instance $25082 m0 *1 91.65,166.53
X$25082 326 637 327 644 645 cell_1rw
* cell instance $25083 r0 *1 91.65,166.53
X$25083 326 636 327 644 645 cell_1rw
* cell instance $25084 m0 *1 91.65,169.26
X$25084 326 639 327 644 645 cell_1rw
* cell instance $25085 r0 *1 91.65,169.26
X$25085 326 638 327 644 645 cell_1rw
* cell instance $25086 m0 *1 91.65,171.99
X$25086 326 640 327 644 645 cell_1rw
* cell instance $25087 m0 *1 91.65,174.72
X$25087 326 642 327 644 645 cell_1rw
* cell instance $25088 r0 *1 91.65,171.99
X$25088 326 641 327 644 645 cell_1rw
* cell instance $25089 r0 *1 91.65,174.72
X$25089 326 643 327 644 645 cell_1rw
* cell instance $25090 m0 *1 92.355,90.09
X$25090 328 581 329 644 645 cell_1rw
* cell instance $25091 r0 *1 92.355,90.09
X$25091 328 580 329 644 645 cell_1rw
* cell instance $25092 m0 *1 92.355,92.82
X$25092 328 583 329 644 645 cell_1rw
* cell instance $25093 r0 *1 92.355,92.82
X$25093 328 582 329 644 645 cell_1rw
* cell instance $25094 m0 *1 92.355,95.55
X$25094 328 584 329 644 645 cell_1rw
* cell instance $25095 r0 *1 92.355,95.55
X$25095 328 585 329 644 645 cell_1rw
* cell instance $25096 m0 *1 92.355,98.28
X$25096 328 586 329 644 645 cell_1rw
* cell instance $25097 r0 *1 92.355,98.28
X$25097 328 587 329 644 645 cell_1rw
* cell instance $25098 m0 *1 92.355,101.01
X$25098 328 588 329 644 645 cell_1rw
* cell instance $25099 m0 *1 92.355,103.74
X$25099 328 590 329 644 645 cell_1rw
* cell instance $25100 r0 *1 92.355,101.01
X$25100 328 589 329 644 645 cell_1rw
* cell instance $25101 m0 *1 92.355,106.47
X$25101 328 593 329 644 645 cell_1rw
* cell instance $25102 r0 *1 92.355,103.74
X$25102 328 591 329 644 645 cell_1rw
* cell instance $25103 r0 *1 92.355,106.47
X$25103 328 592 329 644 645 cell_1rw
* cell instance $25104 m0 *1 92.355,109.2
X$25104 328 594 329 644 645 cell_1rw
* cell instance $25105 r0 *1 92.355,109.2
X$25105 328 595 329 644 645 cell_1rw
* cell instance $25106 m0 *1 92.355,111.93
X$25106 328 597 329 644 645 cell_1rw
* cell instance $25107 r0 *1 92.355,111.93
X$25107 328 596 329 644 645 cell_1rw
* cell instance $25108 m0 *1 92.355,114.66
X$25108 328 598 329 644 645 cell_1rw
* cell instance $25109 r0 *1 92.355,114.66
X$25109 328 599 329 644 645 cell_1rw
* cell instance $25110 m0 *1 92.355,117.39
X$25110 328 600 329 644 645 cell_1rw
* cell instance $25111 r0 *1 92.355,117.39
X$25111 328 601 329 644 645 cell_1rw
* cell instance $25112 m0 *1 92.355,120.12
X$25112 328 602 329 644 645 cell_1rw
* cell instance $25113 r0 *1 92.355,120.12
X$25113 328 603 329 644 645 cell_1rw
* cell instance $25114 m0 *1 92.355,122.85
X$25114 328 604 329 644 645 cell_1rw
* cell instance $25115 r0 *1 92.355,122.85
X$25115 328 605 329 644 645 cell_1rw
* cell instance $25116 m0 *1 92.355,125.58
X$25116 328 606 329 644 645 cell_1rw
* cell instance $25117 r0 *1 92.355,125.58
X$25117 328 607 329 644 645 cell_1rw
* cell instance $25118 m0 *1 92.355,128.31
X$25118 328 609 329 644 645 cell_1rw
* cell instance $25119 r0 *1 92.355,128.31
X$25119 328 608 329 644 645 cell_1rw
* cell instance $25120 m0 *1 92.355,131.04
X$25120 328 610 329 644 645 cell_1rw
* cell instance $25121 r0 *1 92.355,131.04
X$25121 328 611 329 644 645 cell_1rw
* cell instance $25122 m0 *1 92.355,133.77
X$25122 328 612 329 644 645 cell_1rw
* cell instance $25123 r0 *1 92.355,133.77
X$25123 328 613 329 644 645 cell_1rw
* cell instance $25124 m0 *1 92.355,136.5
X$25124 328 615 329 644 645 cell_1rw
* cell instance $25125 m0 *1 92.355,139.23
X$25125 328 617 329 644 645 cell_1rw
* cell instance $25126 r0 *1 92.355,136.5
X$25126 328 614 329 644 645 cell_1rw
* cell instance $25127 r0 *1 92.355,139.23
X$25127 328 616 329 644 645 cell_1rw
* cell instance $25128 m0 *1 92.355,141.96
X$25128 328 618 329 644 645 cell_1rw
* cell instance $25129 r0 *1 92.355,141.96
X$25129 328 619 329 644 645 cell_1rw
* cell instance $25130 m0 *1 92.355,144.69
X$25130 328 620 329 644 645 cell_1rw
* cell instance $25131 r0 *1 92.355,144.69
X$25131 328 621 329 644 645 cell_1rw
* cell instance $25132 m0 *1 92.355,147.42
X$25132 328 622 329 644 645 cell_1rw
* cell instance $25133 r0 *1 92.355,147.42
X$25133 328 623 329 644 645 cell_1rw
* cell instance $25134 m0 *1 92.355,150.15
X$25134 328 624 329 644 645 cell_1rw
* cell instance $25135 r0 *1 92.355,150.15
X$25135 328 625 329 644 645 cell_1rw
* cell instance $25136 m0 *1 92.355,152.88
X$25136 328 626 329 644 645 cell_1rw
* cell instance $25137 r0 *1 92.355,152.88
X$25137 328 627 329 644 645 cell_1rw
* cell instance $25138 m0 *1 92.355,155.61
X$25138 328 628 329 644 645 cell_1rw
* cell instance $25139 r0 *1 92.355,155.61
X$25139 328 629 329 644 645 cell_1rw
* cell instance $25140 m0 *1 92.355,158.34
X$25140 328 630 329 644 645 cell_1rw
* cell instance $25141 r0 *1 92.355,158.34
X$25141 328 631 329 644 645 cell_1rw
* cell instance $25142 m0 *1 92.355,161.07
X$25142 328 632 329 644 645 cell_1rw
* cell instance $25143 r0 *1 92.355,161.07
X$25143 328 633 329 644 645 cell_1rw
* cell instance $25144 m0 *1 92.355,163.8
X$25144 328 634 329 644 645 cell_1rw
* cell instance $25145 r0 *1 92.355,163.8
X$25145 328 635 329 644 645 cell_1rw
* cell instance $25146 m0 *1 92.355,166.53
X$25146 328 637 329 644 645 cell_1rw
* cell instance $25147 r0 *1 92.355,166.53
X$25147 328 636 329 644 645 cell_1rw
* cell instance $25148 m0 *1 92.355,169.26
X$25148 328 639 329 644 645 cell_1rw
* cell instance $25149 r0 *1 92.355,169.26
X$25149 328 638 329 644 645 cell_1rw
* cell instance $25150 m0 *1 92.355,171.99
X$25150 328 640 329 644 645 cell_1rw
* cell instance $25151 r0 *1 92.355,171.99
X$25151 328 641 329 644 645 cell_1rw
* cell instance $25152 m0 *1 92.355,174.72
X$25152 328 642 329 644 645 cell_1rw
* cell instance $25153 r0 *1 92.355,174.72
X$25153 328 643 329 644 645 cell_1rw
* cell instance $25154 m0 *1 93.06,90.09
X$25154 330 581 331 644 645 cell_1rw
* cell instance $25155 r0 *1 93.06,90.09
X$25155 330 580 331 644 645 cell_1rw
* cell instance $25156 m0 *1 93.06,92.82
X$25156 330 583 331 644 645 cell_1rw
* cell instance $25157 r0 *1 93.06,92.82
X$25157 330 582 331 644 645 cell_1rw
* cell instance $25158 m0 *1 93.06,95.55
X$25158 330 584 331 644 645 cell_1rw
* cell instance $25159 m0 *1 93.06,98.28
X$25159 330 586 331 644 645 cell_1rw
* cell instance $25160 r0 *1 93.06,95.55
X$25160 330 585 331 644 645 cell_1rw
* cell instance $25161 r0 *1 93.06,98.28
X$25161 330 587 331 644 645 cell_1rw
* cell instance $25162 m0 *1 93.06,101.01
X$25162 330 588 331 644 645 cell_1rw
* cell instance $25163 r0 *1 93.06,101.01
X$25163 330 589 331 644 645 cell_1rw
* cell instance $25164 m0 *1 93.06,103.74
X$25164 330 590 331 644 645 cell_1rw
* cell instance $25165 r0 *1 93.06,103.74
X$25165 330 591 331 644 645 cell_1rw
* cell instance $25166 m0 *1 93.06,106.47
X$25166 330 593 331 644 645 cell_1rw
* cell instance $25167 r0 *1 93.06,106.47
X$25167 330 592 331 644 645 cell_1rw
* cell instance $25168 m0 *1 93.06,109.2
X$25168 330 594 331 644 645 cell_1rw
* cell instance $25169 m0 *1 93.06,111.93
X$25169 330 597 331 644 645 cell_1rw
* cell instance $25170 r0 *1 93.06,109.2
X$25170 330 595 331 644 645 cell_1rw
* cell instance $25171 r0 *1 93.06,111.93
X$25171 330 596 331 644 645 cell_1rw
* cell instance $25172 m0 *1 93.06,114.66
X$25172 330 598 331 644 645 cell_1rw
* cell instance $25173 r0 *1 93.06,114.66
X$25173 330 599 331 644 645 cell_1rw
* cell instance $25174 m0 *1 93.06,117.39
X$25174 330 600 331 644 645 cell_1rw
* cell instance $25175 r0 *1 93.06,117.39
X$25175 330 601 331 644 645 cell_1rw
* cell instance $25176 m0 *1 93.06,120.12
X$25176 330 602 331 644 645 cell_1rw
* cell instance $25177 r0 *1 93.06,120.12
X$25177 330 603 331 644 645 cell_1rw
* cell instance $25178 m0 *1 93.06,122.85
X$25178 330 604 331 644 645 cell_1rw
* cell instance $25179 r0 *1 93.06,122.85
X$25179 330 605 331 644 645 cell_1rw
* cell instance $25180 m0 *1 93.06,125.58
X$25180 330 606 331 644 645 cell_1rw
* cell instance $25181 r0 *1 93.06,125.58
X$25181 330 607 331 644 645 cell_1rw
* cell instance $25182 m0 *1 93.06,128.31
X$25182 330 609 331 644 645 cell_1rw
* cell instance $25183 r0 *1 93.06,128.31
X$25183 330 608 331 644 645 cell_1rw
* cell instance $25184 m0 *1 93.06,131.04
X$25184 330 610 331 644 645 cell_1rw
* cell instance $25185 r0 *1 93.06,131.04
X$25185 330 611 331 644 645 cell_1rw
* cell instance $25186 m0 *1 93.06,133.77
X$25186 330 612 331 644 645 cell_1rw
* cell instance $25187 r0 *1 93.06,133.77
X$25187 330 613 331 644 645 cell_1rw
* cell instance $25188 m0 *1 93.06,136.5
X$25188 330 615 331 644 645 cell_1rw
* cell instance $25189 r0 *1 93.06,136.5
X$25189 330 614 331 644 645 cell_1rw
* cell instance $25190 m0 *1 93.06,139.23
X$25190 330 617 331 644 645 cell_1rw
* cell instance $25191 r0 *1 93.06,139.23
X$25191 330 616 331 644 645 cell_1rw
* cell instance $25192 m0 *1 93.06,141.96
X$25192 330 618 331 644 645 cell_1rw
* cell instance $25193 r0 *1 93.06,141.96
X$25193 330 619 331 644 645 cell_1rw
* cell instance $25194 m0 *1 93.06,144.69
X$25194 330 620 331 644 645 cell_1rw
* cell instance $25195 r0 *1 93.06,144.69
X$25195 330 621 331 644 645 cell_1rw
* cell instance $25196 m0 *1 93.06,147.42
X$25196 330 622 331 644 645 cell_1rw
* cell instance $25197 m0 *1 93.06,150.15
X$25197 330 624 331 644 645 cell_1rw
* cell instance $25198 r0 *1 93.06,147.42
X$25198 330 623 331 644 645 cell_1rw
* cell instance $25199 r0 *1 93.06,150.15
X$25199 330 625 331 644 645 cell_1rw
* cell instance $25200 m0 *1 93.06,152.88
X$25200 330 626 331 644 645 cell_1rw
* cell instance $25201 r0 *1 93.06,152.88
X$25201 330 627 331 644 645 cell_1rw
* cell instance $25202 m0 *1 93.06,155.61
X$25202 330 628 331 644 645 cell_1rw
* cell instance $25203 r0 *1 93.06,155.61
X$25203 330 629 331 644 645 cell_1rw
* cell instance $25204 m0 *1 93.06,158.34
X$25204 330 630 331 644 645 cell_1rw
* cell instance $25205 r0 *1 93.06,158.34
X$25205 330 631 331 644 645 cell_1rw
* cell instance $25206 m0 *1 93.06,161.07
X$25206 330 632 331 644 645 cell_1rw
* cell instance $25207 m0 *1 93.06,163.8
X$25207 330 634 331 644 645 cell_1rw
* cell instance $25208 r0 *1 93.06,161.07
X$25208 330 633 331 644 645 cell_1rw
* cell instance $25209 m0 *1 93.06,166.53
X$25209 330 637 331 644 645 cell_1rw
* cell instance $25210 r0 *1 93.06,163.8
X$25210 330 635 331 644 645 cell_1rw
* cell instance $25211 r0 *1 93.06,166.53
X$25211 330 636 331 644 645 cell_1rw
* cell instance $25212 m0 *1 93.06,169.26
X$25212 330 639 331 644 645 cell_1rw
* cell instance $25213 m0 *1 93.06,171.99
X$25213 330 640 331 644 645 cell_1rw
* cell instance $25214 r0 *1 93.06,169.26
X$25214 330 638 331 644 645 cell_1rw
* cell instance $25215 m0 *1 93.06,174.72
X$25215 330 642 331 644 645 cell_1rw
* cell instance $25216 r0 *1 93.06,171.99
X$25216 330 641 331 644 645 cell_1rw
* cell instance $25217 r0 *1 93.06,174.72
X$25217 330 643 331 644 645 cell_1rw
* cell instance $25218 m0 *1 93.765,90.09
X$25218 332 581 333 644 645 cell_1rw
* cell instance $25219 r0 *1 93.765,90.09
X$25219 332 580 333 644 645 cell_1rw
* cell instance $25220 m0 *1 93.765,92.82
X$25220 332 583 333 644 645 cell_1rw
* cell instance $25221 r0 *1 93.765,92.82
X$25221 332 582 333 644 645 cell_1rw
* cell instance $25222 m0 *1 93.765,95.55
X$25222 332 584 333 644 645 cell_1rw
* cell instance $25223 r0 *1 93.765,95.55
X$25223 332 585 333 644 645 cell_1rw
* cell instance $25224 m0 *1 93.765,98.28
X$25224 332 586 333 644 645 cell_1rw
* cell instance $25225 r0 *1 93.765,98.28
X$25225 332 587 333 644 645 cell_1rw
* cell instance $25226 m0 *1 93.765,101.01
X$25226 332 588 333 644 645 cell_1rw
* cell instance $25227 r0 *1 93.765,101.01
X$25227 332 589 333 644 645 cell_1rw
* cell instance $25228 m0 *1 93.765,103.74
X$25228 332 590 333 644 645 cell_1rw
* cell instance $25229 m0 *1 93.765,106.47
X$25229 332 593 333 644 645 cell_1rw
* cell instance $25230 r0 *1 93.765,103.74
X$25230 332 591 333 644 645 cell_1rw
* cell instance $25231 r0 *1 93.765,106.47
X$25231 332 592 333 644 645 cell_1rw
* cell instance $25232 m0 *1 93.765,109.2
X$25232 332 594 333 644 645 cell_1rw
* cell instance $25233 r0 *1 93.765,109.2
X$25233 332 595 333 644 645 cell_1rw
* cell instance $25234 m0 *1 93.765,111.93
X$25234 332 597 333 644 645 cell_1rw
* cell instance $25235 r0 *1 93.765,111.93
X$25235 332 596 333 644 645 cell_1rw
* cell instance $25236 m0 *1 93.765,114.66
X$25236 332 598 333 644 645 cell_1rw
* cell instance $25237 m0 *1 93.765,117.39
X$25237 332 600 333 644 645 cell_1rw
* cell instance $25238 r0 *1 93.765,114.66
X$25238 332 599 333 644 645 cell_1rw
* cell instance $25239 r0 *1 93.765,117.39
X$25239 332 601 333 644 645 cell_1rw
* cell instance $25240 m0 *1 93.765,120.12
X$25240 332 602 333 644 645 cell_1rw
* cell instance $25241 r0 *1 93.765,120.12
X$25241 332 603 333 644 645 cell_1rw
* cell instance $25242 m0 *1 93.765,122.85
X$25242 332 604 333 644 645 cell_1rw
* cell instance $25243 r0 *1 93.765,122.85
X$25243 332 605 333 644 645 cell_1rw
* cell instance $25244 m0 *1 93.765,125.58
X$25244 332 606 333 644 645 cell_1rw
* cell instance $25245 r0 *1 93.765,125.58
X$25245 332 607 333 644 645 cell_1rw
* cell instance $25246 m0 *1 93.765,128.31
X$25246 332 609 333 644 645 cell_1rw
* cell instance $25247 r0 *1 93.765,128.31
X$25247 332 608 333 644 645 cell_1rw
* cell instance $25248 m0 *1 93.765,131.04
X$25248 332 610 333 644 645 cell_1rw
* cell instance $25249 r0 *1 93.765,131.04
X$25249 332 611 333 644 645 cell_1rw
* cell instance $25250 m0 *1 93.765,133.77
X$25250 332 612 333 644 645 cell_1rw
* cell instance $25251 m0 *1 93.765,136.5
X$25251 332 615 333 644 645 cell_1rw
* cell instance $25252 r0 *1 93.765,133.77
X$25252 332 613 333 644 645 cell_1rw
* cell instance $25253 r0 *1 93.765,136.5
X$25253 332 614 333 644 645 cell_1rw
* cell instance $25254 m0 *1 93.765,139.23
X$25254 332 617 333 644 645 cell_1rw
* cell instance $25255 m0 *1 93.765,141.96
X$25255 332 618 333 644 645 cell_1rw
* cell instance $25256 r0 *1 93.765,139.23
X$25256 332 616 333 644 645 cell_1rw
* cell instance $25257 r0 *1 93.765,141.96
X$25257 332 619 333 644 645 cell_1rw
* cell instance $25258 m0 *1 93.765,144.69
X$25258 332 620 333 644 645 cell_1rw
* cell instance $25259 r0 *1 93.765,144.69
X$25259 332 621 333 644 645 cell_1rw
* cell instance $25260 m0 *1 93.765,147.42
X$25260 332 622 333 644 645 cell_1rw
* cell instance $25261 r0 *1 93.765,147.42
X$25261 332 623 333 644 645 cell_1rw
* cell instance $25262 m0 *1 93.765,150.15
X$25262 332 624 333 644 645 cell_1rw
* cell instance $25263 r0 *1 93.765,150.15
X$25263 332 625 333 644 645 cell_1rw
* cell instance $25264 m0 *1 93.765,152.88
X$25264 332 626 333 644 645 cell_1rw
* cell instance $25265 m0 *1 93.765,155.61
X$25265 332 628 333 644 645 cell_1rw
* cell instance $25266 r0 *1 93.765,152.88
X$25266 332 627 333 644 645 cell_1rw
* cell instance $25267 r0 *1 93.765,155.61
X$25267 332 629 333 644 645 cell_1rw
* cell instance $25268 m0 *1 93.765,158.34
X$25268 332 630 333 644 645 cell_1rw
* cell instance $25269 r0 *1 93.765,158.34
X$25269 332 631 333 644 645 cell_1rw
* cell instance $25270 m0 *1 93.765,161.07
X$25270 332 632 333 644 645 cell_1rw
* cell instance $25271 r0 *1 93.765,161.07
X$25271 332 633 333 644 645 cell_1rw
* cell instance $25272 m0 *1 93.765,163.8
X$25272 332 634 333 644 645 cell_1rw
* cell instance $25273 r0 *1 93.765,163.8
X$25273 332 635 333 644 645 cell_1rw
* cell instance $25274 m0 *1 93.765,166.53
X$25274 332 637 333 644 645 cell_1rw
* cell instance $25275 r0 *1 93.765,166.53
X$25275 332 636 333 644 645 cell_1rw
* cell instance $25276 m0 *1 93.765,169.26
X$25276 332 639 333 644 645 cell_1rw
* cell instance $25277 r0 *1 93.765,169.26
X$25277 332 638 333 644 645 cell_1rw
* cell instance $25278 m0 *1 93.765,171.99
X$25278 332 640 333 644 645 cell_1rw
* cell instance $25279 r0 *1 93.765,171.99
X$25279 332 641 333 644 645 cell_1rw
* cell instance $25280 m0 *1 93.765,174.72
X$25280 332 642 333 644 645 cell_1rw
* cell instance $25281 r0 *1 93.765,174.72
X$25281 332 643 333 644 645 cell_1rw
* cell instance $25282 m0 *1 94.47,90.09
X$25282 334 581 335 644 645 cell_1rw
* cell instance $25283 r0 *1 94.47,90.09
X$25283 334 580 335 644 645 cell_1rw
* cell instance $25284 m0 *1 94.47,92.82
X$25284 334 583 335 644 645 cell_1rw
* cell instance $25285 r0 *1 94.47,92.82
X$25285 334 582 335 644 645 cell_1rw
* cell instance $25286 m0 *1 94.47,95.55
X$25286 334 584 335 644 645 cell_1rw
* cell instance $25287 r0 *1 94.47,95.55
X$25287 334 585 335 644 645 cell_1rw
* cell instance $25288 m0 *1 94.47,98.28
X$25288 334 586 335 644 645 cell_1rw
* cell instance $25289 r0 *1 94.47,98.28
X$25289 334 587 335 644 645 cell_1rw
* cell instance $25290 m0 *1 94.47,101.01
X$25290 334 588 335 644 645 cell_1rw
* cell instance $25291 r0 *1 94.47,101.01
X$25291 334 589 335 644 645 cell_1rw
* cell instance $25292 m0 *1 94.47,103.74
X$25292 334 590 335 644 645 cell_1rw
* cell instance $25293 r0 *1 94.47,103.74
X$25293 334 591 335 644 645 cell_1rw
* cell instance $25294 m0 *1 94.47,106.47
X$25294 334 593 335 644 645 cell_1rw
* cell instance $25295 r0 *1 94.47,106.47
X$25295 334 592 335 644 645 cell_1rw
* cell instance $25296 m0 *1 94.47,109.2
X$25296 334 594 335 644 645 cell_1rw
* cell instance $25297 m0 *1 94.47,111.93
X$25297 334 597 335 644 645 cell_1rw
* cell instance $25298 r0 *1 94.47,109.2
X$25298 334 595 335 644 645 cell_1rw
* cell instance $25299 m0 *1 94.47,114.66
X$25299 334 598 335 644 645 cell_1rw
* cell instance $25300 r0 *1 94.47,111.93
X$25300 334 596 335 644 645 cell_1rw
* cell instance $25301 r0 *1 94.47,114.66
X$25301 334 599 335 644 645 cell_1rw
* cell instance $25302 m0 *1 94.47,117.39
X$25302 334 600 335 644 645 cell_1rw
* cell instance $25303 r0 *1 94.47,117.39
X$25303 334 601 335 644 645 cell_1rw
* cell instance $25304 m0 *1 94.47,120.12
X$25304 334 602 335 644 645 cell_1rw
* cell instance $25305 m0 *1 94.47,122.85
X$25305 334 604 335 644 645 cell_1rw
* cell instance $25306 r0 *1 94.47,120.12
X$25306 334 603 335 644 645 cell_1rw
* cell instance $25307 r0 *1 94.47,122.85
X$25307 334 605 335 644 645 cell_1rw
* cell instance $25308 m0 *1 94.47,125.58
X$25308 334 606 335 644 645 cell_1rw
* cell instance $25309 r0 *1 94.47,125.58
X$25309 334 607 335 644 645 cell_1rw
* cell instance $25310 m0 *1 94.47,128.31
X$25310 334 609 335 644 645 cell_1rw
* cell instance $25311 m0 *1 94.47,131.04
X$25311 334 610 335 644 645 cell_1rw
* cell instance $25312 r0 *1 94.47,128.31
X$25312 334 608 335 644 645 cell_1rw
* cell instance $25313 r0 *1 94.47,131.04
X$25313 334 611 335 644 645 cell_1rw
* cell instance $25314 m0 *1 94.47,133.77
X$25314 334 612 335 644 645 cell_1rw
* cell instance $25315 m0 *1 94.47,136.5
X$25315 334 615 335 644 645 cell_1rw
* cell instance $25316 r0 *1 94.47,133.77
X$25316 334 613 335 644 645 cell_1rw
* cell instance $25317 m0 *1 94.47,139.23
X$25317 334 617 335 644 645 cell_1rw
* cell instance $25318 r0 *1 94.47,136.5
X$25318 334 614 335 644 645 cell_1rw
* cell instance $25319 m0 *1 94.47,141.96
X$25319 334 618 335 644 645 cell_1rw
* cell instance $25320 r0 *1 94.47,139.23
X$25320 334 616 335 644 645 cell_1rw
* cell instance $25321 r0 *1 94.47,141.96
X$25321 334 619 335 644 645 cell_1rw
* cell instance $25322 m0 *1 94.47,144.69
X$25322 334 620 335 644 645 cell_1rw
* cell instance $25323 r0 *1 94.47,144.69
X$25323 334 621 335 644 645 cell_1rw
* cell instance $25324 m0 *1 94.47,147.42
X$25324 334 622 335 644 645 cell_1rw
* cell instance $25325 r0 *1 94.47,147.42
X$25325 334 623 335 644 645 cell_1rw
* cell instance $25326 m0 *1 94.47,150.15
X$25326 334 624 335 644 645 cell_1rw
* cell instance $25327 r0 *1 94.47,150.15
X$25327 334 625 335 644 645 cell_1rw
* cell instance $25328 m0 *1 94.47,152.88
X$25328 334 626 335 644 645 cell_1rw
* cell instance $25329 r0 *1 94.47,152.88
X$25329 334 627 335 644 645 cell_1rw
* cell instance $25330 m0 *1 94.47,155.61
X$25330 334 628 335 644 645 cell_1rw
* cell instance $25331 r0 *1 94.47,155.61
X$25331 334 629 335 644 645 cell_1rw
* cell instance $25332 m0 *1 94.47,158.34
X$25332 334 630 335 644 645 cell_1rw
* cell instance $25333 r0 *1 94.47,158.34
X$25333 334 631 335 644 645 cell_1rw
* cell instance $25334 m0 *1 94.47,161.07
X$25334 334 632 335 644 645 cell_1rw
* cell instance $25335 m0 *1 94.47,163.8
X$25335 334 634 335 644 645 cell_1rw
* cell instance $25336 r0 *1 94.47,161.07
X$25336 334 633 335 644 645 cell_1rw
* cell instance $25337 r0 *1 94.47,163.8
X$25337 334 635 335 644 645 cell_1rw
* cell instance $25338 m0 *1 94.47,166.53
X$25338 334 637 335 644 645 cell_1rw
* cell instance $25339 r0 *1 94.47,166.53
X$25339 334 636 335 644 645 cell_1rw
* cell instance $25340 m0 *1 94.47,169.26
X$25340 334 639 335 644 645 cell_1rw
* cell instance $25341 r0 *1 94.47,169.26
X$25341 334 638 335 644 645 cell_1rw
* cell instance $25342 m0 *1 94.47,171.99
X$25342 334 640 335 644 645 cell_1rw
* cell instance $25343 r0 *1 94.47,171.99
X$25343 334 641 335 644 645 cell_1rw
* cell instance $25344 m0 *1 94.47,174.72
X$25344 334 642 335 644 645 cell_1rw
* cell instance $25345 r0 *1 94.47,174.72
X$25345 334 643 335 644 645 cell_1rw
* cell instance $25346 m0 *1 95.175,90.09
X$25346 336 581 337 644 645 cell_1rw
* cell instance $25347 r0 *1 95.175,90.09
X$25347 336 580 337 644 645 cell_1rw
* cell instance $25348 m0 *1 95.175,92.82
X$25348 336 583 337 644 645 cell_1rw
* cell instance $25349 r0 *1 95.175,92.82
X$25349 336 582 337 644 645 cell_1rw
* cell instance $25350 m0 *1 95.175,95.55
X$25350 336 584 337 644 645 cell_1rw
* cell instance $25351 r0 *1 95.175,95.55
X$25351 336 585 337 644 645 cell_1rw
* cell instance $25352 m0 *1 95.175,98.28
X$25352 336 586 337 644 645 cell_1rw
* cell instance $25353 r0 *1 95.175,98.28
X$25353 336 587 337 644 645 cell_1rw
* cell instance $25354 m0 *1 95.175,101.01
X$25354 336 588 337 644 645 cell_1rw
* cell instance $25355 m0 *1 95.175,103.74
X$25355 336 590 337 644 645 cell_1rw
* cell instance $25356 r0 *1 95.175,101.01
X$25356 336 589 337 644 645 cell_1rw
* cell instance $25357 r0 *1 95.175,103.74
X$25357 336 591 337 644 645 cell_1rw
* cell instance $25358 m0 *1 95.175,106.47
X$25358 336 593 337 644 645 cell_1rw
* cell instance $25359 r0 *1 95.175,106.47
X$25359 336 592 337 644 645 cell_1rw
* cell instance $25360 m0 *1 95.175,109.2
X$25360 336 594 337 644 645 cell_1rw
* cell instance $25361 r0 *1 95.175,109.2
X$25361 336 595 337 644 645 cell_1rw
* cell instance $25362 m0 *1 95.175,111.93
X$25362 336 597 337 644 645 cell_1rw
* cell instance $25363 r0 *1 95.175,111.93
X$25363 336 596 337 644 645 cell_1rw
* cell instance $25364 m0 *1 95.175,114.66
X$25364 336 598 337 644 645 cell_1rw
* cell instance $25365 r0 *1 95.175,114.66
X$25365 336 599 337 644 645 cell_1rw
* cell instance $25366 m0 *1 95.175,117.39
X$25366 336 600 337 644 645 cell_1rw
* cell instance $25367 r0 *1 95.175,117.39
X$25367 336 601 337 644 645 cell_1rw
* cell instance $25368 m0 *1 95.175,120.12
X$25368 336 602 337 644 645 cell_1rw
* cell instance $25369 m0 *1 95.175,122.85
X$25369 336 604 337 644 645 cell_1rw
* cell instance $25370 r0 *1 95.175,120.12
X$25370 336 603 337 644 645 cell_1rw
* cell instance $25371 r0 *1 95.175,122.85
X$25371 336 605 337 644 645 cell_1rw
* cell instance $25372 m0 *1 95.175,125.58
X$25372 336 606 337 644 645 cell_1rw
* cell instance $25373 r0 *1 95.175,125.58
X$25373 336 607 337 644 645 cell_1rw
* cell instance $25374 m0 *1 95.175,128.31
X$25374 336 609 337 644 645 cell_1rw
* cell instance $25375 r0 *1 95.175,128.31
X$25375 336 608 337 644 645 cell_1rw
* cell instance $25376 m0 *1 95.175,131.04
X$25376 336 610 337 644 645 cell_1rw
* cell instance $25377 r0 *1 95.175,131.04
X$25377 336 611 337 644 645 cell_1rw
* cell instance $25378 m0 *1 95.175,133.77
X$25378 336 612 337 644 645 cell_1rw
* cell instance $25379 r0 *1 95.175,133.77
X$25379 336 613 337 644 645 cell_1rw
* cell instance $25380 m0 *1 95.175,136.5
X$25380 336 615 337 644 645 cell_1rw
* cell instance $25381 m0 *1 95.175,139.23
X$25381 336 617 337 644 645 cell_1rw
* cell instance $25382 r0 *1 95.175,136.5
X$25382 336 614 337 644 645 cell_1rw
* cell instance $25383 r0 *1 95.175,139.23
X$25383 336 616 337 644 645 cell_1rw
* cell instance $25384 m0 *1 95.175,141.96
X$25384 336 618 337 644 645 cell_1rw
* cell instance $25385 r0 *1 95.175,141.96
X$25385 336 619 337 644 645 cell_1rw
* cell instance $25386 m0 *1 95.175,144.69
X$25386 336 620 337 644 645 cell_1rw
* cell instance $25387 r0 *1 95.175,144.69
X$25387 336 621 337 644 645 cell_1rw
* cell instance $25388 m0 *1 95.175,147.42
X$25388 336 622 337 644 645 cell_1rw
* cell instance $25389 m0 *1 95.175,150.15
X$25389 336 624 337 644 645 cell_1rw
* cell instance $25390 r0 *1 95.175,147.42
X$25390 336 623 337 644 645 cell_1rw
* cell instance $25391 r0 *1 95.175,150.15
X$25391 336 625 337 644 645 cell_1rw
* cell instance $25392 m0 *1 95.175,152.88
X$25392 336 626 337 644 645 cell_1rw
* cell instance $25393 r0 *1 95.175,152.88
X$25393 336 627 337 644 645 cell_1rw
* cell instance $25394 m0 *1 95.175,155.61
X$25394 336 628 337 644 645 cell_1rw
* cell instance $25395 r0 *1 95.175,155.61
X$25395 336 629 337 644 645 cell_1rw
* cell instance $25396 m0 *1 95.175,158.34
X$25396 336 630 337 644 645 cell_1rw
* cell instance $25397 r0 *1 95.175,158.34
X$25397 336 631 337 644 645 cell_1rw
* cell instance $25398 m0 *1 95.175,161.07
X$25398 336 632 337 644 645 cell_1rw
* cell instance $25399 r0 *1 95.175,161.07
X$25399 336 633 337 644 645 cell_1rw
* cell instance $25400 m0 *1 95.175,163.8
X$25400 336 634 337 644 645 cell_1rw
* cell instance $25401 r0 *1 95.175,163.8
X$25401 336 635 337 644 645 cell_1rw
* cell instance $25402 m0 *1 95.175,166.53
X$25402 336 637 337 644 645 cell_1rw
* cell instance $25403 r0 *1 95.175,166.53
X$25403 336 636 337 644 645 cell_1rw
* cell instance $25404 m0 *1 95.175,169.26
X$25404 336 639 337 644 645 cell_1rw
* cell instance $25405 m0 *1 95.175,171.99
X$25405 336 640 337 644 645 cell_1rw
* cell instance $25406 r0 *1 95.175,169.26
X$25406 336 638 337 644 645 cell_1rw
* cell instance $25407 r0 *1 95.175,171.99
X$25407 336 641 337 644 645 cell_1rw
* cell instance $25408 m0 *1 95.175,174.72
X$25408 336 642 337 644 645 cell_1rw
* cell instance $25409 r0 *1 95.175,174.72
X$25409 336 643 337 644 645 cell_1rw
* cell instance $25410 m0 *1 95.88,90.09
X$25410 338 581 339 644 645 cell_1rw
* cell instance $25411 m0 *1 95.88,92.82
X$25411 338 583 339 644 645 cell_1rw
* cell instance $25412 r0 *1 95.88,90.09
X$25412 338 580 339 644 645 cell_1rw
* cell instance $25413 r0 *1 95.88,92.82
X$25413 338 582 339 644 645 cell_1rw
* cell instance $25414 m0 *1 95.88,95.55
X$25414 338 584 339 644 645 cell_1rw
* cell instance $25415 r0 *1 95.88,95.55
X$25415 338 585 339 644 645 cell_1rw
* cell instance $25416 m0 *1 95.88,98.28
X$25416 338 586 339 644 645 cell_1rw
* cell instance $25417 r0 *1 95.88,98.28
X$25417 338 587 339 644 645 cell_1rw
* cell instance $25418 m0 *1 95.88,101.01
X$25418 338 588 339 644 645 cell_1rw
* cell instance $25419 r0 *1 95.88,101.01
X$25419 338 589 339 644 645 cell_1rw
* cell instance $25420 m0 *1 95.88,103.74
X$25420 338 590 339 644 645 cell_1rw
* cell instance $25421 r0 *1 95.88,103.74
X$25421 338 591 339 644 645 cell_1rw
* cell instance $25422 m0 *1 95.88,106.47
X$25422 338 593 339 644 645 cell_1rw
* cell instance $25423 m0 *1 95.88,109.2
X$25423 338 594 339 644 645 cell_1rw
* cell instance $25424 r0 *1 95.88,106.47
X$25424 338 592 339 644 645 cell_1rw
* cell instance $25425 r0 *1 95.88,109.2
X$25425 338 595 339 644 645 cell_1rw
* cell instance $25426 m0 *1 95.88,111.93
X$25426 338 597 339 644 645 cell_1rw
* cell instance $25427 r0 *1 95.88,111.93
X$25427 338 596 339 644 645 cell_1rw
* cell instance $25428 m0 *1 95.88,114.66
X$25428 338 598 339 644 645 cell_1rw
* cell instance $25429 r0 *1 95.88,114.66
X$25429 338 599 339 644 645 cell_1rw
* cell instance $25430 m0 *1 95.88,117.39
X$25430 338 600 339 644 645 cell_1rw
* cell instance $25431 r0 *1 95.88,117.39
X$25431 338 601 339 644 645 cell_1rw
* cell instance $25432 m0 *1 95.88,120.12
X$25432 338 602 339 644 645 cell_1rw
* cell instance $25433 r0 *1 95.88,120.12
X$25433 338 603 339 644 645 cell_1rw
* cell instance $25434 m0 *1 95.88,122.85
X$25434 338 604 339 644 645 cell_1rw
* cell instance $25435 r0 *1 95.88,122.85
X$25435 338 605 339 644 645 cell_1rw
* cell instance $25436 m0 *1 95.88,125.58
X$25436 338 606 339 644 645 cell_1rw
* cell instance $25437 m0 *1 95.88,128.31
X$25437 338 609 339 644 645 cell_1rw
* cell instance $25438 r0 *1 95.88,125.58
X$25438 338 607 339 644 645 cell_1rw
* cell instance $25439 m0 *1 95.88,131.04
X$25439 338 610 339 644 645 cell_1rw
* cell instance $25440 r0 *1 95.88,128.31
X$25440 338 608 339 644 645 cell_1rw
* cell instance $25441 r0 *1 95.88,131.04
X$25441 338 611 339 644 645 cell_1rw
* cell instance $25442 m0 *1 95.88,133.77
X$25442 338 612 339 644 645 cell_1rw
* cell instance $25443 m0 *1 95.88,136.5
X$25443 338 615 339 644 645 cell_1rw
* cell instance $25444 r0 *1 95.88,133.77
X$25444 338 613 339 644 645 cell_1rw
* cell instance $25445 r0 *1 95.88,136.5
X$25445 338 614 339 644 645 cell_1rw
* cell instance $25446 m0 *1 95.88,139.23
X$25446 338 617 339 644 645 cell_1rw
* cell instance $25447 r0 *1 95.88,139.23
X$25447 338 616 339 644 645 cell_1rw
* cell instance $25448 m0 *1 95.88,141.96
X$25448 338 618 339 644 645 cell_1rw
* cell instance $25449 r0 *1 95.88,141.96
X$25449 338 619 339 644 645 cell_1rw
* cell instance $25450 m0 *1 95.88,144.69
X$25450 338 620 339 644 645 cell_1rw
* cell instance $25451 m0 *1 95.88,147.42
X$25451 338 622 339 644 645 cell_1rw
* cell instance $25452 r0 *1 95.88,144.69
X$25452 338 621 339 644 645 cell_1rw
* cell instance $25453 r0 *1 95.88,147.42
X$25453 338 623 339 644 645 cell_1rw
* cell instance $25454 m0 *1 95.88,150.15
X$25454 338 624 339 644 645 cell_1rw
* cell instance $25455 r0 *1 95.88,150.15
X$25455 338 625 339 644 645 cell_1rw
* cell instance $25456 m0 *1 95.88,152.88
X$25456 338 626 339 644 645 cell_1rw
* cell instance $25457 r0 *1 95.88,152.88
X$25457 338 627 339 644 645 cell_1rw
* cell instance $25458 m0 *1 95.88,155.61
X$25458 338 628 339 644 645 cell_1rw
* cell instance $25459 r0 *1 95.88,155.61
X$25459 338 629 339 644 645 cell_1rw
* cell instance $25460 m0 *1 95.88,158.34
X$25460 338 630 339 644 645 cell_1rw
* cell instance $25461 r0 *1 95.88,158.34
X$25461 338 631 339 644 645 cell_1rw
* cell instance $25462 m0 *1 95.88,161.07
X$25462 338 632 339 644 645 cell_1rw
* cell instance $25463 r0 *1 95.88,161.07
X$25463 338 633 339 644 645 cell_1rw
* cell instance $25464 m0 *1 95.88,163.8
X$25464 338 634 339 644 645 cell_1rw
* cell instance $25465 r0 *1 95.88,163.8
X$25465 338 635 339 644 645 cell_1rw
* cell instance $25466 m0 *1 95.88,166.53
X$25466 338 637 339 644 645 cell_1rw
* cell instance $25467 r0 *1 95.88,166.53
X$25467 338 636 339 644 645 cell_1rw
* cell instance $25468 m0 *1 95.88,169.26
X$25468 338 639 339 644 645 cell_1rw
* cell instance $25469 r0 *1 95.88,169.26
X$25469 338 638 339 644 645 cell_1rw
* cell instance $25470 m0 *1 95.88,171.99
X$25470 338 640 339 644 645 cell_1rw
* cell instance $25471 r0 *1 95.88,171.99
X$25471 338 641 339 644 645 cell_1rw
* cell instance $25472 m0 *1 95.88,174.72
X$25472 338 642 339 644 645 cell_1rw
* cell instance $25473 r0 *1 95.88,174.72
X$25473 338 643 339 644 645 cell_1rw
* cell instance $25474 m0 *1 96.585,90.09
X$25474 340 581 341 644 645 cell_1rw
* cell instance $25475 m0 *1 96.585,92.82
X$25475 340 583 341 644 645 cell_1rw
* cell instance $25476 r0 *1 96.585,90.09
X$25476 340 580 341 644 645 cell_1rw
* cell instance $25477 r0 *1 96.585,92.82
X$25477 340 582 341 644 645 cell_1rw
* cell instance $25478 m0 *1 96.585,95.55
X$25478 340 584 341 644 645 cell_1rw
* cell instance $25479 m0 *1 96.585,98.28
X$25479 340 586 341 644 645 cell_1rw
* cell instance $25480 r0 *1 96.585,95.55
X$25480 340 585 341 644 645 cell_1rw
* cell instance $25481 m0 *1 96.585,101.01
X$25481 340 588 341 644 645 cell_1rw
* cell instance $25482 r0 *1 96.585,98.28
X$25482 340 587 341 644 645 cell_1rw
* cell instance $25483 r0 *1 96.585,101.01
X$25483 340 589 341 644 645 cell_1rw
* cell instance $25484 m0 *1 96.585,103.74
X$25484 340 590 341 644 645 cell_1rw
* cell instance $25485 r0 *1 96.585,103.74
X$25485 340 591 341 644 645 cell_1rw
* cell instance $25486 m0 *1 96.585,106.47
X$25486 340 593 341 644 645 cell_1rw
* cell instance $25487 r0 *1 96.585,106.47
X$25487 340 592 341 644 645 cell_1rw
* cell instance $25488 m0 *1 96.585,109.2
X$25488 340 594 341 644 645 cell_1rw
* cell instance $25489 r0 *1 96.585,109.2
X$25489 340 595 341 644 645 cell_1rw
* cell instance $25490 m0 *1 96.585,111.93
X$25490 340 597 341 644 645 cell_1rw
* cell instance $25491 r0 *1 96.585,111.93
X$25491 340 596 341 644 645 cell_1rw
* cell instance $25492 m0 *1 96.585,114.66
X$25492 340 598 341 644 645 cell_1rw
* cell instance $25493 r0 *1 96.585,114.66
X$25493 340 599 341 644 645 cell_1rw
* cell instance $25494 m0 *1 96.585,117.39
X$25494 340 600 341 644 645 cell_1rw
* cell instance $25495 r0 *1 96.585,117.39
X$25495 340 601 341 644 645 cell_1rw
* cell instance $25496 m0 *1 96.585,120.12
X$25496 340 602 341 644 645 cell_1rw
* cell instance $25497 r0 *1 96.585,120.12
X$25497 340 603 341 644 645 cell_1rw
* cell instance $25498 m0 *1 96.585,122.85
X$25498 340 604 341 644 645 cell_1rw
* cell instance $25499 r0 *1 96.585,122.85
X$25499 340 605 341 644 645 cell_1rw
* cell instance $25500 m0 *1 96.585,125.58
X$25500 340 606 341 644 645 cell_1rw
* cell instance $25501 r0 *1 96.585,125.58
X$25501 340 607 341 644 645 cell_1rw
* cell instance $25502 m0 *1 96.585,128.31
X$25502 340 609 341 644 645 cell_1rw
* cell instance $25503 r0 *1 96.585,128.31
X$25503 340 608 341 644 645 cell_1rw
* cell instance $25504 m0 *1 96.585,131.04
X$25504 340 610 341 644 645 cell_1rw
* cell instance $25505 r0 *1 96.585,131.04
X$25505 340 611 341 644 645 cell_1rw
* cell instance $25506 m0 *1 96.585,133.77
X$25506 340 612 341 644 645 cell_1rw
* cell instance $25507 r0 *1 96.585,133.77
X$25507 340 613 341 644 645 cell_1rw
* cell instance $25508 m0 *1 96.585,136.5
X$25508 340 615 341 644 645 cell_1rw
* cell instance $25509 r0 *1 96.585,136.5
X$25509 340 614 341 644 645 cell_1rw
* cell instance $25510 m0 *1 96.585,139.23
X$25510 340 617 341 644 645 cell_1rw
* cell instance $25511 r0 *1 96.585,139.23
X$25511 340 616 341 644 645 cell_1rw
* cell instance $25512 m0 *1 96.585,141.96
X$25512 340 618 341 644 645 cell_1rw
* cell instance $25513 r0 *1 96.585,141.96
X$25513 340 619 341 644 645 cell_1rw
* cell instance $25514 m0 *1 96.585,144.69
X$25514 340 620 341 644 645 cell_1rw
* cell instance $25515 r0 *1 96.585,144.69
X$25515 340 621 341 644 645 cell_1rw
* cell instance $25516 m0 *1 96.585,147.42
X$25516 340 622 341 644 645 cell_1rw
* cell instance $25517 r0 *1 96.585,147.42
X$25517 340 623 341 644 645 cell_1rw
* cell instance $25518 m0 *1 96.585,150.15
X$25518 340 624 341 644 645 cell_1rw
* cell instance $25519 r0 *1 96.585,150.15
X$25519 340 625 341 644 645 cell_1rw
* cell instance $25520 m0 *1 96.585,152.88
X$25520 340 626 341 644 645 cell_1rw
* cell instance $25521 r0 *1 96.585,152.88
X$25521 340 627 341 644 645 cell_1rw
* cell instance $25522 m0 *1 96.585,155.61
X$25522 340 628 341 644 645 cell_1rw
* cell instance $25523 r0 *1 96.585,155.61
X$25523 340 629 341 644 645 cell_1rw
* cell instance $25524 m0 *1 96.585,158.34
X$25524 340 630 341 644 645 cell_1rw
* cell instance $25525 m0 *1 96.585,161.07
X$25525 340 632 341 644 645 cell_1rw
* cell instance $25526 r0 *1 96.585,158.34
X$25526 340 631 341 644 645 cell_1rw
* cell instance $25527 r0 *1 96.585,161.07
X$25527 340 633 341 644 645 cell_1rw
* cell instance $25528 m0 *1 96.585,163.8
X$25528 340 634 341 644 645 cell_1rw
* cell instance $25529 r0 *1 96.585,163.8
X$25529 340 635 341 644 645 cell_1rw
* cell instance $25530 m0 *1 96.585,166.53
X$25530 340 637 341 644 645 cell_1rw
* cell instance $25531 m0 *1 96.585,169.26
X$25531 340 639 341 644 645 cell_1rw
* cell instance $25532 r0 *1 96.585,166.53
X$25532 340 636 341 644 645 cell_1rw
* cell instance $25533 m0 *1 96.585,171.99
X$25533 340 640 341 644 645 cell_1rw
* cell instance $25534 r0 *1 96.585,169.26
X$25534 340 638 341 644 645 cell_1rw
* cell instance $25535 r0 *1 96.585,171.99
X$25535 340 641 341 644 645 cell_1rw
* cell instance $25536 m0 *1 96.585,174.72
X$25536 340 642 341 644 645 cell_1rw
* cell instance $25537 r0 *1 96.585,174.72
X$25537 340 643 341 644 645 cell_1rw
* cell instance $25538 m0 *1 97.29,90.09
X$25538 342 581 343 644 645 cell_1rw
* cell instance $25539 r0 *1 97.29,90.09
X$25539 342 580 343 644 645 cell_1rw
* cell instance $25540 m0 *1 97.29,92.82
X$25540 342 583 343 644 645 cell_1rw
* cell instance $25541 r0 *1 97.29,92.82
X$25541 342 582 343 644 645 cell_1rw
* cell instance $25542 m0 *1 97.29,95.55
X$25542 342 584 343 644 645 cell_1rw
* cell instance $25543 r0 *1 97.29,95.55
X$25543 342 585 343 644 645 cell_1rw
* cell instance $25544 m0 *1 97.29,98.28
X$25544 342 586 343 644 645 cell_1rw
* cell instance $25545 r0 *1 97.29,98.28
X$25545 342 587 343 644 645 cell_1rw
* cell instance $25546 m0 *1 97.29,101.01
X$25546 342 588 343 644 645 cell_1rw
* cell instance $25547 m0 *1 97.29,103.74
X$25547 342 590 343 644 645 cell_1rw
* cell instance $25548 r0 *1 97.29,101.01
X$25548 342 589 343 644 645 cell_1rw
* cell instance $25549 r0 *1 97.29,103.74
X$25549 342 591 343 644 645 cell_1rw
* cell instance $25550 m0 *1 97.29,106.47
X$25550 342 593 343 644 645 cell_1rw
* cell instance $25551 r0 *1 97.29,106.47
X$25551 342 592 343 644 645 cell_1rw
* cell instance $25552 m0 *1 97.29,109.2
X$25552 342 594 343 644 645 cell_1rw
* cell instance $25553 r0 *1 97.29,109.2
X$25553 342 595 343 644 645 cell_1rw
* cell instance $25554 m0 *1 97.29,111.93
X$25554 342 597 343 644 645 cell_1rw
* cell instance $25555 r0 *1 97.29,111.93
X$25555 342 596 343 644 645 cell_1rw
* cell instance $25556 m0 *1 97.29,114.66
X$25556 342 598 343 644 645 cell_1rw
* cell instance $25557 r0 *1 97.29,114.66
X$25557 342 599 343 644 645 cell_1rw
* cell instance $25558 m0 *1 97.29,117.39
X$25558 342 600 343 644 645 cell_1rw
* cell instance $25559 r0 *1 97.29,117.39
X$25559 342 601 343 644 645 cell_1rw
* cell instance $25560 m0 *1 97.29,120.12
X$25560 342 602 343 644 645 cell_1rw
* cell instance $25561 r0 *1 97.29,120.12
X$25561 342 603 343 644 645 cell_1rw
* cell instance $25562 m0 *1 97.29,122.85
X$25562 342 604 343 644 645 cell_1rw
* cell instance $25563 r0 *1 97.29,122.85
X$25563 342 605 343 644 645 cell_1rw
* cell instance $25564 m0 *1 97.29,125.58
X$25564 342 606 343 644 645 cell_1rw
* cell instance $25565 r0 *1 97.29,125.58
X$25565 342 607 343 644 645 cell_1rw
* cell instance $25566 m0 *1 97.29,128.31
X$25566 342 609 343 644 645 cell_1rw
* cell instance $25567 r0 *1 97.29,128.31
X$25567 342 608 343 644 645 cell_1rw
* cell instance $25568 m0 *1 97.29,131.04
X$25568 342 610 343 644 645 cell_1rw
* cell instance $25569 r0 *1 97.29,131.04
X$25569 342 611 343 644 645 cell_1rw
* cell instance $25570 m0 *1 97.29,133.77
X$25570 342 612 343 644 645 cell_1rw
* cell instance $25571 r0 *1 97.29,133.77
X$25571 342 613 343 644 645 cell_1rw
* cell instance $25572 m0 *1 97.29,136.5
X$25572 342 615 343 644 645 cell_1rw
* cell instance $25573 r0 *1 97.29,136.5
X$25573 342 614 343 644 645 cell_1rw
* cell instance $25574 m0 *1 97.29,139.23
X$25574 342 617 343 644 645 cell_1rw
* cell instance $25575 r0 *1 97.29,139.23
X$25575 342 616 343 644 645 cell_1rw
* cell instance $25576 m0 *1 97.29,141.96
X$25576 342 618 343 644 645 cell_1rw
* cell instance $25577 r0 *1 97.29,141.96
X$25577 342 619 343 644 645 cell_1rw
* cell instance $25578 m0 *1 97.29,144.69
X$25578 342 620 343 644 645 cell_1rw
* cell instance $25579 r0 *1 97.29,144.69
X$25579 342 621 343 644 645 cell_1rw
* cell instance $25580 m0 *1 97.29,147.42
X$25580 342 622 343 644 645 cell_1rw
* cell instance $25581 r0 *1 97.29,147.42
X$25581 342 623 343 644 645 cell_1rw
* cell instance $25582 m0 *1 97.29,150.15
X$25582 342 624 343 644 645 cell_1rw
* cell instance $25583 r0 *1 97.29,150.15
X$25583 342 625 343 644 645 cell_1rw
* cell instance $25584 m0 *1 97.29,152.88
X$25584 342 626 343 644 645 cell_1rw
* cell instance $25585 r0 *1 97.29,152.88
X$25585 342 627 343 644 645 cell_1rw
* cell instance $25586 m0 *1 97.29,155.61
X$25586 342 628 343 644 645 cell_1rw
* cell instance $25587 m0 *1 97.29,158.34
X$25587 342 630 343 644 645 cell_1rw
* cell instance $25588 r0 *1 97.29,155.61
X$25588 342 629 343 644 645 cell_1rw
* cell instance $25589 r0 *1 97.29,158.34
X$25589 342 631 343 644 645 cell_1rw
* cell instance $25590 m0 *1 97.29,161.07
X$25590 342 632 343 644 645 cell_1rw
* cell instance $25591 r0 *1 97.29,161.07
X$25591 342 633 343 644 645 cell_1rw
* cell instance $25592 m0 *1 97.29,163.8
X$25592 342 634 343 644 645 cell_1rw
* cell instance $25593 r0 *1 97.29,163.8
X$25593 342 635 343 644 645 cell_1rw
* cell instance $25594 m0 *1 97.29,166.53
X$25594 342 637 343 644 645 cell_1rw
* cell instance $25595 r0 *1 97.29,166.53
X$25595 342 636 343 644 645 cell_1rw
* cell instance $25596 m0 *1 97.29,169.26
X$25596 342 639 343 644 645 cell_1rw
* cell instance $25597 m0 *1 97.29,171.99
X$25597 342 640 343 644 645 cell_1rw
* cell instance $25598 r0 *1 97.29,169.26
X$25598 342 638 343 644 645 cell_1rw
* cell instance $25599 r0 *1 97.29,171.99
X$25599 342 641 343 644 645 cell_1rw
* cell instance $25600 m0 *1 97.29,174.72
X$25600 342 642 343 644 645 cell_1rw
* cell instance $25601 r0 *1 97.29,174.72
X$25601 342 643 343 644 645 cell_1rw
* cell instance $25602 m0 *1 97.995,90.09
X$25602 344 581 345 644 645 cell_1rw
* cell instance $25603 r0 *1 97.995,90.09
X$25603 344 580 345 644 645 cell_1rw
* cell instance $25604 m0 *1 97.995,92.82
X$25604 344 583 345 644 645 cell_1rw
* cell instance $25605 r0 *1 97.995,92.82
X$25605 344 582 345 644 645 cell_1rw
* cell instance $25606 m0 *1 97.995,95.55
X$25606 344 584 345 644 645 cell_1rw
* cell instance $25607 r0 *1 97.995,95.55
X$25607 344 585 345 644 645 cell_1rw
* cell instance $25608 m0 *1 97.995,98.28
X$25608 344 586 345 644 645 cell_1rw
* cell instance $25609 r0 *1 97.995,98.28
X$25609 344 587 345 644 645 cell_1rw
* cell instance $25610 m0 *1 97.995,101.01
X$25610 344 588 345 644 645 cell_1rw
* cell instance $25611 r0 *1 97.995,101.01
X$25611 344 589 345 644 645 cell_1rw
* cell instance $25612 m0 *1 97.995,103.74
X$25612 344 590 345 644 645 cell_1rw
* cell instance $25613 r0 *1 97.995,103.74
X$25613 344 591 345 644 645 cell_1rw
* cell instance $25614 m0 *1 97.995,106.47
X$25614 344 593 345 644 645 cell_1rw
* cell instance $25615 r0 *1 97.995,106.47
X$25615 344 592 345 644 645 cell_1rw
* cell instance $25616 m0 *1 97.995,109.2
X$25616 344 594 345 644 645 cell_1rw
* cell instance $25617 r0 *1 97.995,109.2
X$25617 344 595 345 644 645 cell_1rw
* cell instance $25618 m0 *1 97.995,111.93
X$25618 344 597 345 644 645 cell_1rw
* cell instance $25619 r0 *1 97.995,111.93
X$25619 344 596 345 644 645 cell_1rw
* cell instance $25620 m0 *1 97.995,114.66
X$25620 344 598 345 644 645 cell_1rw
* cell instance $25621 r0 *1 97.995,114.66
X$25621 344 599 345 644 645 cell_1rw
* cell instance $25622 m0 *1 97.995,117.39
X$25622 344 600 345 644 645 cell_1rw
* cell instance $25623 m0 *1 97.995,120.12
X$25623 344 602 345 644 645 cell_1rw
* cell instance $25624 r0 *1 97.995,117.39
X$25624 344 601 345 644 645 cell_1rw
* cell instance $25625 r0 *1 97.995,120.12
X$25625 344 603 345 644 645 cell_1rw
* cell instance $25626 m0 *1 97.995,122.85
X$25626 344 604 345 644 645 cell_1rw
* cell instance $25627 r0 *1 97.995,122.85
X$25627 344 605 345 644 645 cell_1rw
* cell instance $25628 m0 *1 97.995,125.58
X$25628 344 606 345 644 645 cell_1rw
* cell instance $25629 r0 *1 97.995,125.58
X$25629 344 607 345 644 645 cell_1rw
* cell instance $25630 m0 *1 97.995,128.31
X$25630 344 609 345 644 645 cell_1rw
* cell instance $25631 r0 *1 97.995,128.31
X$25631 344 608 345 644 645 cell_1rw
* cell instance $25632 m0 *1 97.995,131.04
X$25632 344 610 345 644 645 cell_1rw
* cell instance $25633 r0 *1 97.995,131.04
X$25633 344 611 345 644 645 cell_1rw
* cell instance $25634 m0 *1 97.995,133.77
X$25634 344 612 345 644 645 cell_1rw
* cell instance $25635 r0 *1 97.995,133.77
X$25635 344 613 345 644 645 cell_1rw
* cell instance $25636 m0 *1 97.995,136.5
X$25636 344 615 345 644 645 cell_1rw
* cell instance $25637 m0 *1 97.995,139.23
X$25637 344 617 345 644 645 cell_1rw
* cell instance $25638 r0 *1 97.995,136.5
X$25638 344 614 345 644 645 cell_1rw
* cell instance $25639 m0 *1 97.995,141.96
X$25639 344 618 345 644 645 cell_1rw
* cell instance $25640 r0 *1 97.995,139.23
X$25640 344 616 345 644 645 cell_1rw
* cell instance $25641 r0 *1 97.995,141.96
X$25641 344 619 345 644 645 cell_1rw
* cell instance $25642 m0 *1 97.995,144.69
X$25642 344 620 345 644 645 cell_1rw
* cell instance $25643 r0 *1 97.995,144.69
X$25643 344 621 345 644 645 cell_1rw
* cell instance $25644 m0 *1 97.995,147.42
X$25644 344 622 345 644 645 cell_1rw
* cell instance $25645 r0 *1 97.995,147.42
X$25645 344 623 345 644 645 cell_1rw
* cell instance $25646 m0 *1 97.995,150.15
X$25646 344 624 345 644 645 cell_1rw
* cell instance $25647 r0 *1 97.995,150.15
X$25647 344 625 345 644 645 cell_1rw
* cell instance $25648 m0 *1 97.995,152.88
X$25648 344 626 345 644 645 cell_1rw
* cell instance $25649 r0 *1 97.995,152.88
X$25649 344 627 345 644 645 cell_1rw
* cell instance $25650 m0 *1 97.995,155.61
X$25650 344 628 345 644 645 cell_1rw
* cell instance $25651 m0 *1 97.995,158.34
X$25651 344 630 345 644 645 cell_1rw
* cell instance $25652 r0 *1 97.995,155.61
X$25652 344 629 345 644 645 cell_1rw
* cell instance $25653 r0 *1 97.995,158.34
X$25653 344 631 345 644 645 cell_1rw
* cell instance $25654 m0 *1 97.995,161.07
X$25654 344 632 345 644 645 cell_1rw
* cell instance $25655 r0 *1 97.995,161.07
X$25655 344 633 345 644 645 cell_1rw
* cell instance $25656 m0 *1 97.995,163.8
X$25656 344 634 345 644 645 cell_1rw
* cell instance $25657 r0 *1 97.995,163.8
X$25657 344 635 345 644 645 cell_1rw
* cell instance $25658 m0 *1 97.995,166.53
X$25658 344 637 345 644 645 cell_1rw
* cell instance $25659 r0 *1 97.995,166.53
X$25659 344 636 345 644 645 cell_1rw
* cell instance $25660 m0 *1 97.995,169.26
X$25660 344 639 345 644 645 cell_1rw
* cell instance $25661 r0 *1 97.995,169.26
X$25661 344 638 345 644 645 cell_1rw
* cell instance $25662 m0 *1 97.995,171.99
X$25662 344 640 345 644 645 cell_1rw
* cell instance $25663 r0 *1 97.995,171.99
X$25663 344 641 345 644 645 cell_1rw
* cell instance $25664 m0 *1 97.995,174.72
X$25664 344 642 345 644 645 cell_1rw
* cell instance $25665 r0 *1 97.995,174.72
X$25665 344 643 345 644 645 cell_1rw
* cell instance $25666 m0 *1 98.7,90.09
X$25666 346 581 347 644 645 cell_1rw
* cell instance $25667 r0 *1 98.7,90.09
X$25667 346 580 347 644 645 cell_1rw
* cell instance $25668 m0 *1 98.7,92.82
X$25668 346 583 347 644 645 cell_1rw
* cell instance $25669 r0 *1 98.7,92.82
X$25669 346 582 347 644 645 cell_1rw
* cell instance $25670 m0 *1 98.7,95.55
X$25670 346 584 347 644 645 cell_1rw
* cell instance $25671 r0 *1 98.7,95.55
X$25671 346 585 347 644 645 cell_1rw
* cell instance $25672 m0 *1 98.7,98.28
X$25672 346 586 347 644 645 cell_1rw
* cell instance $25673 m0 *1 98.7,101.01
X$25673 346 588 347 644 645 cell_1rw
* cell instance $25674 r0 *1 98.7,98.28
X$25674 346 587 347 644 645 cell_1rw
* cell instance $25675 r0 *1 98.7,101.01
X$25675 346 589 347 644 645 cell_1rw
* cell instance $25676 m0 *1 98.7,103.74
X$25676 346 590 347 644 645 cell_1rw
* cell instance $25677 m0 *1 98.7,106.47
X$25677 346 593 347 644 645 cell_1rw
* cell instance $25678 r0 *1 98.7,103.74
X$25678 346 591 347 644 645 cell_1rw
* cell instance $25679 r0 *1 98.7,106.47
X$25679 346 592 347 644 645 cell_1rw
* cell instance $25680 m0 *1 98.7,109.2
X$25680 346 594 347 644 645 cell_1rw
* cell instance $25681 r0 *1 98.7,109.2
X$25681 346 595 347 644 645 cell_1rw
* cell instance $25682 m0 *1 98.7,111.93
X$25682 346 597 347 644 645 cell_1rw
* cell instance $25683 m0 *1 98.7,114.66
X$25683 346 598 347 644 645 cell_1rw
* cell instance $25684 r0 *1 98.7,111.93
X$25684 346 596 347 644 645 cell_1rw
* cell instance $25685 r0 *1 98.7,114.66
X$25685 346 599 347 644 645 cell_1rw
* cell instance $25686 m0 *1 98.7,117.39
X$25686 346 600 347 644 645 cell_1rw
* cell instance $25687 r0 *1 98.7,117.39
X$25687 346 601 347 644 645 cell_1rw
* cell instance $25688 m0 *1 98.7,120.12
X$25688 346 602 347 644 645 cell_1rw
* cell instance $25689 r0 *1 98.7,120.12
X$25689 346 603 347 644 645 cell_1rw
* cell instance $25690 m0 *1 98.7,122.85
X$25690 346 604 347 644 645 cell_1rw
* cell instance $25691 r0 *1 98.7,122.85
X$25691 346 605 347 644 645 cell_1rw
* cell instance $25692 m0 *1 98.7,125.58
X$25692 346 606 347 644 645 cell_1rw
* cell instance $25693 r0 *1 98.7,125.58
X$25693 346 607 347 644 645 cell_1rw
* cell instance $25694 m0 *1 98.7,128.31
X$25694 346 609 347 644 645 cell_1rw
* cell instance $25695 r0 *1 98.7,128.31
X$25695 346 608 347 644 645 cell_1rw
* cell instance $25696 m0 *1 98.7,131.04
X$25696 346 610 347 644 645 cell_1rw
* cell instance $25697 m0 *1 98.7,133.77
X$25697 346 612 347 644 645 cell_1rw
* cell instance $25698 r0 *1 98.7,131.04
X$25698 346 611 347 644 645 cell_1rw
* cell instance $25699 r0 *1 98.7,133.77
X$25699 346 613 347 644 645 cell_1rw
* cell instance $25700 m0 *1 98.7,136.5
X$25700 346 615 347 644 645 cell_1rw
* cell instance $25701 r0 *1 98.7,136.5
X$25701 346 614 347 644 645 cell_1rw
* cell instance $25702 m0 *1 98.7,139.23
X$25702 346 617 347 644 645 cell_1rw
* cell instance $25703 r0 *1 98.7,139.23
X$25703 346 616 347 644 645 cell_1rw
* cell instance $25704 m0 *1 98.7,141.96
X$25704 346 618 347 644 645 cell_1rw
* cell instance $25705 m0 *1 98.7,144.69
X$25705 346 620 347 644 645 cell_1rw
* cell instance $25706 r0 *1 98.7,141.96
X$25706 346 619 347 644 645 cell_1rw
* cell instance $25707 r0 *1 98.7,144.69
X$25707 346 621 347 644 645 cell_1rw
* cell instance $25708 m0 *1 98.7,147.42
X$25708 346 622 347 644 645 cell_1rw
* cell instance $25709 r0 *1 98.7,147.42
X$25709 346 623 347 644 645 cell_1rw
* cell instance $25710 m0 *1 98.7,150.15
X$25710 346 624 347 644 645 cell_1rw
* cell instance $25711 m0 *1 98.7,152.88
X$25711 346 626 347 644 645 cell_1rw
* cell instance $25712 r0 *1 98.7,150.15
X$25712 346 625 347 644 645 cell_1rw
* cell instance $25713 r0 *1 98.7,152.88
X$25713 346 627 347 644 645 cell_1rw
* cell instance $25714 m0 *1 98.7,155.61
X$25714 346 628 347 644 645 cell_1rw
* cell instance $25715 r0 *1 98.7,155.61
X$25715 346 629 347 644 645 cell_1rw
* cell instance $25716 m0 *1 98.7,158.34
X$25716 346 630 347 644 645 cell_1rw
* cell instance $25717 r0 *1 98.7,158.34
X$25717 346 631 347 644 645 cell_1rw
* cell instance $25718 m0 *1 98.7,161.07
X$25718 346 632 347 644 645 cell_1rw
* cell instance $25719 r0 *1 98.7,161.07
X$25719 346 633 347 644 645 cell_1rw
* cell instance $25720 m0 *1 98.7,163.8
X$25720 346 634 347 644 645 cell_1rw
* cell instance $25721 r0 *1 98.7,163.8
X$25721 346 635 347 644 645 cell_1rw
* cell instance $25722 m0 *1 98.7,166.53
X$25722 346 637 347 644 645 cell_1rw
* cell instance $25723 r0 *1 98.7,166.53
X$25723 346 636 347 644 645 cell_1rw
* cell instance $25724 m0 *1 98.7,169.26
X$25724 346 639 347 644 645 cell_1rw
* cell instance $25725 r0 *1 98.7,169.26
X$25725 346 638 347 644 645 cell_1rw
* cell instance $25726 m0 *1 98.7,171.99
X$25726 346 640 347 644 645 cell_1rw
* cell instance $25727 r0 *1 98.7,171.99
X$25727 346 641 347 644 645 cell_1rw
* cell instance $25728 m0 *1 98.7,174.72
X$25728 346 642 347 644 645 cell_1rw
* cell instance $25729 r0 *1 98.7,174.72
X$25729 346 643 347 644 645 cell_1rw
* cell instance $25730 m0 *1 99.405,90.09
X$25730 348 581 349 644 645 cell_1rw
* cell instance $25731 m0 *1 99.405,92.82
X$25731 348 583 349 644 645 cell_1rw
* cell instance $25732 r0 *1 99.405,90.09
X$25732 348 580 349 644 645 cell_1rw
* cell instance $25733 m0 *1 99.405,95.55
X$25733 348 584 349 644 645 cell_1rw
* cell instance $25734 r0 *1 99.405,92.82
X$25734 348 582 349 644 645 cell_1rw
* cell instance $25735 m0 *1 99.405,98.28
X$25735 348 586 349 644 645 cell_1rw
* cell instance $25736 r0 *1 99.405,95.55
X$25736 348 585 349 644 645 cell_1rw
* cell instance $25737 r0 *1 99.405,98.28
X$25737 348 587 349 644 645 cell_1rw
* cell instance $25738 m0 *1 99.405,101.01
X$25738 348 588 349 644 645 cell_1rw
* cell instance $25739 m0 *1 99.405,103.74
X$25739 348 590 349 644 645 cell_1rw
* cell instance $25740 r0 *1 99.405,101.01
X$25740 348 589 349 644 645 cell_1rw
* cell instance $25741 m0 *1 99.405,106.47
X$25741 348 593 349 644 645 cell_1rw
* cell instance $25742 r0 *1 99.405,103.74
X$25742 348 591 349 644 645 cell_1rw
* cell instance $25743 r0 *1 99.405,106.47
X$25743 348 592 349 644 645 cell_1rw
* cell instance $25744 m0 *1 99.405,109.2
X$25744 348 594 349 644 645 cell_1rw
* cell instance $25745 r0 *1 99.405,109.2
X$25745 348 595 349 644 645 cell_1rw
* cell instance $25746 m0 *1 99.405,111.93
X$25746 348 597 349 644 645 cell_1rw
* cell instance $25747 m0 *1 99.405,114.66
X$25747 348 598 349 644 645 cell_1rw
* cell instance $25748 r0 *1 99.405,111.93
X$25748 348 596 349 644 645 cell_1rw
* cell instance $25749 r0 *1 99.405,114.66
X$25749 348 599 349 644 645 cell_1rw
* cell instance $25750 m0 *1 99.405,117.39
X$25750 348 600 349 644 645 cell_1rw
* cell instance $25751 r0 *1 99.405,117.39
X$25751 348 601 349 644 645 cell_1rw
* cell instance $25752 m0 *1 99.405,120.12
X$25752 348 602 349 644 645 cell_1rw
* cell instance $25753 r0 *1 99.405,120.12
X$25753 348 603 349 644 645 cell_1rw
* cell instance $25754 m0 *1 99.405,122.85
X$25754 348 604 349 644 645 cell_1rw
* cell instance $25755 r0 *1 99.405,122.85
X$25755 348 605 349 644 645 cell_1rw
* cell instance $25756 m0 *1 99.405,125.58
X$25756 348 606 349 644 645 cell_1rw
* cell instance $25757 r0 *1 99.405,125.58
X$25757 348 607 349 644 645 cell_1rw
* cell instance $25758 m0 *1 99.405,128.31
X$25758 348 609 349 644 645 cell_1rw
* cell instance $25759 r0 *1 99.405,128.31
X$25759 348 608 349 644 645 cell_1rw
* cell instance $25760 m0 *1 99.405,131.04
X$25760 348 610 349 644 645 cell_1rw
* cell instance $25761 r0 *1 99.405,131.04
X$25761 348 611 349 644 645 cell_1rw
* cell instance $25762 m0 *1 99.405,133.77
X$25762 348 612 349 644 645 cell_1rw
* cell instance $25763 r0 *1 99.405,133.77
X$25763 348 613 349 644 645 cell_1rw
* cell instance $25764 m0 *1 99.405,136.5
X$25764 348 615 349 644 645 cell_1rw
* cell instance $25765 r0 *1 99.405,136.5
X$25765 348 614 349 644 645 cell_1rw
* cell instance $25766 m0 *1 99.405,139.23
X$25766 348 617 349 644 645 cell_1rw
* cell instance $25767 r0 *1 99.405,139.23
X$25767 348 616 349 644 645 cell_1rw
* cell instance $25768 m0 *1 99.405,141.96
X$25768 348 618 349 644 645 cell_1rw
* cell instance $25769 r0 *1 99.405,141.96
X$25769 348 619 349 644 645 cell_1rw
* cell instance $25770 m0 *1 99.405,144.69
X$25770 348 620 349 644 645 cell_1rw
* cell instance $25771 r0 *1 99.405,144.69
X$25771 348 621 349 644 645 cell_1rw
* cell instance $25772 m0 *1 99.405,147.42
X$25772 348 622 349 644 645 cell_1rw
* cell instance $25773 m0 *1 99.405,150.15
X$25773 348 624 349 644 645 cell_1rw
* cell instance $25774 r0 *1 99.405,147.42
X$25774 348 623 349 644 645 cell_1rw
* cell instance $25775 m0 *1 99.405,152.88
X$25775 348 626 349 644 645 cell_1rw
* cell instance $25776 r0 *1 99.405,150.15
X$25776 348 625 349 644 645 cell_1rw
* cell instance $25777 r0 *1 99.405,152.88
X$25777 348 627 349 644 645 cell_1rw
* cell instance $25778 m0 *1 99.405,155.61
X$25778 348 628 349 644 645 cell_1rw
* cell instance $25779 m0 *1 99.405,158.34
X$25779 348 630 349 644 645 cell_1rw
* cell instance $25780 r0 *1 99.405,155.61
X$25780 348 629 349 644 645 cell_1rw
* cell instance $25781 r0 *1 99.405,158.34
X$25781 348 631 349 644 645 cell_1rw
* cell instance $25782 m0 *1 99.405,161.07
X$25782 348 632 349 644 645 cell_1rw
* cell instance $25783 r0 *1 99.405,161.07
X$25783 348 633 349 644 645 cell_1rw
* cell instance $25784 m0 *1 99.405,163.8
X$25784 348 634 349 644 645 cell_1rw
* cell instance $25785 r0 *1 99.405,163.8
X$25785 348 635 349 644 645 cell_1rw
* cell instance $25786 m0 *1 99.405,166.53
X$25786 348 637 349 644 645 cell_1rw
* cell instance $25787 r0 *1 99.405,166.53
X$25787 348 636 349 644 645 cell_1rw
* cell instance $25788 m0 *1 99.405,169.26
X$25788 348 639 349 644 645 cell_1rw
* cell instance $25789 m0 *1 99.405,171.99
X$25789 348 640 349 644 645 cell_1rw
* cell instance $25790 r0 *1 99.405,169.26
X$25790 348 638 349 644 645 cell_1rw
* cell instance $25791 r0 *1 99.405,171.99
X$25791 348 641 349 644 645 cell_1rw
* cell instance $25792 m0 *1 99.405,174.72
X$25792 348 642 349 644 645 cell_1rw
* cell instance $25793 r0 *1 99.405,174.72
X$25793 348 643 349 644 645 cell_1rw
* cell instance $25794 m0 *1 100.11,90.09
X$25794 350 581 351 644 645 cell_1rw
* cell instance $25795 r0 *1 100.11,90.09
X$25795 350 580 351 644 645 cell_1rw
* cell instance $25796 m0 *1 100.11,92.82
X$25796 350 583 351 644 645 cell_1rw
* cell instance $25797 r0 *1 100.11,92.82
X$25797 350 582 351 644 645 cell_1rw
* cell instance $25798 m0 *1 100.11,95.55
X$25798 350 584 351 644 645 cell_1rw
* cell instance $25799 m0 *1 100.11,98.28
X$25799 350 586 351 644 645 cell_1rw
* cell instance $25800 r0 *1 100.11,95.55
X$25800 350 585 351 644 645 cell_1rw
* cell instance $25801 r0 *1 100.11,98.28
X$25801 350 587 351 644 645 cell_1rw
* cell instance $25802 m0 *1 100.11,101.01
X$25802 350 588 351 644 645 cell_1rw
* cell instance $25803 r0 *1 100.11,101.01
X$25803 350 589 351 644 645 cell_1rw
* cell instance $25804 m0 *1 100.11,103.74
X$25804 350 590 351 644 645 cell_1rw
* cell instance $25805 r0 *1 100.11,103.74
X$25805 350 591 351 644 645 cell_1rw
* cell instance $25806 m0 *1 100.11,106.47
X$25806 350 593 351 644 645 cell_1rw
* cell instance $25807 r0 *1 100.11,106.47
X$25807 350 592 351 644 645 cell_1rw
* cell instance $25808 m0 *1 100.11,109.2
X$25808 350 594 351 644 645 cell_1rw
* cell instance $25809 r0 *1 100.11,109.2
X$25809 350 595 351 644 645 cell_1rw
* cell instance $25810 m0 *1 100.11,111.93
X$25810 350 597 351 644 645 cell_1rw
* cell instance $25811 r0 *1 100.11,111.93
X$25811 350 596 351 644 645 cell_1rw
* cell instance $25812 m0 *1 100.11,114.66
X$25812 350 598 351 644 645 cell_1rw
* cell instance $25813 r0 *1 100.11,114.66
X$25813 350 599 351 644 645 cell_1rw
* cell instance $25814 m0 *1 100.11,117.39
X$25814 350 600 351 644 645 cell_1rw
* cell instance $25815 r0 *1 100.11,117.39
X$25815 350 601 351 644 645 cell_1rw
* cell instance $25816 m0 *1 100.11,120.12
X$25816 350 602 351 644 645 cell_1rw
* cell instance $25817 r0 *1 100.11,120.12
X$25817 350 603 351 644 645 cell_1rw
* cell instance $25818 m0 *1 100.11,122.85
X$25818 350 604 351 644 645 cell_1rw
* cell instance $25819 r0 *1 100.11,122.85
X$25819 350 605 351 644 645 cell_1rw
* cell instance $25820 m0 *1 100.11,125.58
X$25820 350 606 351 644 645 cell_1rw
* cell instance $25821 r0 *1 100.11,125.58
X$25821 350 607 351 644 645 cell_1rw
* cell instance $25822 m0 *1 100.11,128.31
X$25822 350 609 351 644 645 cell_1rw
* cell instance $25823 r0 *1 100.11,128.31
X$25823 350 608 351 644 645 cell_1rw
* cell instance $25824 m0 *1 100.11,131.04
X$25824 350 610 351 644 645 cell_1rw
* cell instance $25825 r0 *1 100.11,131.04
X$25825 350 611 351 644 645 cell_1rw
* cell instance $25826 m0 *1 100.11,133.77
X$25826 350 612 351 644 645 cell_1rw
* cell instance $25827 r0 *1 100.11,133.77
X$25827 350 613 351 644 645 cell_1rw
* cell instance $25828 m0 *1 100.11,136.5
X$25828 350 615 351 644 645 cell_1rw
* cell instance $25829 m0 *1 100.11,139.23
X$25829 350 617 351 644 645 cell_1rw
* cell instance $25830 r0 *1 100.11,136.5
X$25830 350 614 351 644 645 cell_1rw
* cell instance $25831 r0 *1 100.11,139.23
X$25831 350 616 351 644 645 cell_1rw
* cell instance $25832 m0 *1 100.11,141.96
X$25832 350 618 351 644 645 cell_1rw
* cell instance $25833 m0 *1 100.11,144.69
X$25833 350 620 351 644 645 cell_1rw
* cell instance $25834 r0 *1 100.11,141.96
X$25834 350 619 351 644 645 cell_1rw
* cell instance $25835 r0 *1 100.11,144.69
X$25835 350 621 351 644 645 cell_1rw
* cell instance $25836 m0 *1 100.11,147.42
X$25836 350 622 351 644 645 cell_1rw
* cell instance $25837 r0 *1 100.11,147.42
X$25837 350 623 351 644 645 cell_1rw
* cell instance $25838 m0 *1 100.11,150.15
X$25838 350 624 351 644 645 cell_1rw
* cell instance $25839 r0 *1 100.11,150.15
X$25839 350 625 351 644 645 cell_1rw
* cell instance $25840 m0 *1 100.11,152.88
X$25840 350 626 351 644 645 cell_1rw
* cell instance $25841 r0 *1 100.11,152.88
X$25841 350 627 351 644 645 cell_1rw
* cell instance $25842 m0 *1 100.11,155.61
X$25842 350 628 351 644 645 cell_1rw
* cell instance $25843 m0 *1 100.11,158.34
X$25843 350 630 351 644 645 cell_1rw
* cell instance $25844 r0 *1 100.11,155.61
X$25844 350 629 351 644 645 cell_1rw
* cell instance $25845 r0 *1 100.11,158.34
X$25845 350 631 351 644 645 cell_1rw
* cell instance $25846 m0 *1 100.11,161.07
X$25846 350 632 351 644 645 cell_1rw
* cell instance $25847 r0 *1 100.11,161.07
X$25847 350 633 351 644 645 cell_1rw
* cell instance $25848 m0 *1 100.11,163.8
X$25848 350 634 351 644 645 cell_1rw
* cell instance $25849 m0 *1 100.11,166.53
X$25849 350 637 351 644 645 cell_1rw
* cell instance $25850 r0 *1 100.11,163.8
X$25850 350 635 351 644 645 cell_1rw
* cell instance $25851 r0 *1 100.11,166.53
X$25851 350 636 351 644 645 cell_1rw
* cell instance $25852 m0 *1 100.11,169.26
X$25852 350 639 351 644 645 cell_1rw
* cell instance $25853 r0 *1 100.11,169.26
X$25853 350 638 351 644 645 cell_1rw
* cell instance $25854 m0 *1 100.11,171.99
X$25854 350 640 351 644 645 cell_1rw
* cell instance $25855 m0 *1 100.11,174.72
X$25855 350 642 351 644 645 cell_1rw
* cell instance $25856 r0 *1 100.11,171.99
X$25856 350 641 351 644 645 cell_1rw
* cell instance $25857 r0 *1 100.11,174.72
X$25857 350 643 351 644 645 cell_1rw
* cell instance $25858 m0 *1 100.815,90.09
X$25858 352 581 353 644 645 cell_1rw
* cell instance $25859 r0 *1 100.815,90.09
X$25859 352 580 353 644 645 cell_1rw
* cell instance $25860 m0 *1 100.815,92.82
X$25860 352 583 353 644 645 cell_1rw
* cell instance $25861 r0 *1 100.815,92.82
X$25861 352 582 353 644 645 cell_1rw
* cell instance $25862 m0 *1 100.815,95.55
X$25862 352 584 353 644 645 cell_1rw
* cell instance $25863 r0 *1 100.815,95.55
X$25863 352 585 353 644 645 cell_1rw
* cell instance $25864 m0 *1 100.815,98.28
X$25864 352 586 353 644 645 cell_1rw
* cell instance $25865 r0 *1 100.815,98.28
X$25865 352 587 353 644 645 cell_1rw
* cell instance $25866 m0 *1 100.815,101.01
X$25866 352 588 353 644 645 cell_1rw
* cell instance $25867 r0 *1 100.815,101.01
X$25867 352 589 353 644 645 cell_1rw
* cell instance $25868 m0 *1 100.815,103.74
X$25868 352 590 353 644 645 cell_1rw
* cell instance $25869 r0 *1 100.815,103.74
X$25869 352 591 353 644 645 cell_1rw
* cell instance $25870 m0 *1 100.815,106.47
X$25870 352 593 353 644 645 cell_1rw
* cell instance $25871 r0 *1 100.815,106.47
X$25871 352 592 353 644 645 cell_1rw
* cell instance $25872 m0 *1 100.815,109.2
X$25872 352 594 353 644 645 cell_1rw
* cell instance $25873 r0 *1 100.815,109.2
X$25873 352 595 353 644 645 cell_1rw
* cell instance $25874 m0 *1 100.815,111.93
X$25874 352 597 353 644 645 cell_1rw
* cell instance $25875 r0 *1 100.815,111.93
X$25875 352 596 353 644 645 cell_1rw
* cell instance $25876 m0 *1 100.815,114.66
X$25876 352 598 353 644 645 cell_1rw
* cell instance $25877 r0 *1 100.815,114.66
X$25877 352 599 353 644 645 cell_1rw
* cell instance $25878 m0 *1 100.815,117.39
X$25878 352 600 353 644 645 cell_1rw
* cell instance $25879 m0 *1 100.815,120.12
X$25879 352 602 353 644 645 cell_1rw
* cell instance $25880 r0 *1 100.815,117.39
X$25880 352 601 353 644 645 cell_1rw
* cell instance $25881 r0 *1 100.815,120.12
X$25881 352 603 353 644 645 cell_1rw
* cell instance $25882 m0 *1 100.815,122.85
X$25882 352 604 353 644 645 cell_1rw
* cell instance $25883 r0 *1 100.815,122.85
X$25883 352 605 353 644 645 cell_1rw
* cell instance $25884 m0 *1 100.815,125.58
X$25884 352 606 353 644 645 cell_1rw
* cell instance $25885 m0 *1 100.815,128.31
X$25885 352 609 353 644 645 cell_1rw
* cell instance $25886 r0 *1 100.815,125.58
X$25886 352 607 353 644 645 cell_1rw
* cell instance $25887 m0 *1 100.815,131.04
X$25887 352 610 353 644 645 cell_1rw
* cell instance $25888 r0 *1 100.815,128.31
X$25888 352 608 353 644 645 cell_1rw
* cell instance $25889 r0 *1 100.815,131.04
X$25889 352 611 353 644 645 cell_1rw
* cell instance $25890 m0 *1 100.815,133.77
X$25890 352 612 353 644 645 cell_1rw
* cell instance $25891 m0 *1 100.815,136.5
X$25891 352 615 353 644 645 cell_1rw
* cell instance $25892 r0 *1 100.815,133.77
X$25892 352 613 353 644 645 cell_1rw
* cell instance $25893 r0 *1 100.815,136.5
X$25893 352 614 353 644 645 cell_1rw
* cell instance $25894 m0 *1 100.815,139.23
X$25894 352 617 353 644 645 cell_1rw
* cell instance $25895 r0 *1 100.815,139.23
X$25895 352 616 353 644 645 cell_1rw
* cell instance $25896 m0 *1 100.815,141.96
X$25896 352 618 353 644 645 cell_1rw
* cell instance $25897 r0 *1 100.815,141.96
X$25897 352 619 353 644 645 cell_1rw
* cell instance $25898 m0 *1 100.815,144.69
X$25898 352 620 353 644 645 cell_1rw
* cell instance $25899 r0 *1 100.815,144.69
X$25899 352 621 353 644 645 cell_1rw
* cell instance $25900 m0 *1 100.815,147.42
X$25900 352 622 353 644 645 cell_1rw
* cell instance $25901 m0 *1 100.815,150.15
X$25901 352 624 353 644 645 cell_1rw
* cell instance $25902 r0 *1 100.815,147.42
X$25902 352 623 353 644 645 cell_1rw
* cell instance $25903 m0 *1 100.815,152.88
X$25903 352 626 353 644 645 cell_1rw
* cell instance $25904 r0 *1 100.815,150.15
X$25904 352 625 353 644 645 cell_1rw
* cell instance $25905 r0 *1 100.815,152.88
X$25905 352 627 353 644 645 cell_1rw
* cell instance $25906 m0 *1 100.815,155.61
X$25906 352 628 353 644 645 cell_1rw
* cell instance $25907 r0 *1 100.815,155.61
X$25907 352 629 353 644 645 cell_1rw
* cell instance $25908 m0 *1 100.815,158.34
X$25908 352 630 353 644 645 cell_1rw
* cell instance $25909 r0 *1 100.815,158.34
X$25909 352 631 353 644 645 cell_1rw
* cell instance $25910 m0 *1 100.815,161.07
X$25910 352 632 353 644 645 cell_1rw
* cell instance $25911 r0 *1 100.815,161.07
X$25911 352 633 353 644 645 cell_1rw
* cell instance $25912 m0 *1 100.815,163.8
X$25912 352 634 353 644 645 cell_1rw
* cell instance $25913 r0 *1 100.815,163.8
X$25913 352 635 353 644 645 cell_1rw
* cell instance $25914 m0 *1 100.815,166.53
X$25914 352 637 353 644 645 cell_1rw
* cell instance $25915 r0 *1 100.815,166.53
X$25915 352 636 353 644 645 cell_1rw
* cell instance $25916 m0 *1 100.815,169.26
X$25916 352 639 353 644 645 cell_1rw
* cell instance $25917 r0 *1 100.815,169.26
X$25917 352 638 353 644 645 cell_1rw
* cell instance $25918 m0 *1 100.815,171.99
X$25918 352 640 353 644 645 cell_1rw
* cell instance $25919 m0 *1 100.815,174.72
X$25919 352 642 353 644 645 cell_1rw
* cell instance $25920 r0 *1 100.815,171.99
X$25920 352 641 353 644 645 cell_1rw
* cell instance $25921 r0 *1 100.815,174.72
X$25921 352 643 353 644 645 cell_1rw
* cell instance $25922 m0 *1 101.52,90.09
X$25922 354 581 355 644 645 cell_1rw
* cell instance $25923 r0 *1 101.52,90.09
X$25923 354 580 355 644 645 cell_1rw
* cell instance $25924 m0 *1 101.52,92.82
X$25924 354 583 355 644 645 cell_1rw
* cell instance $25925 r0 *1 101.52,92.82
X$25925 354 582 355 644 645 cell_1rw
* cell instance $25926 m0 *1 101.52,95.55
X$25926 354 584 355 644 645 cell_1rw
* cell instance $25927 r0 *1 101.52,95.55
X$25927 354 585 355 644 645 cell_1rw
* cell instance $25928 m0 *1 101.52,98.28
X$25928 354 586 355 644 645 cell_1rw
* cell instance $25929 r0 *1 101.52,98.28
X$25929 354 587 355 644 645 cell_1rw
* cell instance $25930 m0 *1 101.52,101.01
X$25930 354 588 355 644 645 cell_1rw
* cell instance $25931 r0 *1 101.52,101.01
X$25931 354 589 355 644 645 cell_1rw
* cell instance $25932 m0 *1 101.52,103.74
X$25932 354 590 355 644 645 cell_1rw
* cell instance $25933 r0 *1 101.52,103.74
X$25933 354 591 355 644 645 cell_1rw
* cell instance $25934 m0 *1 101.52,106.47
X$25934 354 593 355 644 645 cell_1rw
* cell instance $25935 m0 *1 101.52,109.2
X$25935 354 594 355 644 645 cell_1rw
* cell instance $25936 r0 *1 101.52,106.47
X$25936 354 592 355 644 645 cell_1rw
* cell instance $25937 r0 *1 101.52,109.2
X$25937 354 595 355 644 645 cell_1rw
* cell instance $25938 m0 *1 101.52,111.93
X$25938 354 597 355 644 645 cell_1rw
* cell instance $25939 m0 *1 101.52,114.66
X$25939 354 598 355 644 645 cell_1rw
* cell instance $25940 r0 *1 101.52,111.93
X$25940 354 596 355 644 645 cell_1rw
* cell instance $25941 r0 *1 101.52,114.66
X$25941 354 599 355 644 645 cell_1rw
* cell instance $25942 m0 *1 101.52,117.39
X$25942 354 600 355 644 645 cell_1rw
* cell instance $25943 m0 *1 101.52,120.12
X$25943 354 602 355 644 645 cell_1rw
* cell instance $25944 r0 *1 101.52,117.39
X$25944 354 601 355 644 645 cell_1rw
* cell instance $25945 r0 *1 101.52,120.12
X$25945 354 603 355 644 645 cell_1rw
* cell instance $25946 m0 *1 101.52,122.85
X$25946 354 604 355 644 645 cell_1rw
* cell instance $25947 r0 *1 101.52,122.85
X$25947 354 605 355 644 645 cell_1rw
* cell instance $25948 m0 *1 101.52,125.58
X$25948 354 606 355 644 645 cell_1rw
* cell instance $25949 r0 *1 101.52,125.58
X$25949 354 607 355 644 645 cell_1rw
* cell instance $25950 m0 *1 101.52,128.31
X$25950 354 609 355 644 645 cell_1rw
* cell instance $25951 r0 *1 101.52,128.31
X$25951 354 608 355 644 645 cell_1rw
* cell instance $25952 m0 *1 101.52,131.04
X$25952 354 610 355 644 645 cell_1rw
* cell instance $25953 r0 *1 101.52,131.04
X$25953 354 611 355 644 645 cell_1rw
* cell instance $25954 m0 *1 101.52,133.77
X$25954 354 612 355 644 645 cell_1rw
* cell instance $25955 r0 *1 101.52,133.77
X$25955 354 613 355 644 645 cell_1rw
* cell instance $25956 m0 *1 101.52,136.5
X$25956 354 615 355 644 645 cell_1rw
* cell instance $25957 r0 *1 101.52,136.5
X$25957 354 614 355 644 645 cell_1rw
* cell instance $25958 m0 *1 101.52,139.23
X$25958 354 617 355 644 645 cell_1rw
* cell instance $25959 r0 *1 101.52,139.23
X$25959 354 616 355 644 645 cell_1rw
* cell instance $25960 m0 *1 101.52,141.96
X$25960 354 618 355 644 645 cell_1rw
* cell instance $25961 r0 *1 101.52,141.96
X$25961 354 619 355 644 645 cell_1rw
* cell instance $25962 m0 *1 101.52,144.69
X$25962 354 620 355 644 645 cell_1rw
* cell instance $25963 r0 *1 101.52,144.69
X$25963 354 621 355 644 645 cell_1rw
* cell instance $25964 m0 *1 101.52,147.42
X$25964 354 622 355 644 645 cell_1rw
* cell instance $25965 r0 *1 101.52,147.42
X$25965 354 623 355 644 645 cell_1rw
* cell instance $25966 m0 *1 101.52,150.15
X$25966 354 624 355 644 645 cell_1rw
* cell instance $25967 m0 *1 101.52,152.88
X$25967 354 626 355 644 645 cell_1rw
* cell instance $25968 r0 *1 101.52,150.15
X$25968 354 625 355 644 645 cell_1rw
* cell instance $25969 r0 *1 101.52,152.88
X$25969 354 627 355 644 645 cell_1rw
* cell instance $25970 m0 *1 101.52,155.61
X$25970 354 628 355 644 645 cell_1rw
* cell instance $25971 m0 *1 101.52,158.34
X$25971 354 630 355 644 645 cell_1rw
* cell instance $25972 r0 *1 101.52,155.61
X$25972 354 629 355 644 645 cell_1rw
* cell instance $25973 r0 *1 101.52,158.34
X$25973 354 631 355 644 645 cell_1rw
* cell instance $25974 m0 *1 101.52,161.07
X$25974 354 632 355 644 645 cell_1rw
* cell instance $25975 r0 *1 101.52,161.07
X$25975 354 633 355 644 645 cell_1rw
* cell instance $25976 m0 *1 101.52,163.8
X$25976 354 634 355 644 645 cell_1rw
* cell instance $25977 r0 *1 101.52,163.8
X$25977 354 635 355 644 645 cell_1rw
* cell instance $25978 m0 *1 101.52,166.53
X$25978 354 637 355 644 645 cell_1rw
* cell instance $25979 r0 *1 101.52,166.53
X$25979 354 636 355 644 645 cell_1rw
* cell instance $25980 m0 *1 101.52,169.26
X$25980 354 639 355 644 645 cell_1rw
* cell instance $25981 r0 *1 101.52,169.26
X$25981 354 638 355 644 645 cell_1rw
* cell instance $25982 m0 *1 101.52,171.99
X$25982 354 640 355 644 645 cell_1rw
* cell instance $25983 r0 *1 101.52,171.99
X$25983 354 641 355 644 645 cell_1rw
* cell instance $25984 m0 *1 101.52,174.72
X$25984 354 642 355 644 645 cell_1rw
* cell instance $25985 r0 *1 101.52,174.72
X$25985 354 643 355 644 645 cell_1rw
* cell instance $25986 m0 *1 102.225,90.09
X$25986 356 581 357 644 645 cell_1rw
* cell instance $25987 r0 *1 102.225,90.09
X$25987 356 580 357 644 645 cell_1rw
* cell instance $25988 m0 *1 102.225,92.82
X$25988 356 583 357 644 645 cell_1rw
* cell instance $25989 r0 *1 102.225,92.82
X$25989 356 582 357 644 645 cell_1rw
* cell instance $25990 m0 *1 102.225,95.55
X$25990 356 584 357 644 645 cell_1rw
* cell instance $25991 r0 *1 102.225,95.55
X$25991 356 585 357 644 645 cell_1rw
* cell instance $25992 m0 *1 102.225,98.28
X$25992 356 586 357 644 645 cell_1rw
* cell instance $25993 r0 *1 102.225,98.28
X$25993 356 587 357 644 645 cell_1rw
* cell instance $25994 m0 *1 102.225,101.01
X$25994 356 588 357 644 645 cell_1rw
* cell instance $25995 m0 *1 102.225,103.74
X$25995 356 590 357 644 645 cell_1rw
* cell instance $25996 r0 *1 102.225,101.01
X$25996 356 589 357 644 645 cell_1rw
* cell instance $25997 r0 *1 102.225,103.74
X$25997 356 591 357 644 645 cell_1rw
* cell instance $25998 m0 *1 102.225,106.47
X$25998 356 593 357 644 645 cell_1rw
* cell instance $25999 r0 *1 102.225,106.47
X$25999 356 592 357 644 645 cell_1rw
* cell instance $26000 m0 *1 102.225,109.2
X$26000 356 594 357 644 645 cell_1rw
* cell instance $26001 r0 *1 102.225,109.2
X$26001 356 595 357 644 645 cell_1rw
* cell instance $26002 m0 *1 102.225,111.93
X$26002 356 597 357 644 645 cell_1rw
* cell instance $26003 r0 *1 102.225,111.93
X$26003 356 596 357 644 645 cell_1rw
* cell instance $26004 m0 *1 102.225,114.66
X$26004 356 598 357 644 645 cell_1rw
* cell instance $26005 r0 *1 102.225,114.66
X$26005 356 599 357 644 645 cell_1rw
* cell instance $26006 m0 *1 102.225,117.39
X$26006 356 600 357 644 645 cell_1rw
* cell instance $26007 r0 *1 102.225,117.39
X$26007 356 601 357 644 645 cell_1rw
* cell instance $26008 m0 *1 102.225,120.12
X$26008 356 602 357 644 645 cell_1rw
* cell instance $26009 r0 *1 102.225,120.12
X$26009 356 603 357 644 645 cell_1rw
* cell instance $26010 m0 *1 102.225,122.85
X$26010 356 604 357 644 645 cell_1rw
* cell instance $26011 r0 *1 102.225,122.85
X$26011 356 605 357 644 645 cell_1rw
* cell instance $26012 m0 *1 102.225,125.58
X$26012 356 606 357 644 645 cell_1rw
* cell instance $26013 m0 *1 102.225,128.31
X$26013 356 609 357 644 645 cell_1rw
* cell instance $26014 r0 *1 102.225,125.58
X$26014 356 607 357 644 645 cell_1rw
* cell instance $26015 r0 *1 102.225,128.31
X$26015 356 608 357 644 645 cell_1rw
* cell instance $26016 m0 *1 102.225,131.04
X$26016 356 610 357 644 645 cell_1rw
* cell instance $26017 r0 *1 102.225,131.04
X$26017 356 611 357 644 645 cell_1rw
* cell instance $26018 m0 *1 102.225,133.77
X$26018 356 612 357 644 645 cell_1rw
* cell instance $26019 r0 *1 102.225,133.77
X$26019 356 613 357 644 645 cell_1rw
* cell instance $26020 m0 *1 102.225,136.5
X$26020 356 615 357 644 645 cell_1rw
* cell instance $26021 r0 *1 102.225,136.5
X$26021 356 614 357 644 645 cell_1rw
* cell instance $26022 m0 *1 102.225,139.23
X$26022 356 617 357 644 645 cell_1rw
* cell instance $26023 r0 *1 102.225,139.23
X$26023 356 616 357 644 645 cell_1rw
* cell instance $26024 m0 *1 102.225,141.96
X$26024 356 618 357 644 645 cell_1rw
* cell instance $26025 r0 *1 102.225,141.96
X$26025 356 619 357 644 645 cell_1rw
* cell instance $26026 m0 *1 102.225,144.69
X$26026 356 620 357 644 645 cell_1rw
* cell instance $26027 m0 *1 102.225,147.42
X$26027 356 622 357 644 645 cell_1rw
* cell instance $26028 r0 *1 102.225,144.69
X$26028 356 621 357 644 645 cell_1rw
* cell instance $26029 r0 *1 102.225,147.42
X$26029 356 623 357 644 645 cell_1rw
* cell instance $26030 m0 *1 102.225,150.15
X$26030 356 624 357 644 645 cell_1rw
* cell instance $26031 r0 *1 102.225,150.15
X$26031 356 625 357 644 645 cell_1rw
* cell instance $26032 m0 *1 102.225,152.88
X$26032 356 626 357 644 645 cell_1rw
* cell instance $26033 r0 *1 102.225,152.88
X$26033 356 627 357 644 645 cell_1rw
* cell instance $26034 m0 *1 102.225,155.61
X$26034 356 628 357 644 645 cell_1rw
* cell instance $26035 m0 *1 102.225,158.34
X$26035 356 630 357 644 645 cell_1rw
* cell instance $26036 r0 *1 102.225,155.61
X$26036 356 629 357 644 645 cell_1rw
* cell instance $26037 r0 *1 102.225,158.34
X$26037 356 631 357 644 645 cell_1rw
* cell instance $26038 m0 *1 102.225,161.07
X$26038 356 632 357 644 645 cell_1rw
* cell instance $26039 m0 *1 102.225,163.8
X$26039 356 634 357 644 645 cell_1rw
* cell instance $26040 r0 *1 102.225,161.07
X$26040 356 633 357 644 645 cell_1rw
* cell instance $26041 r0 *1 102.225,163.8
X$26041 356 635 357 644 645 cell_1rw
* cell instance $26042 m0 *1 102.225,166.53
X$26042 356 637 357 644 645 cell_1rw
* cell instance $26043 r0 *1 102.225,166.53
X$26043 356 636 357 644 645 cell_1rw
* cell instance $26044 m0 *1 102.225,169.26
X$26044 356 639 357 644 645 cell_1rw
* cell instance $26045 r0 *1 102.225,169.26
X$26045 356 638 357 644 645 cell_1rw
* cell instance $26046 m0 *1 102.225,171.99
X$26046 356 640 357 644 645 cell_1rw
* cell instance $26047 m0 *1 102.225,174.72
X$26047 356 642 357 644 645 cell_1rw
* cell instance $26048 r0 *1 102.225,171.99
X$26048 356 641 357 644 645 cell_1rw
* cell instance $26049 r0 *1 102.225,174.72
X$26049 356 643 357 644 645 cell_1rw
* cell instance $26050 m0 *1 102.93,90.09
X$26050 358 581 359 644 645 cell_1rw
* cell instance $26051 r0 *1 102.93,90.09
X$26051 358 580 359 644 645 cell_1rw
* cell instance $26052 m0 *1 102.93,92.82
X$26052 358 583 359 644 645 cell_1rw
* cell instance $26053 r0 *1 102.93,92.82
X$26053 358 582 359 644 645 cell_1rw
* cell instance $26054 m0 *1 102.93,95.55
X$26054 358 584 359 644 645 cell_1rw
* cell instance $26055 r0 *1 102.93,95.55
X$26055 358 585 359 644 645 cell_1rw
* cell instance $26056 m0 *1 102.93,98.28
X$26056 358 586 359 644 645 cell_1rw
* cell instance $26057 m0 *1 102.93,101.01
X$26057 358 588 359 644 645 cell_1rw
* cell instance $26058 r0 *1 102.93,98.28
X$26058 358 587 359 644 645 cell_1rw
* cell instance $26059 r0 *1 102.93,101.01
X$26059 358 589 359 644 645 cell_1rw
* cell instance $26060 m0 *1 102.93,103.74
X$26060 358 590 359 644 645 cell_1rw
* cell instance $26061 r0 *1 102.93,103.74
X$26061 358 591 359 644 645 cell_1rw
* cell instance $26062 m0 *1 102.93,106.47
X$26062 358 593 359 644 645 cell_1rw
* cell instance $26063 r0 *1 102.93,106.47
X$26063 358 592 359 644 645 cell_1rw
* cell instance $26064 m0 *1 102.93,109.2
X$26064 358 594 359 644 645 cell_1rw
* cell instance $26065 r0 *1 102.93,109.2
X$26065 358 595 359 644 645 cell_1rw
* cell instance $26066 m0 *1 102.93,111.93
X$26066 358 597 359 644 645 cell_1rw
* cell instance $26067 r0 *1 102.93,111.93
X$26067 358 596 359 644 645 cell_1rw
* cell instance $26068 m0 *1 102.93,114.66
X$26068 358 598 359 644 645 cell_1rw
* cell instance $26069 r0 *1 102.93,114.66
X$26069 358 599 359 644 645 cell_1rw
* cell instance $26070 m0 *1 102.93,117.39
X$26070 358 600 359 644 645 cell_1rw
* cell instance $26071 r0 *1 102.93,117.39
X$26071 358 601 359 644 645 cell_1rw
* cell instance $26072 m0 *1 102.93,120.12
X$26072 358 602 359 644 645 cell_1rw
* cell instance $26073 r0 *1 102.93,120.12
X$26073 358 603 359 644 645 cell_1rw
* cell instance $26074 m0 *1 102.93,122.85
X$26074 358 604 359 644 645 cell_1rw
* cell instance $26075 r0 *1 102.93,122.85
X$26075 358 605 359 644 645 cell_1rw
* cell instance $26076 m0 *1 102.93,125.58
X$26076 358 606 359 644 645 cell_1rw
* cell instance $26077 r0 *1 102.93,125.58
X$26077 358 607 359 644 645 cell_1rw
* cell instance $26078 m0 *1 102.93,128.31
X$26078 358 609 359 644 645 cell_1rw
* cell instance $26079 r0 *1 102.93,128.31
X$26079 358 608 359 644 645 cell_1rw
* cell instance $26080 m0 *1 102.93,131.04
X$26080 358 610 359 644 645 cell_1rw
* cell instance $26081 r0 *1 102.93,131.04
X$26081 358 611 359 644 645 cell_1rw
* cell instance $26082 m0 *1 102.93,133.77
X$26082 358 612 359 644 645 cell_1rw
* cell instance $26083 r0 *1 102.93,133.77
X$26083 358 613 359 644 645 cell_1rw
* cell instance $26084 m0 *1 102.93,136.5
X$26084 358 615 359 644 645 cell_1rw
* cell instance $26085 r0 *1 102.93,136.5
X$26085 358 614 359 644 645 cell_1rw
* cell instance $26086 m0 *1 102.93,139.23
X$26086 358 617 359 644 645 cell_1rw
* cell instance $26087 m0 *1 102.93,141.96
X$26087 358 618 359 644 645 cell_1rw
* cell instance $26088 r0 *1 102.93,139.23
X$26088 358 616 359 644 645 cell_1rw
* cell instance $26089 r0 *1 102.93,141.96
X$26089 358 619 359 644 645 cell_1rw
* cell instance $26090 m0 *1 102.93,144.69
X$26090 358 620 359 644 645 cell_1rw
* cell instance $26091 r0 *1 102.93,144.69
X$26091 358 621 359 644 645 cell_1rw
* cell instance $26092 m0 *1 102.93,147.42
X$26092 358 622 359 644 645 cell_1rw
* cell instance $26093 m0 *1 102.93,150.15
X$26093 358 624 359 644 645 cell_1rw
* cell instance $26094 r0 *1 102.93,147.42
X$26094 358 623 359 644 645 cell_1rw
* cell instance $26095 r0 *1 102.93,150.15
X$26095 358 625 359 644 645 cell_1rw
* cell instance $26096 m0 *1 102.93,152.88
X$26096 358 626 359 644 645 cell_1rw
* cell instance $26097 r0 *1 102.93,152.88
X$26097 358 627 359 644 645 cell_1rw
* cell instance $26098 m0 *1 102.93,155.61
X$26098 358 628 359 644 645 cell_1rw
* cell instance $26099 m0 *1 102.93,158.34
X$26099 358 630 359 644 645 cell_1rw
* cell instance $26100 r0 *1 102.93,155.61
X$26100 358 629 359 644 645 cell_1rw
* cell instance $26101 r0 *1 102.93,158.34
X$26101 358 631 359 644 645 cell_1rw
* cell instance $26102 m0 *1 102.93,161.07
X$26102 358 632 359 644 645 cell_1rw
* cell instance $26103 m0 *1 102.93,163.8
X$26103 358 634 359 644 645 cell_1rw
* cell instance $26104 r0 *1 102.93,161.07
X$26104 358 633 359 644 645 cell_1rw
* cell instance $26105 r0 *1 102.93,163.8
X$26105 358 635 359 644 645 cell_1rw
* cell instance $26106 m0 *1 102.93,166.53
X$26106 358 637 359 644 645 cell_1rw
* cell instance $26107 r0 *1 102.93,166.53
X$26107 358 636 359 644 645 cell_1rw
* cell instance $26108 m0 *1 102.93,169.26
X$26108 358 639 359 644 645 cell_1rw
* cell instance $26109 r0 *1 102.93,169.26
X$26109 358 638 359 644 645 cell_1rw
* cell instance $26110 m0 *1 102.93,171.99
X$26110 358 640 359 644 645 cell_1rw
* cell instance $26111 r0 *1 102.93,171.99
X$26111 358 641 359 644 645 cell_1rw
* cell instance $26112 m0 *1 102.93,174.72
X$26112 358 642 359 644 645 cell_1rw
* cell instance $26113 r0 *1 102.93,174.72
X$26113 358 643 359 644 645 cell_1rw
* cell instance $26114 m0 *1 103.635,90.09
X$26114 360 581 361 644 645 cell_1rw
* cell instance $26115 r0 *1 103.635,90.09
X$26115 360 580 361 644 645 cell_1rw
* cell instance $26116 m0 *1 103.635,92.82
X$26116 360 583 361 644 645 cell_1rw
* cell instance $26117 r0 *1 103.635,92.82
X$26117 360 582 361 644 645 cell_1rw
* cell instance $26118 m0 *1 103.635,95.55
X$26118 360 584 361 644 645 cell_1rw
* cell instance $26119 m0 *1 103.635,98.28
X$26119 360 586 361 644 645 cell_1rw
* cell instance $26120 r0 *1 103.635,95.55
X$26120 360 585 361 644 645 cell_1rw
* cell instance $26121 r0 *1 103.635,98.28
X$26121 360 587 361 644 645 cell_1rw
* cell instance $26122 m0 *1 103.635,101.01
X$26122 360 588 361 644 645 cell_1rw
* cell instance $26123 r0 *1 103.635,101.01
X$26123 360 589 361 644 645 cell_1rw
* cell instance $26124 m0 *1 103.635,103.74
X$26124 360 590 361 644 645 cell_1rw
* cell instance $26125 r0 *1 103.635,103.74
X$26125 360 591 361 644 645 cell_1rw
* cell instance $26126 m0 *1 103.635,106.47
X$26126 360 593 361 644 645 cell_1rw
* cell instance $26127 m0 *1 103.635,109.2
X$26127 360 594 361 644 645 cell_1rw
* cell instance $26128 r0 *1 103.635,106.47
X$26128 360 592 361 644 645 cell_1rw
* cell instance $26129 r0 *1 103.635,109.2
X$26129 360 595 361 644 645 cell_1rw
* cell instance $26130 m0 *1 103.635,111.93
X$26130 360 597 361 644 645 cell_1rw
* cell instance $26131 r0 *1 103.635,111.93
X$26131 360 596 361 644 645 cell_1rw
* cell instance $26132 m0 *1 103.635,114.66
X$26132 360 598 361 644 645 cell_1rw
* cell instance $26133 r0 *1 103.635,114.66
X$26133 360 599 361 644 645 cell_1rw
* cell instance $26134 m0 *1 103.635,117.39
X$26134 360 600 361 644 645 cell_1rw
* cell instance $26135 r0 *1 103.635,117.39
X$26135 360 601 361 644 645 cell_1rw
* cell instance $26136 m0 *1 103.635,120.12
X$26136 360 602 361 644 645 cell_1rw
* cell instance $26137 r0 *1 103.635,120.12
X$26137 360 603 361 644 645 cell_1rw
* cell instance $26138 m0 *1 103.635,122.85
X$26138 360 604 361 644 645 cell_1rw
* cell instance $26139 r0 *1 103.635,122.85
X$26139 360 605 361 644 645 cell_1rw
* cell instance $26140 m0 *1 103.635,125.58
X$26140 360 606 361 644 645 cell_1rw
* cell instance $26141 r0 *1 103.635,125.58
X$26141 360 607 361 644 645 cell_1rw
* cell instance $26142 m0 *1 103.635,128.31
X$26142 360 609 361 644 645 cell_1rw
* cell instance $26143 r0 *1 103.635,128.31
X$26143 360 608 361 644 645 cell_1rw
* cell instance $26144 m0 *1 103.635,131.04
X$26144 360 610 361 644 645 cell_1rw
* cell instance $26145 r0 *1 103.635,131.04
X$26145 360 611 361 644 645 cell_1rw
* cell instance $26146 m0 *1 103.635,133.77
X$26146 360 612 361 644 645 cell_1rw
* cell instance $26147 m0 *1 103.635,136.5
X$26147 360 615 361 644 645 cell_1rw
* cell instance $26148 r0 *1 103.635,133.77
X$26148 360 613 361 644 645 cell_1rw
* cell instance $26149 r0 *1 103.635,136.5
X$26149 360 614 361 644 645 cell_1rw
* cell instance $26150 m0 *1 103.635,139.23
X$26150 360 617 361 644 645 cell_1rw
* cell instance $26151 r0 *1 103.635,139.23
X$26151 360 616 361 644 645 cell_1rw
* cell instance $26152 m0 *1 103.635,141.96
X$26152 360 618 361 644 645 cell_1rw
* cell instance $26153 r0 *1 103.635,141.96
X$26153 360 619 361 644 645 cell_1rw
* cell instance $26154 m0 *1 103.635,144.69
X$26154 360 620 361 644 645 cell_1rw
* cell instance $26155 r0 *1 103.635,144.69
X$26155 360 621 361 644 645 cell_1rw
* cell instance $26156 m0 *1 103.635,147.42
X$26156 360 622 361 644 645 cell_1rw
* cell instance $26157 m0 *1 103.635,150.15
X$26157 360 624 361 644 645 cell_1rw
* cell instance $26158 r0 *1 103.635,147.42
X$26158 360 623 361 644 645 cell_1rw
* cell instance $26159 r0 *1 103.635,150.15
X$26159 360 625 361 644 645 cell_1rw
* cell instance $26160 m0 *1 103.635,152.88
X$26160 360 626 361 644 645 cell_1rw
* cell instance $26161 r0 *1 103.635,152.88
X$26161 360 627 361 644 645 cell_1rw
* cell instance $26162 m0 *1 103.635,155.61
X$26162 360 628 361 644 645 cell_1rw
* cell instance $26163 r0 *1 103.635,155.61
X$26163 360 629 361 644 645 cell_1rw
* cell instance $26164 m0 *1 103.635,158.34
X$26164 360 630 361 644 645 cell_1rw
* cell instance $26165 r0 *1 103.635,158.34
X$26165 360 631 361 644 645 cell_1rw
* cell instance $26166 m0 *1 103.635,161.07
X$26166 360 632 361 644 645 cell_1rw
* cell instance $26167 r0 *1 103.635,161.07
X$26167 360 633 361 644 645 cell_1rw
* cell instance $26168 m0 *1 103.635,163.8
X$26168 360 634 361 644 645 cell_1rw
* cell instance $26169 r0 *1 103.635,163.8
X$26169 360 635 361 644 645 cell_1rw
* cell instance $26170 m0 *1 103.635,166.53
X$26170 360 637 361 644 645 cell_1rw
* cell instance $26171 r0 *1 103.635,166.53
X$26171 360 636 361 644 645 cell_1rw
* cell instance $26172 m0 *1 103.635,169.26
X$26172 360 639 361 644 645 cell_1rw
* cell instance $26173 r0 *1 103.635,169.26
X$26173 360 638 361 644 645 cell_1rw
* cell instance $26174 m0 *1 103.635,171.99
X$26174 360 640 361 644 645 cell_1rw
* cell instance $26175 r0 *1 103.635,171.99
X$26175 360 641 361 644 645 cell_1rw
* cell instance $26176 m0 *1 103.635,174.72
X$26176 360 642 361 644 645 cell_1rw
* cell instance $26177 r0 *1 103.635,174.72
X$26177 360 643 361 644 645 cell_1rw
* cell instance $26178 m0 *1 104.34,90.09
X$26178 362 581 363 644 645 cell_1rw
* cell instance $26179 r0 *1 104.34,90.09
X$26179 362 580 363 644 645 cell_1rw
* cell instance $26180 m0 *1 104.34,92.82
X$26180 362 583 363 644 645 cell_1rw
* cell instance $26181 r0 *1 104.34,92.82
X$26181 362 582 363 644 645 cell_1rw
* cell instance $26182 m0 *1 104.34,95.55
X$26182 362 584 363 644 645 cell_1rw
* cell instance $26183 r0 *1 104.34,95.55
X$26183 362 585 363 644 645 cell_1rw
* cell instance $26184 m0 *1 104.34,98.28
X$26184 362 586 363 644 645 cell_1rw
* cell instance $26185 r0 *1 104.34,98.28
X$26185 362 587 363 644 645 cell_1rw
* cell instance $26186 m0 *1 104.34,101.01
X$26186 362 588 363 644 645 cell_1rw
* cell instance $26187 r0 *1 104.34,101.01
X$26187 362 589 363 644 645 cell_1rw
* cell instance $26188 m0 *1 104.34,103.74
X$26188 362 590 363 644 645 cell_1rw
* cell instance $26189 r0 *1 104.34,103.74
X$26189 362 591 363 644 645 cell_1rw
* cell instance $26190 m0 *1 104.34,106.47
X$26190 362 593 363 644 645 cell_1rw
* cell instance $26191 m0 *1 104.34,109.2
X$26191 362 594 363 644 645 cell_1rw
* cell instance $26192 r0 *1 104.34,106.47
X$26192 362 592 363 644 645 cell_1rw
* cell instance $26193 r0 *1 104.34,109.2
X$26193 362 595 363 644 645 cell_1rw
* cell instance $26194 m0 *1 104.34,111.93
X$26194 362 597 363 644 645 cell_1rw
* cell instance $26195 r0 *1 104.34,111.93
X$26195 362 596 363 644 645 cell_1rw
* cell instance $26196 m0 *1 104.34,114.66
X$26196 362 598 363 644 645 cell_1rw
* cell instance $26197 r0 *1 104.34,114.66
X$26197 362 599 363 644 645 cell_1rw
* cell instance $26198 m0 *1 104.34,117.39
X$26198 362 600 363 644 645 cell_1rw
* cell instance $26199 r0 *1 104.34,117.39
X$26199 362 601 363 644 645 cell_1rw
* cell instance $26200 m0 *1 104.34,120.12
X$26200 362 602 363 644 645 cell_1rw
* cell instance $26201 r0 *1 104.34,120.12
X$26201 362 603 363 644 645 cell_1rw
* cell instance $26202 m0 *1 104.34,122.85
X$26202 362 604 363 644 645 cell_1rw
* cell instance $26203 m0 *1 104.34,125.58
X$26203 362 606 363 644 645 cell_1rw
* cell instance $26204 r0 *1 104.34,122.85
X$26204 362 605 363 644 645 cell_1rw
* cell instance $26205 r0 *1 104.34,125.58
X$26205 362 607 363 644 645 cell_1rw
* cell instance $26206 m0 *1 104.34,128.31
X$26206 362 609 363 644 645 cell_1rw
* cell instance $26207 m0 *1 104.34,131.04
X$26207 362 610 363 644 645 cell_1rw
* cell instance $26208 r0 *1 104.34,128.31
X$26208 362 608 363 644 645 cell_1rw
* cell instance $26209 r0 *1 104.34,131.04
X$26209 362 611 363 644 645 cell_1rw
* cell instance $26210 m0 *1 104.34,133.77
X$26210 362 612 363 644 645 cell_1rw
* cell instance $26211 m0 *1 104.34,136.5
X$26211 362 615 363 644 645 cell_1rw
* cell instance $26212 r0 *1 104.34,133.77
X$26212 362 613 363 644 645 cell_1rw
* cell instance $26213 r0 *1 104.34,136.5
X$26213 362 614 363 644 645 cell_1rw
* cell instance $26214 m0 *1 104.34,139.23
X$26214 362 617 363 644 645 cell_1rw
* cell instance $26215 r0 *1 104.34,139.23
X$26215 362 616 363 644 645 cell_1rw
* cell instance $26216 m0 *1 104.34,141.96
X$26216 362 618 363 644 645 cell_1rw
* cell instance $26217 r0 *1 104.34,141.96
X$26217 362 619 363 644 645 cell_1rw
* cell instance $26218 m0 *1 104.34,144.69
X$26218 362 620 363 644 645 cell_1rw
* cell instance $26219 r0 *1 104.34,144.69
X$26219 362 621 363 644 645 cell_1rw
* cell instance $26220 m0 *1 104.34,147.42
X$26220 362 622 363 644 645 cell_1rw
* cell instance $26221 r0 *1 104.34,147.42
X$26221 362 623 363 644 645 cell_1rw
* cell instance $26222 m0 *1 104.34,150.15
X$26222 362 624 363 644 645 cell_1rw
* cell instance $26223 r0 *1 104.34,150.15
X$26223 362 625 363 644 645 cell_1rw
* cell instance $26224 m0 *1 104.34,152.88
X$26224 362 626 363 644 645 cell_1rw
* cell instance $26225 r0 *1 104.34,152.88
X$26225 362 627 363 644 645 cell_1rw
* cell instance $26226 m0 *1 104.34,155.61
X$26226 362 628 363 644 645 cell_1rw
* cell instance $26227 r0 *1 104.34,155.61
X$26227 362 629 363 644 645 cell_1rw
* cell instance $26228 m0 *1 104.34,158.34
X$26228 362 630 363 644 645 cell_1rw
* cell instance $26229 m0 *1 104.34,161.07
X$26229 362 632 363 644 645 cell_1rw
* cell instance $26230 r0 *1 104.34,158.34
X$26230 362 631 363 644 645 cell_1rw
* cell instance $26231 m0 *1 104.34,163.8
X$26231 362 634 363 644 645 cell_1rw
* cell instance $26232 r0 *1 104.34,161.07
X$26232 362 633 363 644 645 cell_1rw
* cell instance $26233 r0 *1 104.34,163.8
X$26233 362 635 363 644 645 cell_1rw
* cell instance $26234 m0 *1 104.34,166.53
X$26234 362 637 363 644 645 cell_1rw
* cell instance $26235 r0 *1 104.34,166.53
X$26235 362 636 363 644 645 cell_1rw
* cell instance $26236 m0 *1 104.34,169.26
X$26236 362 639 363 644 645 cell_1rw
* cell instance $26237 m0 *1 104.34,171.99
X$26237 362 640 363 644 645 cell_1rw
* cell instance $26238 r0 *1 104.34,169.26
X$26238 362 638 363 644 645 cell_1rw
* cell instance $26239 r0 *1 104.34,171.99
X$26239 362 641 363 644 645 cell_1rw
* cell instance $26240 m0 *1 104.34,174.72
X$26240 362 642 363 644 645 cell_1rw
* cell instance $26241 r0 *1 104.34,174.72
X$26241 362 643 363 644 645 cell_1rw
* cell instance $26242 m0 *1 105.045,90.09
X$26242 364 581 365 644 645 cell_1rw
* cell instance $26243 r0 *1 105.045,90.09
X$26243 364 580 365 644 645 cell_1rw
* cell instance $26244 m0 *1 105.045,92.82
X$26244 364 583 365 644 645 cell_1rw
* cell instance $26245 r0 *1 105.045,92.82
X$26245 364 582 365 644 645 cell_1rw
* cell instance $26246 m0 *1 105.045,95.55
X$26246 364 584 365 644 645 cell_1rw
* cell instance $26247 m0 *1 105.045,98.28
X$26247 364 586 365 644 645 cell_1rw
* cell instance $26248 r0 *1 105.045,95.55
X$26248 364 585 365 644 645 cell_1rw
* cell instance $26249 r0 *1 105.045,98.28
X$26249 364 587 365 644 645 cell_1rw
* cell instance $26250 m0 *1 105.045,101.01
X$26250 364 588 365 644 645 cell_1rw
* cell instance $26251 r0 *1 105.045,101.01
X$26251 364 589 365 644 645 cell_1rw
* cell instance $26252 m0 *1 105.045,103.74
X$26252 364 590 365 644 645 cell_1rw
* cell instance $26253 r0 *1 105.045,103.74
X$26253 364 591 365 644 645 cell_1rw
* cell instance $26254 m0 *1 105.045,106.47
X$26254 364 593 365 644 645 cell_1rw
* cell instance $26255 m0 *1 105.045,109.2
X$26255 364 594 365 644 645 cell_1rw
* cell instance $26256 r0 *1 105.045,106.47
X$26256 364 592 365 644 645 cell_1rw
* cell instance $26257 m0 *1 105.045,111.93
X$26257 364 597 365 644 645 cell_1rw
* cell instance $26258 r0 *1 105.045,109.2
X$26258 364 595 365 644 645 cell_1rw
* cell instance $26259 m0 *1 105.045,114.66
X$26259 364 598 365 644 645 cell_1rw
* cell instance $26260 r0 *1 105.045,111.93
X$26260 364 596 365 644 645 cell_1rw
* cell instance $26261 r0 *1 105.045,114.66
X$26261 364 599 365 644 645 cell_1rw
* cell instance $26262 m0 *1 105.045,117.39
X$26262 364 600 365 644 645 cell_1rw
* cell instance $26263 r0 *1 105.045,117.39
X$26263 364 601 365 644 645 cell_1rw
* cell instance $26264 m0 *1 105.045,120.12
X$26264 364 602 365 644 645 cell_1rw
* cell instance $26265 r0 *1 105.045,120.12
X$26265 364 603 365 644 645 cell_1rw
* cell instance $26266 m0 *1 105.045,122.85
X$26266 364 604 365 644 645 cell_1rw
* cell instance $26267 r0 *1 105.045,122.85
X$26267 364 605 365 644 645 cell_1rw
* cell instance $26268 m0 *1 105.045,125.58
X$26268 364 606 365 644 645 cell_1rw
* cell instance $26269 r0 *1 105.045,125.58
X$26269 364 607 365 644 645 cell_1rw
* cell instance $26270 m0 *1 105.045,128.31
X$26270 364 609 365 644 645 cell_1rw
* cell instance $26271 r0 *1 105.045,128.31
X$26271 364 608 365 644 645 cell_1rw
* cell instance $26272 m0 *1 105.045,131.04
X$26272 364 610 365 644 645 cell_1rw
* cell instance $26273 r0 *1 105.045,131.04
X$26273 364 611 365 644 645 cell_1rw
* cell instance $26274 m0 *1 105.045,133.77
X$26274 364 612 365 644 645 cell_1rw
* cell instance $26275 r0 *1 105.045,133.77
X$26275 364 613 365 644 645 cell_1rw
* cell instance $26276 m0 *1 105.045,136.5
X$26276 364 615 365 644 645 cell_1rw
* cell instance $26277 r0 *1 105.045,136.5
X$26277 364 614 365 644 645 cell_1rw
* cell instance $26278 m0 *1 105.045,139.23
X$26278 364 617 365 644 645 cell_1rw
* cell instance $26279 r0 *1 105.045,139.23
X$26279 364 616 365 644 645 cell_1rw
* cell instance $26280 m0 *1 105.045,141.96
X$26280 364 618 365 644 645 cell_1rw
* cell instance $26281 m0 *1 105.045,144.69
X$26281 364 620 365 644 645 cell_1rw
* cell instance $26282 r0 *1 105.045,141.96
X$26282 364 619 365 644 645 cell_1rw
* cell instance $26283 m0 *1 105.045,147.42
X$26283 364 622 365 644 645 cell_1rw
* cell instance $26284 r0 *1 105.045,144.69
X$26284 364 621 365 644 645 cell_1rw
* cell instance $26285 r0 *1 105.045,147.42
X$26285 364 623 365 644 645 cell_1rw
* cell instance $26286 m0 *1 105.045,150.15
X$26286 364 624 365 644 645 cell_1rw
* cell instance $26287 r0 *1 105.045,150.15
X$26287 364 625 365 644 645 cell_1rw
* cell instance $26288 m0 *1 105.045,152.88
X$26288 364 626 365 644 645 cell_1rw
* cell instance $26289 r0 *1 105.045,152.88
X$26289 364 627 365 644 645 cell_1rw
* cell instance $26290 m0 *1 105.045,155.61
X$26290 364 628 365 644 645 cell_1rw
* cell instance $26291 r0 *1 105.045,155.61
X$26291 364 629 365 644 645 cell_1rw
* cell instance $26292 m0 *1 105.045,158.34
X$26292 364 630 365 644 645 cell_1rw
* cell instance $26293 r0 *1 105.045,158.34
X$26293 364 631 365 644 645 cell_1rw
* cell instance $26294 m0 *1 105.045,161.07
X$26294 364 632 365 644 645 cell_1rw
* cell instance $26295 r0 *1 105.045,161.07
X$26295 364 633 365 644 645 cell_1rw
* cell instance $26296 m0 *1 105.045,163.8
X$26296 364 634 365 644 645 cell_1rw
* cell instance $26297 r0 *1 105.045,163.8
X$26297 364 635 365 644 645 cell_1rw
* cell instance $26298 m0 *1 105.045,166.53
X$26298 364 637 365 644 645 cell_1rw
* cell instance $26299 r0 *1 105.045,166.53
X$26299 364 636 365 644 645 cell_1rw
* cell instance $26300 m0 *1 105.045,169.26
X$26300 364 639 365 644 645 cell_1rw
* cell instance $26301 r0 *1 105.045,169.26
X$26301 364 638 365 644 645 cell_1rw
* cell instance $26302 m0 *1 105.045,171.99
X$26302 364 640 365 644 645 cell_1rw
* cell instance $26303 m0 *1 105.045,174.72
X$26303 364 642 365 644 645 cell_1rw
* cell instance $26304 r0 *1 105.045,171.99
X$26304 364 641 365 644 645 cell_1rw
* cell instance $26305 r0 *1 105.045,174.72
X$26305 364 643 365 644 645 cell_1rw
* cell instance $26306 m0 *1 105.75,90.09
X$26306 366 581 367 644 645 cell_1rw
* cell instance $26307 r0 *1 105.75,90.09
X$26307 366 580 367 644 645 cell_1rw
* cell instance $26308 m0 *1 105.75,92.82
X$26308 366 583 367 644 645 cell_1rw
* cell instance $26309 r0 *1 105.75,92.82
X$26309 366 582 367 644 645 cell_1rw
* cell instance $26310 m0 *1 105.75,95.55
X$26310 366 584 367 644 645 cell_1rw
* cell instance $26311 r0 *1 105.75,95.55
X$26311 366 585 367 644 645 cell_1rw
* cell instance $26312 m0 *1 105.75,98.28
X$26312 366 586 367 644 645 cell_1rw
* cell instance $26313 m0 *1 105.75,101.01
X$26313 366 588 367 644 645 cell_1rw
* cell instance $26314 r0 *1 105.75,98.28
X$26314 366 587 367 644 645 cell_1rw
* cell instance $26315 m0 *1 105.75,103.74
X$26315 366 590 367 644 645 cell_1rw
* cell instance $26316 r0 *1 105.75,101.01
X$26316 366 589 367 644 645 cell_1rw
* cell instance $26317 r0 *1 105.75,103.74
X$26317 366 591 367 644 645 cell_1rw
* cell instance $26318 m0 *1 105.75,106.47
X$26318 366 593 367 644 645 cell_1rw
* cell instance $26319 r0 *1 105.75,106.47
X$26319 366 592 367 644 645 cell_1rw
* cell instance $26320 m0 *1 105.75,109.2
X$26320 366 594 367 644 645 cell_1rw
* cell instance $26321 r0 *1 105.75,109.2
X$26321 366 595 367 644 645 cell_1rw
* cell instance $26322 m0 *1 105.75,111.93
X$26322 366 597 367 644 645 cell_1rw
* cell instance $26323 m0 *1 105.75,114.66
X$26323 366 598 367 644 645 cell_1rw
* cell instance $26324 r0 *1 105.75,111.93
X$26324 366 596 367 644 645 cell_1rw
* cell instance $26325 r0 *1 105.75,114.66
X$26325 366 599 367 644 645 cell_1rw
* cell instance $26326 m0 *1 105.75,117.39
X$26326 366 600 367 644 645 cell_1rw
* cell instance $26327 r0 *1 105.75,117.39
X$26327 366 601 367 644 645 cell_1rw
* cell instance $26328 m0 *1 105.75,120.12
X$26328 366 602 367 644 645 cell_1rw
* cell instance $26329 r0 *1 105.75,120.12
X$26329 366 603 367 644 645 cell_1rw
* cell instance $26330 m0 *1 105.75,122.85
X$26330 366 604 367 644 645 cell_1rw
* cell instance $26331 r0 *1 105.75,122.85
X$26331 366 605 367 644 645 cell_1rw
* cell instance $26332 m0 *1 105.75,125.58
X$26332 366 606 367 644 645 cell_1rw
* cell instance $26333 r0 *1 105.75,125.58
X$26333 366 607 367 644 645 cell_1rw
* cell instance $26334 m0 *1 105.75,128.31
X$26334 366 609 367 644 645 cell_1rw
* cell instance $26335 r0 *1 105.75,128.31
X$26335 366 608 367 644 645 cell_1rw
* cell instance $26336 m0 *1 105.75,131.04
X$26336 366 610 367 644 645 cell_1rw
* cell instance $26337 r0 *1 105.75,131.04
X$26337 366 611 367 644 645 cell_1rw
* cell instance $26338 m0 *1 105.75,133.77
X$26338 366 612 367 644 645 cell_1rw
* cell instance $26339 m0 *1 105.75,136.5
X$26339 366 615 367 644 645 cell_1rw
* cell instance $26340 r0 *1 105.75,133.77
X$26340 366 613 367 644 645 cell_1rw
* cell instance $26341 r0 *1 105.75,136.5
X$26341 366 614 367 644 645 cell_1rw
* cell instance $26342 m0 *1 105.75,139.23
X$26342 366 617 367 644 645 cell_1rw
* cell instance $26343 m0 *1 105.75,141.96
X$26343 366 618 367 644 645 cell_1rw
* cell instance $26344 r0 *1 105.75,139.23
X$26344 366 616 367 644 645 cell_1rw
* cell instance $26345 r0 *1 105.75,141.96
X$26345 366 619 367 644 645 cell_1rw
* cell instance $26346 m0 *1 105.75,144.69
X$26346 366 620 367 644 645 cell_1rw
* cell instance $26347 r0 *1 105.75,144.69
X$26347 366 621 367 644 645 cell_1rw
* cell instance $26348 m0 *1 105.75,147.42
X$26348 366 622 367 644 645 cell_1rw
* cell instance $26349 r0 *1 105.75,147.42
X$26349 366 623 367 644 645 cell_1rw
* cell instance $26350 m0 *1 105.75,150.15
X$26350 366 624 367 644 645 cell_1rw
* cell instance $26351 r0 *1 105.75,150.15
X$26351 366 625 367 644 645 cell_1rw
* cell instance $26352 m0 *1 105.75,152.88
X$26352 366 626 367 644 645 cell_1rw
* cell instance $26353 r0 *1 105.75,152.88
X$26353 366 627 367 644 645 cell_1rw
* cell instance $26354 m0 *1 105.75,155.61
X$26354 366 628 367 644 645 cell_1rw
* cell instance $26355 r0 *1 105.75,155.61
X$26355 366 629 367 644 645 cell_1rw
* cell instance $26356 m0 *1 105.75,158.34
X$26356 366 630 367 644 645 cell_1rw
* cell instance $26357 r0 *1 105.75,158.34
X$26357 366 631 367 644 645 cell_1rw
* cell instance $26358 m0 *1 105.75,161.07
X$26358 366 632 367 644 645 cell_1rw
* cell instance $26359 r0 *1 105.75,161.07
X$26359 366 633 367 644 645 cell_1rw
* cell instance $26360 m0 *1 105.75,163.8
X$26360 366 634 367 644 645 cell_1rw
* cell instance $26361 m0 *1 105.75,166.53
X$26361 366 637 367 644 645 cell_1rw
* cell instance $26362 r0 *1 105.75,163.8
X$26362 366 635 367 644 645 cell_1rw
* cell instance $26363 r0 *1 105.75,166.53
X$26363 366 636 367 644 645 cell_1rw
* cell instance $26364 m0 *1 105.75,169.26
X$26364 366 639 367 644 645 cell_1rw
* cell instance $26365 r0 *1 105.75,169.26
X$26365 366 638 367 644 645 cell_1rw
* cell instance $26366 m0 *1 105.75,171.99
X$26366 366 640 367 644 645 cell_1rw
* cell instance $26367 r0 *1 105.75,171.99
X$26367 366 641 367 644 645 cell_1rw
* cell instance $26368 m0 *1 105.75,174.72
X$26368 366 642 367 644 645 cell_1rw
* cell instance $26369 r0 *1 105.75,174.72
X$26369 366 643 367 644 645 cell_1rw
* cell instance $26370 m0 *1 106.455,90.09
X$26370 368 581 369 644 645 cell_1rw
* cell instance $26371 r0 *1 106.455,90.09
X$26371 368 580 369 644 645 cell_1rw
* cell instance $26372 m0 *1 106.455,92.82
X$26372 368 583 369 644 645 cell_1rw
* cell instance $26373 r0 *1 106.455,92.82
X$26373 368 582 369 644 645 cell_1rw
* cell instance $26374 m0 *1 106.455,95.55
X$26374 368 584 369 644 645 cell_1rw
* cell instance $26375 r0 *1 106.455,95.55
X$26375 368 585 369 644 645 cell_1rw
* cell instance $26376 m0 *1 106.455,98.28
X$26376 368 586 369 644 645 cell_1rw
* cell instance $26377 r0 *1 106.455,98.28
X$26377 368 587 369 644 645 cell_1rw
* cell instance $26378 m0 *1 106.455,101.01
X$26378 368 588 369 644 645 cell_1rw
* cell instance $26379 r0 *1 106.455,101.01
X$26379 368 589 369 644 645 cell_1rw
* cell instance $26380 m0 *1 106.455,103.74
X$26380 368 590 369 644 645 cell_1rw
* cell instance $26381 m0 *1 106.455,106.47
X$26381 368 593 369 644 645 cell_1rw
* cell instance $26382 r0 *1 106.455,103.74
X$26382 368 591 369 644 645 cell_1rw
* cell instance $26383 r0 *1 106.455,106.47
X$26383 368 592 369 644 645 cell_1rw
* cell instance $26384 m0 *1 106.455,109.2
X$26384 368 594 369 644 645 cell_1rw
* cell instance $26385 r0 *1 106.455,109.2
X$26385 368 595 369 644 645 cell_1rw
* cell instance $26386 m0 *1 106.455,111.93
X$26386 368 597 369 644 645 cell_1rw
* cell instance $26387 r0 *1 106.455,111.93
X$26387 368 596 369 644 645 cell_1rw
* cell instance $26388 m0 *1 106.455,114.66
X$26388 368 598 369 644 645 cell_1rw
* cell instance $26389 r0 *1 106.455,114.66
X$26389 368 599 369 644 645 cell_1rw
* cell instance $26390 m0 *1 106.455,117.39
X$26390 368 600 369 644 645 cell_1rw
* cell instance $26391 r0 *1 106.455,117.39
X$26391 368 601 369 644 645 cell_1rw
* cell instance $26392 m0 *1 106.455,120.12
X$26392 368 602 369 644 645 cell_1rw
* cell instance $26393 r0 *1 106.455,120.12
X$26393 368 603 369 644 645 cell_1rw
* cell instance $26394 m0 *1 106.455,122.85
X$26394 368 604 369 644 645 cell_1rw
* cell instance $26395 r0 *1 106.455,122.85
X$26395 368 605 369 644 645 cell_1rw
* cell instance $26396 m0 *1 106.455,125.58
X$26396 368 606 369 644 645 cell_1rw
* cell instance $26397 m0 *1 106.455,128.31
X$26397 368 609 369 644 645 cell_1rw
* cell instance $26398 r0 *1 106.455,125.58
X$26398 368 607 369 644 645 cell_1rw
* cell instance $26399 r0 *1 106.455,128.31
X$26399 368 608 369 644 645 cell_1rw
* cell instance $26400 m0 *1 106.455,131.04
X$26400 368 610 369 644 645 cell_1rw
* cell instance $26401 r0 *1 106.455,131.04
X$26401 368 611 369 644 645 cell_1rw
* cell instance $26402 m0 *1 106.455,133.77
X$26402 368 612 369 644 645 cell_1rw
* cell instance $26403 r0 *1 106.455,133.77
X$26403 368 613 369 644 645 cell_1rw
* cell instance $26404 m0 *1 106.455,136.5
X$26404 368 615 369 644 645 cell_1rw
* cell instance $26405 r0 *1 106.455,136.5
X$26405 368 614 369 644 645 cell_1rw
* cell instance $26406 m0 *1 106.455,139.23
X$26406 368 617 369 644 645 cell_1rw
* cell instance $26407 r0 *1 106.455,139.23
X$26407 368 616 369 644 645 cell_1rw
* cell instance $26408 m0 *1 106.455,141.96
X$26408 368 618 369 644 645 cell_1rw
* cell instance $26409 r0 *1 106.455,141.96
X$26409 368 619 369 644 645 cell_1rw
* cell instance $26410 m0 *1 106.455,144.69
X$26410 368 620 369 644 645 cell_1rw
* cell instance $26411 r0 *1 106.455,144.69
X$26411 368 621 369 644 645 cell_1rw
* cell instance $26412 m0 *1 106.455,147.42
X$26412 368 622 369 644 645 cell_1rw
* cell instance $26413 m0 *1 106.455,150.15
X$26413 368 624 369 644 645 cell_1rw
* cell instance $26414 r0 *1 106.455,147.42
X$26414 368 623 369 644 645 cell_1rw
* cell instance $26415 m0 *1 106.455,152.88
X$26415 368 626 369 644 645 cell_1rw
* cell instance $26416 r0 *1 106.455,150.15
X$26416 368 625 369 644 645 cell_1rw
* cell instance $26417 m0 *1 106.455,155.61
X$26417 368 628 369 644 645 cell_1rw
* cell instance $26418 r0 *1 106.455,152.88
X$26418 368 627 369 644 645 cell_1rw
* cell instance $26419 r0 *1 106.455,155.61
X$26419 368 629 369 644 645 cell_1rw
* cell instance $26420 m0 *1 106.455,158.34
X$26420 368 630 369 644 645 cell_1rw
* cell instance $26421 r0 *1 106.455,158.34
X$26421 368 631 369 644 645 cell_1rw
* cell instance $26422 m0 *1 106.455,161.07
X$26422 368 632 369 644 645 cell_1rw
* cell instance $26423 r0 *1 106.455,161.07
X$26423 368 633 369 644 645 cell_1rw
* cell instance $26424 m0 *1 106.455,163.8
X$26424 368 634 369 644 645 cell_1rw
* cell instance $26425 r0 *1 106.455,163.8
X$26425 368 635 369 644 645 cell_1rw
* cell instance $26426 m0 *1 106.455,166.53
X$26426 368 637 369 644 645 cell_1rw
* cell instance $26427 r0 *1 106.455,166.53
X$26427 368 636 369 644 645 cell_1rw
* cell instance $26428 m0 *1 106.455,169.26
X$26428 368 639 369 644 645 cell_1rw
* cell instance $26429 r0 *1 106.455,169.26
X$26429 368 638 369 644 645 cell_1rw
* cell instance $26430 m0 *1 106.455,171.99
X$26430 368 640 369 644 645 cell_1rw
* cell instance $26431 r0 *1 106.455,171.99
X$26431 368 641 369 644 645 cell_1rw
* cell instance $26432 m0 *1 106.455,174.72
X$26432 368 642 369 644 645 cell_1rw
* cell instance $26433 r0 *1 106.455,174.72
X$26433 368 643 369 644 645 cell_1rw
* cell instance $26434 m0 *1 107.16,90.09
X$26434 370 581 371 644 645 cell_1rw
* cell instance $26435 r0 *1 107.16,90.09
X$26435 370 580 371 644 645 cell_1rw
* cell instance $26436 m0 *1 107.16,92.82
X$26436 370 583 371 644 645 cell_1rw
* cell instance $26437 r0 *1 107.16,92.82
X$26437 370 582 371 644 645 cell_1rw
* cell instance $26438 m0 *1 107.16,95.55
X$26438 370 584 371 644 645 cell_1rw
* cell instance $26439 r0 *1 107.16,95.55
X$26439 370 585 371 644 645 cell_1rw
* cell instance $26440 m0 *1 107.16,98.28
X$26440 370 586 371 644 645 cell_1rw
* cell instance $26441 m0 *1 107.16,101.01
X$26441 370 588 371 644 645 cell_1rw
* cell instance $26442 r0 *1 107.16,98.28
X$26442 370 587 371 644 645 cell_1rw
* cell instance $26443 r0 *1 107.16,101.01
X$26443 370 589 371 644 645 cell_1rw
* cell instance $26444 m0 *1 107.16,103.74
X$26444 370 590 371 644 645 cell_1rw
* cell instance $26445 r0 *1 107.16,103.74
X$26445 370 591 371 644 645 cell_1rw
* cell instance $26446 m0 *1 107.16,106.47
X$26446 370 593 371 644 645 cell_1rw
* cell instance $26447 m0 *1 107.16,109.2
X$26447 370 594 371 644 645 cell_1rw
* cell instance $26448 r0 *1 107.16,106.47
X$26448 370 592 371 644 645 cell_1rw
* cell instance $26449 r0 *1 107.16,109.2
X$26449 370 595 371 644 645 cell_1rw
* cell instance $26450 m0 *1 107.16,111.93
X$26450 370 597 371 644 645 cell_1rw
* cell instance $26451 r0 *1 107.16,111.93
X$26451 370 596 371 644 645 cell_1rw
* cell instance $26452 m0 *1 107.16,114.66
X$26452 370 598 371 644 645 cell_1rw
* cell instance $26453 m0 *1 107.16,117.39
X$26453 370 600 371 644 645 cell_1rw
* cell instance $26454 r0 *1 107.16,114.66
X$26454 370 599 371 644 645 cell_1rw
* cell instance $26455 r0 *1 107.16,117.39
X$26455 370 601 371 644 645 cell_1rw
* cell instance $26456 m0 *1 107.16,120.12
X$26456 370 602 371 644 645 cell_1rw
* cell instance $26457 r0 *1 107.16,120.12
X$26457 370 603 371 644 645 cell_1rw
* cell instance $26458 m0 *1 107.16,122.85
X$26458 370 604 371 644 645 cell_1rw
* cell instance $26459 r0 *1 107.16,122.85
X$26459 370 605 371 644 645 cell_1rw
* cell instance $26460 m0 *1 107.16,125.58
X$26460 370 606 371 644 645 cell_1rw
* cell instance $26461 r0 *1 107.16,125.58
X$26461 370 607 371 644 645 cell_1rw
* cell instance $26462 m0 *1 107.16,128.31
X$26462 370 609 371 644 645 cell_1rw
* cell instance $26463 r0 *1 107.16,128.31
X$26463 370 608 371 644 645 cell_1rw
* cell instance $26464 m0 *1 107.16,131.04
X$26464 370 610 371 644 645 cell_1rw
* cell instance $26465 r0 *1 107.16,131.04
X$26465 370 611 371 644 645 cell_1rw
* cell instance $26466 m0 *1 107.16,133.77
X$26466 370 612 371 644 645 cell_1rw
* cell instance $26467 r0 *1 107.16,133.77
X$26467 370 613 371 644 645 cell_1rw
* cell instance $26468 m0 *1 107.16,136.5
X$26468 370 615 371 644 645 cell_1rw
* cell instance $26469 r0 *1 107.16,136.5
X$26469 370 614 371 644 645 cell_1rw
* cell instance $26470 m0 *1 107.16,139.23
X$26470 370 617 371 644 645 cell_1rw
* cell instance $26471 r0 *1 107.16,139.23
X$26471 370 616 371 644 645 cell_1rw
* cell instance $26472 m0 *1 107.16,141.96
X$26472 370 618 371 644 645 cell_1rw
* cell instance $26473 r0 *1 107.16,141.96
X$26473 370 619 371 644 645 cell_1rw
* cell instance $26474 m0 *1 107.16,144.69
X$26474 370 620 371 644 645 cell_1rw
* cell instance $26475 r0 *1 107.16,144.69
X$26475 370 621 371 644 645 cell_1rw
* cell instance $26476 m0 *1 107.16,147.42
X$26476 370 622 371 644 645 cell_1rw
* cell instance $26477 r0 *1 107.16,147.42
X$26477 370 623 371 644 645 cell_1rw
* cell instance $26478 m0 *1 107.16,150.15
X$26478 370 624 371 644 645 cell_1rw
* cell instance $26479 r0 *1 107.16,150.15
X$26479 370 625 371 644 645 cell_1rw
* cell instance $26480 m0 *1 107.16,152.88
X$26480 370 626 371 644 645 cell_1rw
* cell instance $26481 r0 *1 107.16,152.88
X$26481 370 627 371 644 645 cell_1rw
* cell instance $26482 m0 *1 107.16,155.61
X$26482 370 628 371 644 645 cell_1rw
* cell instance $26483 r0 *1 107.16,155.61
X$26483 370 629 371 644 645 cell_1rw
* cell instance $26484 m0 *1 107.16,158.34
X$26484 370 630 371 644 645 cell_1rw
* cell instance $26485 r0 *1 107.16,158.34
X$26485 370 631 371 644 645 cell_1rw
* cell instance $26486 m0 *1 107.16,161.07
X$26486 370 632 371 644 645 cell_1rw
* cell instance $26487 r0 *1 107.16,161.07
X$26487 370 633 371 644 645 cell_1rw
* cell instance $26488 m0 *1 107.16,163.8
X$26488 370 634 371 644 645 cell_1rw
* cell instance $26489 r0 *1 107.16,163.8
X$26489 370 635 371 644 645 cell_1rw
* cell instance $26490 m0 *1 107.16,166.53
X$26490 370 637 371 644 645 cell_1rw
* cell instance $26491 r0 *1 107.16,166.53
X$26491 370 636 371 644 645 cell_1rw
* cell instance $26492 m0 *1 107.16,169.26
X$26492 370 639 371 644 645 cell_1rw
* cell instance $26493 r0 *1 107.16,169.26
X$26493 370 638 371 644 645 cell_1rw
* cell instance $26494 m0 *1 107.16,171.99
X$26494 370 640 371 644 645 cell_1rw
* cell instance $26495 r0 *1 107.16,171.99
X$26495 370 641 371 644 645 cell_1rw
* cell instance $26496 m0 *1 107.16,174.72
X$26496 370 642 371 644 645 cell_1rw
* cell instance $26497 r0 *1 107.16,174.72
X$26497 370 643 371 644 645 cell_1rw
* cell instance $26498 m0 *1 107.865,90.09
X$26498 372 581 373 644 645 cell_1rw
* cell instance $26499 r0 *1 107.865,90.09
X$26499 372 580 373 644 645 cell_1rw
* cell instance $26500 m0 *1 107.865,92.82
X$26500 372 583 373 644 645 cell_1rw
* cell instance $26501 r0 *1 107.865,92.82
X$26501 372 582 373 644 645 cell_1rw
* cell instance $26502 m0 *1 107.865,95.55
X$26502 372 584 373 644 645 cell_1rw
* cell instance $26503 r0 *1 107.865,95.55
X$26503 372 585 373 644 645 cell_1rw
* cell instance $26504 m0 *1 107.865,98.28
X$26504 372 586 373 644 645 cell_1rw
* cell instance $26505 r0 *1 107.865,98.28
X$26505 372 587 373 644 645 cell_1rw
* cell instance $26506 m0 *1 107.865,101.01
X$26506 372 588 373 644 645 cell_1rw
* cell instance $26507 r0 *1 107.865,101.01
X$26507 372 589 373 644 645 cell_1rw
* cell instance $26508 m0 *1 107.865,103.74
X$26508 372 590 373 644 645 cell_1rw
* cell instance $26509 r0 *1 107.865,103.74
X$26509 372 591 373 644 645 cell_1rw
* cell instance $26510 m0 *1 107.865,106.47
X$26510 372 593 373 644 645 cell_1rw
* cell instance $26511 m0 *1 107.865,109.2
X$26511 372 594 373 644 645 cell_1rw
* cell instance $26512 r0 *1 107.865,106.47
X$26512 372 592 373 644 645 cell_1rw
* cell instance $26513 m0 *1 107.865,111.93
X$26513 372 597 373 644 645 cell_1rw
* cell instance $26514 r0 *1 107.865,109.2
X$26514 372 595 373 644 645 cell_1rw
* cell instance $26515 r0 *1 107.865,111.93
X$26515 372 596 373 644 645 cell_1rw
* cell instance $26516 m0 *1 107.865,114.66
X$26516 372 598 373 644 645 cell_1rw
* cell instance $26517 m0 *1 107.865,117.39
X$26517 372 600 373 644 645 cell_1rw
* cell instance $26518 r0 *1 107.865,114.66
X$26518 372 599 373 644 645 cell_1rw
* cell instance $26519 r0 *1 107.865,117.39
X$26519 372 601 373 644 645 cell_1rw
* cell instance $26520 m0 *1 107.865,120.12
X$26520 372 602 373 644 645 cell_1rw
* cell instance $26521 r0 *1 107.865,120.12
X$26521 372 603 373 644 645 cell_1rw
* cell instance $26522 m0 *1 107.865,122.85
X$26522 372 604 373 644 645 cell_1rw
* cell instance $26523 r0 *1 107.865,122.85
X$26523 372 605 373 644 645 cell_1rw
* cell instance $26524 m0 *1 107.865,125.58
X$26524 372 606 373 644 645 cell_1rw
* cell instance $26525 r0 *1 107.865,125.58
X$26525 372 607 373 644 645 cell_1rw
* cell instance $26526 m0 *1 107.865,128.31
X$26526 372 609 373 644 645 cell_1rw
* cell instance $26527 r0 *1 107.865,128.31
X$26527 372 608 373 644 645 cell_1rw
* cell instance $26528 m0 *1 107.865,131.04
X$26528 372 610 373 644 645 cell_1rw
* cell instance $26529 r0 *1 107.865,131.04
X$26529 372 611 373 644 645 cell_1rw
* cell instance $26530 m0 *1 107.865,133.77
X$26530 372 612 373 644 645 cell_1rw
* cell instance $26531 m0 *1 107.865,136.5
X$26531 372 615 373 644 645 cell_1rw
* cell instance $26532 r0 *1 107.865,133.77
X$26532 372 613 373 644 645 cell_1rw
* cell instance $26533 r0 *1 107.865,136.5
X$26533 372 614 373 644 645 cell_1rw
* cell instance $26534 m0 *1 107.865,139.23
X$26534 372 617 373 644 645 cell_1rw
* cell instance $26535 r0 *1 107.865,139.23
X$26535 372 616 373 644 645 cell_1rw
* cell instance $26536 m0 *1 107.865,141.96
X$26536 372 618 373 644 645 cell_1rw
* cell instance $26537 r0 *1 107.865,141.96
X$26537 372 619 373 644 645 cell_1rw
* cell instance $26538 m0 *1 107.865,144.69
X$26538 372 620 373 644 645 cell_1rw
* cell instance $26539 r0 *1 107.865,144.69
X$26539 372 621 373 644 645 cell_1rw
* cell instance $26540 m0 *1 107.865,147.42
X$26540 372 622 373 644 645 cell_1rw
* cell instance $26541 r0 *1 107.865,147.42
X$26541 372 623 373 644 645 cell_1rw
* cell instance $26542 m0 *1 107.865,150.15
X$26542 372 624 373 644 645 cell_1rw
* cell instance $26543 r0 *1 107.865,150.15
X$26543 372 625 373 644 645 cell_1rw
* cell instance $26544 m0 *1 107.865,152.88
X$26544 372 626 373 644 645 cell_1rw
* cell instance $26545 m0 *1 107.865,155.61
X$26545 372 628 373 644 645 cell_1rw
* cell instance $26546 r0 *1 107.865,152.88
X$26546 372 627 373 644 645 cell_1rw
* cell instance $26547 r0 *1 107.865,155.61
X$26547 372 629 373 644 645 cell_1rw
* cell instance $26548 m0 *1 107.865,158.34
X$26548 372 630 373 644 645 cell_1rw
* cell instance $26549 r0 *1 107.865,158.34
X$26549 372 631 373 644 645 cell_1rw
* cell instance $26550 m0 *1 107.865,161.07
X$26550 372 632 373 644 645 cell_1rw
* cell instance $26551 r0 *1 107.865,161.07
X$26551 372 633 373 644 645 cell_1rw
* cell instance $26552 m0 *1 107.865,163.8
X$26552 372 634 373 644 645 cell_1rw
* cell instance $26553 r0 *1 107.865,163.8
X$26553 372 635 373 644 645 cell_1rw
* cell instance $26554 m0 *1 107.865,166.53
X$26554 372 637 373 644 645 cell_1rw
* cell instance $26555 m0 *1 107.865,169.26
X$26555 372 639 373 644 645 cell_1rw
* cell instance $26556 r0 *1 107.865,166.53
X$26556 372 636 373 644 645 cell_1rw
* cell instance $26557 r0 *1 107.865,169.26
X$26557 372 638 373 644 645 cell_1rw
* cell instance $26558 m0 *1 107.865,171.99
X$26558 372 640 373 644 645 cell_1rw
* cell instance $26559 m0 *1 107.865,174.72
X$26559 372 642 373 644 645 cell_1rw
* cell instance $26560 r0 *1 107.865,171.99
X$26560 372 641 373 644 645 cell_1rw
* cell instance $26561 r0 *1 107.865,174.72
X$26561 372 643 373 644 645 cell_1rw
* cell instance $26562 m0 *1 108.57,90.09
X$26562 374 581 375 644 645 cell_1rw
* cell instance $26563 r0 *1 108.57,90.09
X$26563 374 580 375 644 645 cell_1rw
* cell instance $26564 m0 *1 108.57,92.82
X$26564 374 583 375 644 645 cell_1rw
* cell instance $26565 r0 *1 108.57,92.82
X$26565 374 582 375 644 645 cell_1rw
* cell instance $26566 m0 *1 108.57,95.55
X$26566 374 584 375 644 645 cell_1rw
* cell instance $26567 m0 *1 108.57,98.28
X$26567 374 586 375 644 645 cell_1rw
* cell instance $26568 r0 *1 108.57,95.55
X$26568 374 585 375 644 645 cell_1rw
* cell instance $26569 r0 *1 108.57,98.28
X$26569 374 587 375 644 645 cell_1rw
* cell instance $26570 m0 *1 108.57,101.01
X$26570 374 588 375 644 645 cell_1rw
* cell instance $26571 r0 *1 108.57,101.01
X$26571 374 589 375 644 645 cell_1rw
* cell instance $26572 m0 *1 108.57,103.74
X$26572 374 590 375 644 645 cell_1rw
* cell instance $26573 r0 *1 108.57,103.74
X$26573 374 591 375 644 645 cell_1rw
* cell instance $26574 m0 *1 108.57,106.47
X$26574 374 593 375 644 645 cell_1rw
* cell instance $26575 r0 *1 108.57,106.47
X$26575 374 592 375 644 645 cell_1rw
* cell instance $26576 m0 *1 108.57,109.2
X$26576 374 594 375 644 645 cell_1rw
* cell instance $26577 r0 *1 108.57,109.2
X$26577 374 595 375 644 645 cell_1rw
* cell instance $26578 m0 *1 108.57,111.93
X$26578 374 597 375 644 645 cell_1rw
* cell instance $26579 r0 *1 108.57,111.93
X$26579 374 596 375 644 645 cell_1rw
* cell instance $26580 m0 *1 108.57,114.66
X$26580 374 598 375 644 645 cell_1rw
* cell instance $26581 r0 *1 108.57,114.66
X$26581 374 599 375 644 645 cell_1rw
* cell instance $26582 m0 *1 108.57,117.39
X$26582 374 600 375 644 645 cell_1rw
* cell instance $26583 r0 *1 108.57,117.39
X$26583 374 601 375 644 645 cell_1rw
* cell instance $26584 m0 *1 108.57,120.12
X$26584 374 602 375 644 645 cell_1rw
* cell instance $26585 r0 *1 108.57,120.12
X$26585 374 603 375 644 645 cell_1rw
* cell instance $26586 m0 *1 108.57,122.85
X$26586 374 604 375 644 645 cell_1rw
* cell instance $26587 r0 *1 108.57,122.85
X$26587 374 605 375 644 645 cell_1rw
* cell instance $26588 m0 *1 108.57,125.58
X$26588 374 606 375 644 645 cell_1rw
* cell instance $26589 r0 *1 108.57,125.58
X$26589 374 607 375 644 645 cell_1rw
* cell instance $26590 m0 *1 108.57,128.31
X$26590 374 609 375 644 645 cell_1rw
* cell instance $26591 r0 *1 108.57,128.31
X$26591 374 608 375 644 645 cell_1rw
* cell instance $26592 m0 *1 108.57,131.04
X$26592 374 610 375 644 645 cell_1rw
* cell instance $26593 m0 *1 108.57,133.77
X$26593 374 612 375 644 645 cell_1rw
* cell instance $26594 r0 *1 108.57,131.04
X$26594 374 611 375 644 645 cell_1rw
* cell instance $26595 r0 *1 108.57,133.77
X$26595 374 613 375 644 645 cell_1rw
* cell instance $26596 m0 *1 108.57,136.5
X$26596 374 615 375 644 645 cell_1rw
* cell instance $26597 r0 *1 108.57,136.5
X$26597 374 614 375 644 645 cell_1rw
* cell instance $26598 m0 *1 108.57,139.23
X$26598 374 617 375 644 645 cell_1rw
* cell instance $26599 r0 *1 108.57,139.23
X$26599 374 616 375 644 645 cell_1rw
* cell instance $26600 m0 *1 108.57,141.96
X$26600 374 618 375 644 645 cell_1rw
* cell instance $26601 r0 *1 108.57,141.96
X$26601 374 619 375 644 645 cell_1rw
* cell instance $26602 m0 *1 108.57,144.69
X$26602 374 620 375 644 645 cell_1rw
* cell instance $26603 r0 *1 108.57,144.69
X$26603 374 621 375 644 645 cell_1rw
* cell instance $26604 m0 *1 108.57,147.42
X$26604 374 622 375 644 645 cell_1rw
* cell instance $26605 r0 *1 108.57,147.42
X$26605 374 623 375 644 645 cell_1rw
* cell instance $26606 m0 *1 108.57,150.15
X$26606 374 624 375 644 645 cell_1rw
* cell instance $26607 r0 *1 108.57,150.15
X$26607 374 625 375 644 645 cell_1rw
* cell instance $26608 m0 *1 108.57,152.88
X$26608 374 626 375 644 645 cell_1rw
* cell instance $26609 r0 *1 108.57,152.88
X$26609 374 627 375 644 645 cell_1rw
* cell instance $26610 m0 *1 108.57,155.61
X$26610 374 628 375 644 645 cell_1rw
* cell instance $26611 r0 *1 108.57,155.61
X$26611 374 629 375 644 645 cell_1rw
* cell instance $26612 m0 *1 108.57,158.34
X$26612 374 630 375 644 645 cell_1rw
* cell instance $26613 r0 *1 108.57,158.34
X$26613 374 631 375 644 645 cell_1rw
* cell instance $26614 m0 *1 108.57,161.07
X$26614 374 632 375 644 645 cell_1rw
* cell instance $26615 r0 *1 108.57,161.07
X$26615 374 633 375 644 645 cell_1rw
* cell instance $26616 m0 *1 108.57,163.8
X$26616 374 634 375 644 645 cell_1rw
* cell instance $26617 r0 *1 108.57,163.8
X$26617 374 635 375 644 645 cell_1rw
* cell instance $26618 m0 *1 108.57,166.53
X$26618 374 637 375 644 645 cell_1rw
* cell instance $26619 r0 *1 108.57,166.53
X$26619 374 636 375 644 645 cell_1rw
* cell instance $26620 m0 *1 108.57,169.26
X$26620 374 639 375 644 645 cell_1rw
* cell instance $26621 r0 *1 108.57,169.26
X$26621 374 638 375 644 645 cell_1rw
* cell instance $26622 m0 *1 108.57,171.99
X$26622 374 640 375 644 645 cell_1rw
* cell instance $26623 m0 *1 108.57,174.72
X$26623 374 642 375 644 645 cell_1rw
* cell instance $26624 r0 *1 108.57,171.99
X$26624 374 641 375 644 645 cell_1rw
* cell instance $26625 r0 *1 108.57,174.72
X$26625 374 643 375 644 645 cell_1rw
* cell instance $26626 m0 *1 109.275,90.09
X$26626 376 581 377 644 645 cell_1rw
* cell instance $26627 r0 *1 109.275,90.09
X$26627 376 580 377 644 645 cell_1rw
* cell instance $26628 m0 *1 109.275,92.82
X$26628 376 583 377 644 645 cell_1rw
* cell instance $26629 r0 *1 109.275,92.82
X$26629 376 582 377 644 645 cell_1rw
* cell instance $26630 m0 *1 109.275,95.55
X$26630 376 584 377 644 645 cell_1rw
* cell instance $26631 r0 *1 109.275,95.55
X$26631 376 585 377 644 645 cell_1rw
* cell instance $26632 m0 *1 109.275,98.28
X$26632 376 586 377 644 645 cell_1rw
* cell instance $26633 r0 *1 109.275,98.28
X$26633 376 587 377 644 645 cell_1rw
* cell instance $26634 m0 *1 109.275,101.01
X$26634 376 588 377 644 645 cell_1rw
* cell instance $26635 r0 *1 109.275,101.01
X$26635 376 589 377 644 645 cell_1rw
* cell instance $26636 m0 *1 109.275,103.74
X$26636 376 590 377 644 645 cell_1rw
* cell instance $26637 r0 *1 109.275,103.74
X$26637 376 591 377 644 645 cell_1rw
* cell instance $26638 m0 *1 109.275,106.47
X$26638 376 593 377 644 645 cell_1rw
* cell instance $26639 r0 *1 109.275,106.47
X$26639 376 592 377 644 645 cell_1rw
* cell instance $26640 m0 *1 109.275,109.2
X$26640 376 594 377 644 645 cell_1rw
* cell instance $26641 r0 *1 109.275,109.2
X$26641 376 595 377 644 645 cell_1rw
* cell instance $26642 m0 *1 109.275,111.93
X$26642 376 597 377 644 645 cell_1rw
* cell instance $26643 r0 *1 109.275,111.93
X$26643 376 596 377 644 645 cell_1rw
* cell instance $26644 m0 *1 109.275,114.66
X$26644 376 598 377 644 645 cell_1rw
* cell instance $26645 r0 *1 109.275,114.66
X$26645 376 599 377 644 645 cell_1rw
* cell instance $26646 m0 *1 109.275,117.39
X$26646 376 600 377 644 645 cell_1rw
* cell instance $26647 r0 *1 109.275,117.39
X$26647 376 601 377 644 645 cell_1rw
* cell instance $26648 m0 *1 109.275,120.12
X$26648 376 602 377 644 645 cell_1rw
* cell instance $26649 r0 *1 109.275,120.12
X$26649 376 603 377 644 645 cell_1rw
* cell instance $26650 m0 *1 109.275,122.85
X$26650 376 604 377 644 645 cell_1rw
* cell instance $26651 r0 *1 109.275,122.85
X$26651 376 605 377 644 645 cell_1rw
* cell instance $26652 m0 *1 109.275,125.58
X$26652 376 606 377 644 645 cell_1rw
* cell instance $26653 r0 *1 109.275,125.58
X$26653 376 607 377 644 645 cell_1rw
* cell instance $26654 m0 *1 109.275,128.31
X$26654 376 609 377 644 645 cell_1rw
* cell instance $26655 r0 *1 109.275,128.31
X$26655 376 608 377 644 645 cell_1rw
* cell instance $26656 m0 *1 109.275,131.04
X$26656 376 610 377 644 645 cell_1rw
* cell instance $26657 r0 *1 109.275,131.04
X$26657 376 611 377 644 645 cell_1rw
* cell instance $26658 m0 *1 109.275,133.77
X$26658 376 612 377 644 645 cell_1rw
* cell instance $26659 r0 *1 109.275,133.77
X$26659 376 613 377 644 645 cell_1rw
* cell instance $26660 m0 *1 109.275,136.5
X$26660 376 615 377 644 645 cell_1rw
* cell instance $26661 r0 *1 109.275,136.5
X$26661 376 614 377 644 645 cell_1rw
* cell instance $26662 m0 *1 109.275,139.23
X$26662 376 617 377 644 645 cell_1rw
* cell instance $26663 r0 *1 109.275,139.23
X$26663 376 616 377 644 645 cell_1rw
* cell instance $26664 m0 *1 109.275,141.96
X$26664 376 618 377 644 645 cell_1rw
* cell instance $26665 r0 *1 109.275,141.96
X$26665 376 619 377 644 645 cell_1rw
* cell instance $26666 m0 *1 109.275,144.69
X$26666 376 620 377 644 645 cell_1rw
* cell instance $26667 r0 *1 109.275,144.69
X$26667 376 621 377 644 645 cell_1rw
* cell instance $26668 m0 *1 109.275,147.42
X$26668 376 622 377 644 645 cell_1rw
* cell instance $26669 r0 *1 109.275,147.42
X$26669 376 623 377 644 645 cell_1rw
* cell instance $26670 m0 *1 109.275,150.15
X$26670 376 624 377 644 645 cell_1rw
* cell instance $26671 r0 *1 109.275,150.15
X$26671 376 625 377 644 645 cell_1rw
* cell instance $26672 m0 *1 109.275,152.88
X$26672 376 626 377 644 645 cell_1rw
* cell instance $26673 r0 *1 109.275,152.88
X$26673 376 627 377 644 645 cell_1rw
* cell instance $26674 m0 *1 109.275,155.61
X$26674 376 628 377 644 645 cell_1rw
* cell instance $26675 r0 *1 109.275,155.61
X$26675 376 629 377 644 645 cell_1rw
* cell instance $26676 m0 *1 109.275,158.34
X$26676 376 630 377 644 645 cell_1rw
* cell instance $26677 m0 *1 109.275,161.07
X$26677 376 632 377 644 645 cell_1rw
* cell instance $26678 r0 *1 109.275,158.34
X$26678 376 631 377 644 645 cell_1rw
* cell instance $26679 r0 *1 109.275,161.07
X$26679 376 633 377 644 645 cell_1rw
* cell instance $26680 m0 *1 109.275,163.8
X$26680 376 634 377 644 645 cell_1rw
* cell instance $26681 r0 *1 109.275,163.8
X$26681 376 635 377 644 645 cell_1rw
* cell instance $26682 m0 *1 109.275,166.53
X$26682 376 637 377 644 645 cell_1rw
* cell instance $26683 r0 *1 109.275,166.53
X$26683 376 636 377 644 645 cell_1rw
* cell instance $26684 m0 *1 109.275,169.26
X$26684 376 639 377 644 645 cell_1rw
* cell instance $26685 r0 *1 109.275,169.26
X$26685 376 638 377 644 645 cell_1rw
* cell instance $26686 m0 *1 109.275,171.99
X$26686 376 640 377 644 645 cell_1rw
* cell instance $26687 r0 *1 109.275,171.99
X$26687 376 641 377 644 645 cell_1rw
* cell instance $26688 m0 *1 109.275,174.72
X$26688 376 642 377 644 645 cell_1rw
* cell instance $26689 r0 *1 109.275,174.72
X$26689 376 643 377 644 645 cell_1rw
* cell instance $26690 m0 *1 109.98,90.09
X$26690 378 581 379 644 645 cell_1rw
* cell instance $26691 r0 *1 109.98,90.09
X$26691 378 580 379 644 645 cell_1rw
* cell instance $26692 m0 *1 109.98,92.82
X$26692 378 583 379 644 645 cell_1rw
* cell instance $26693 m0 *1 109.98,95.55
X$26693 378 584 379 644 645 cell_1rw
* cell instance $26694 r0 *1 109.98,92.82
X$26694 378 582 379 644 645 cell_1rw
* cell instance $26695 m0 *1 109.98,98.28
X$26695 378 586 379 644 645 cell_1rw
* cell instance $26696 r0 *1 109.98,95.55
X$26696 378 585 379 644 645 cell_1rw
* cell instance $26697 m0 *1 109.98,101.01
X$26697 378 588 379 644 645 cell_1rw
* cell instance $26698 r0 *1 109.98,98.28
X$26698 378 587 379 644 645 cell_1rw
* cell instance $26699 r0 *1 109.98,101.01
X$26699 378 589 379 644 645 cell_1rw
* cell instance $26700 m0 *1 109.98,103.74
X$26700 378 590 379 644 645 cell_1rw
* cell instance $26701 r0 *1 109.98,103.74
X$26701 378 591 379 644 645 cell_1rw
* cell instance $26702 m0 *1 109.98,106.47
X$26702 378 593 379 644 645 cell_1rw
* cell instance $26703 r0 *1 109.98,106.47
X$26703 378 592 379 644 645 cell_1rw
* cell instance $26704 m0 *1 109.98,109.2
X$26704 378 594 379 644 645 cell_1rw
* cell instance $26705 r0 *1 109.98,109.2
X$26705 378 595 379 644 645 cell_1rw
* cell instance $26706 m0 *1 109.98,111.93
X$26706 378 597 379 644 645 cell_1rw
* cell instance $26707 r0 *1 109.98,111.93
X$26707 378 596 379 644 645 cell_1rw
* cell instance $26708 m0 *1 109.98,114.66
X$26708 378 598 379 644 645 cell_1rw
* cell instance $26709 r0 *1 109.98,114.66
X$26709 378 599 379 644 645 cell_1rw
* cell instance $26710 m0 *1 109.98,117.39
X$26710 378 600 379 644 645 cell_1rw
* cell instance $26711 r0 *1 109.98,117.39
X$26711 378 601 379 644 645 cell_1rw
* cell instance $26712 m0 *1 109.98,120.12
X$26712 378 602 379 644 645 cell_1rw
* cell instance $26713 r0 *1 109.98,120.12
X$26713 378 603 379 644 645 cell_1rw
* cell instance $26714 m0 *1 109.98,122.85
X$26714 378 604 379 644 645 cell_1rw
* cell instance $26715 r0 *1 109.98,122.85
X$26715 378 605 379 644 645 cell_1rw
* cell instance $26716 m0 *1 109.98,125.58
X$26716 378 606 379 644 645 cell_1rw
* cell instance $26717 r0 *1 109.98,125.58
X$26717 378 607 379 644 645 cell_1rw
* cell instance $26718 m0 *1 109.98,128.31
X$26718 378 609 379 644 645 cell_1rw
* cell instance $26719 r0 *1 109.98,128.31
X$26719 378 608 379 644 645 cell_1rw
* cell instance $26720 m0 *1 109.98,131.04
X$26720 378 610 379 644 645 cell_1rw
* cell instance $26721 r0 *1 109.98,131.04
X$26721 378 611 379 644 645 cell_1rw
* cell instance $26722 m0 *1 109.98,133.77
X$26722 378 612 379 644 645 cell_1rw
* cell instance $26723 r0 *1 109.98,133.77
X$26723 378 613 379 644 645 cell_1rw
* cell instance $26724 m0 *1 109.98,136.5
X$26724 378 615 379 644 645 cell_1rw
* cell instance $26725 r0 *1 109.98,136.5
X$26725 378 614 379 644 645 cell_1rw
* cell instance $26726 m0 *1 109.98,139.23
X$26726 378 617 379 644 645 cell_1rw
* cell instance $26727 r0 *1 109.98,139.23
X$26727 378 616 379 644 645 cell_1rw
* cell instance $26728 m0 *1 109.98,141.96
X$26728 378 618 379 644 645 cell_1rw
* cell instance $26729 m0 *1 109.98,144.69
X$26729 378 620 379 644 645 cell_1rw
* cell instance $26730 r0 *1 109.98,141.96
X$26730 378 619 379 644 645 cell_1rw
* cell instance $26731 m0 *1 109.98,147.42
X$26731 378 622 379 644 645 cell_1rw
* cell instance $26732 r0 *1 109.98,144.69
X$26732 378 621 379 644 645 cell_1rw
* cell instance $26733 r0 *1 109.98,147.42
X$26733 378 623 379 644 645 cell_1rw
* cell instance $26734 m0 *1 109.98,150.15
X$26734 378 624 379 644 645 cell_1rw
* cell instance $26735 r0 *1 109.98,150.15
X$26735 378 625 379 644 645 cell_1rw
* cell instance $26736 m0 *1 109.98,152.88
X$26736 378 626 379 644 645 cell_1rw
* cell instance $26737 r0 *1 109.98,152.88
X$26737 378 627 379 644 645 cell_1rw
* cell instance $26738 m0 *1 109.98,155.61
X$26738 378 628 379 644 645 cell_1rw
* cell instance $26739 r0 *1 109.98,155.61
X$26739 378 629 379 644 645 cell_1rw
* cell instance $26740 m0 *1 109.98,158.34
X$26740 378 630 379 644 645 cell_1rw
* cell instance $26741 r0 *1 109.98,158.34
X$26741 378 631 379 644 645 cell_1rw
* cell instance $26742 m0 *1 109.98,161.07
X$26742 378 632 379 644 645 cell_1rw
* cell instance $26743 m0 *1 109.98,163.8
X$26743 378 634 379 644 645 cell_1rw
* cell instance $26744 r0 *1 109.98,161.07
X$26744 378 633 379 644 645 cell_1rw
* cell instance $26745 r0 *1 109.98,163.8
X$26745 378 635 379 644 645 cell_1rw
* cell instance $26746 m0 *1 109.98,166.53
X$26746 378 637 379 644 645 cell_1rw
* cell instance $26747 m0 *1 109.98,169.26
X$26747 378 639 379 644 645 cell_1rw
* cell instance $26748 r0 *1 109.98,166.53
X$26748 378 636 379 644 645 cell_1rw
* cell instance $26749 r0 *1 109.98,169.26
X$26749 378 638 379 644 645 cell_1rw
* cell instance $26750 m0 *1 109.98,171.99
X$26750 378 640 379 644 645 cell_1rw
* cell instance $26751 r0 *1 109.98,171.99
X$26751 378 641 379 644 645 cell_1rw
* cell instance $26752 m0 *1 109.98,174.72
X$26752 378 642 379 644 645 cell_1rw
* cell instance $26753 r0 *1 109.98,174.72
X$26753 378 643 379 644 645 cell_1rw
* cell instance $26754 m0 *1 110.685,90.09
X$26754 380 581 381 644 645 cell_1rw
* cell instance $26755 m0 *1 110.685,92.82
X$26755 380 583 381 644 645 cell_1rw
* cell instance $26756 r0 *1 110.685,90.09
X$26756 380 580 381 644 645 cell_1rw
* cell instance $26757 r0 *1 110.685,92.82
X$26757 380 582 381 644 645 cell_1rw
* cell instance $26758 m0 *1 110.685,95.55
X$26758 380 584 381 644 645 cell_1rw
* cell instance $26759 m0 *1 110.685,98.28
X$26759 380 586 381 644 645 cell_1rw
* cell instance $26760 r0 *1 110.685,95.55
X$26760 380 585 381 644 645 cell_1rw
* cell instance $26761 m0 *1 110.685,101.01
X$26761 380 588 381 644 645 cell_1rw
* cell instance $26762 r0 *1 110.685,98.28
X$26762 380 587 381 644 645 cell_1rw
* cell instance $26763 r0 *1 110.685,101.01
X$26763 380 589 381 644 645 cell_1rw
* cell instance $26764 m0 *1 110.685,103.74
X$26764 380 590 381 644 645 cell_1rw
* cell instance $26765 r0 *1 110.685,103.74
X$26765 380 591 381 644 645 cell_1rw
* cell instance $26766 m0 *1 110.685,106.47
X$26766 380 593 381 644 645 cell_1rw
* cell instance $26767 r0 *1 110.685,106.47
X$26767 380 592 381 644 645 cell_1rw
* cell instance $26768 m0 *1 110.685,109.2
X$26768 380 594 381 644 645 cell_1rw
* cell instance $26769 r0 *1 110.685,109.2
X$26769 380 595 381 644 645 cell_1rw
* cell instance $26770 m0 *1 110.685,111.93
X$26770 380 597 381 644 645 cell_1rw
* cell instance $26771 r0 *1 110.685,111.93
X$26771 380 596 381 644 645 cell_1rw
* cell instance $26772 m0 *1 110.685,114.66
X$26772 380 598 381 644 645 cell_1rw
* cell instance $26773 r0 *1 110.685,114.66
X$26773 380 599 381 644 645 cell_1rw
* cell instance $26774 m0 *1 110.685,117.39
X$26774 380 600 381 644 645 cell_1rw
* cell instance $26775 r0 *1 110.685,117.39
X$26775 380 601 381 644 645 cell_1rw
* cell instance $26776 m0 *1 110.685,120.12
X$26776 380 602 381 644 645 cell_1rw
* cell instance $26777 m0 *1 110.685,122.85
X$26777 380 604 381 644 645 cell_1rw
* cell instance $26778 r0 *1 110.685,120.12
X$26778 380 603 381 644 645 cell_1rw
* cell instance $26779 r0 *1 110.685,122.85
X$26779 380 605 381 644 645 cell_1rw
* cell instance $26780 m0 *1 110.685,125.58
X$26780 380 606 381 644 645 cell_1rw
* cell instance $26781 r0 *1 110.685,125.58
X$26781 380 607 381 644 645 cell_1rw
* cell instance $26782 m0 *1 110.685,128.31
X$26782 380 609 381 644 645 cell_1rw
* cell instance $26783 r0 *1 110.685,128.31
X$26783 380 608 381 644 645 cell_1rw
* cell instance $26784 m0 *1 110.685,131.04
X$26784 380 610 381 644 645 cell_1rw
* cell instance $26785 r0 *1 110.685,131.04
X$26785 380 611 381 644 645 cell_1rw
* cell instance $26786 m0 *1 110.685,133.77
X$26786 380 612 381 644 645 cell_1rw
* cell instance $26787 r0 *1 110.685,133.77
X$26787 380 613 381 644 645 cell_1rw
* cell instance $26788 m0 *1 110.685,136.5
X$26788 380 615 381 644 645 cell_1rw
* cell instance $26789 m0 *1 110.685,139.23
X$26789 380 617 381 644 645 cell_1rw
* cell instance $26790 r0 *1 110.685,136.5
X$26790 380 614 381 644 645 cell_1rw
* cell instance $26791 r0 *1 110.685,139.23
X$26791 380 616 381 644 645 cell_1rw
* cell instance $26792 m0 *1 110.685,141.96
X$26792 380 618 381 644 645 cell_1rw
* cell instance $26793 r0 *1 110.685,141.96
X$26793 380 619 381 644 645 cell_1rw
* cell instance $26794 m0 *1 110.685,144.69
X$26794 380 620 381 644 645 cell_1rw
* cell instance $26795 m0 *1 110.685,147.42
X$26795 380 622 381 644 645 cell_1rw
* cell instance $26796 r0 *1 110.685,144.69
X$26796 380 621 381 644 645 cell_1rw
* cell instance $26797 r0 *1 110.685,147.42
X$26797 380 623 381 644 645 cell_1rw
* cell instance $26798 m0 *1 110.685,150.15
X$26798 380 624 381 644 645 cell_1rw
* cell instance $26799 r0 *1 110.685,150.15
X$26799 380 625 381 644 645 cell_1rw
* cell instance $26800 m0 *1 110.685,152.88
X$26800 380 626 381 644 645 cell_1rw
* cell instance $26801 r0 *1 110.685,152.88
X$26801 380 627 381 644 645 cell_1rw
* cell instance $26802 m0 *1 110.685,155.61
X$26802 380 628 381 644 645 cell_1rw
* cell instance $26803 r0 *1 110.685,155.61
X$26803 380 629 381 644 645 cell_1rw
* cell instance $26804 m0 *1 110.685,158.34
X$26804 380 630 381 644 645 cell_1rw
* cell instance $26805 r0 *1 110.685,158.34
X$26805 380 631 381 644 645 cell_1rw
* cell instance $26806 m0 *1 110.685,161.07
X$26806 380 632 381 644 645 cell_1rw
* cell instance $26807 r0 *1 110.685,161.07
X$26807 380 633 381 644 645 cell_1rw
* cell instance $26808 m0 *1 110.685,163.8
X$26808 380 634 381 644 645 cell_1rw
* cell instance $26809 r0 *1 110.685,163.8
X$26809 380 635 381 644 645 cell_1rw
* cell instance $26810 m0 *1 110.685,166.53
X$26810 380 637 381 644 645 cell_1rw
* cell instance $26811 m0 *1 110.685,169.26
X$26811 380 639 381 644 645 cell_1rw
* cell instance $26812 r0 *1 110.685,166.53
X$26812 380 636 381 644 645 cell_1rw
* cell instance $26813 r0 *1 110.685,169.26
X$26813 380 638 381 644 645 cell_1rw
* cell instance $26814 m0 *1 110.685,171.99
X$26814 380 640 381 644 645 cell_1rw
* cell instance $26815 m0 *1 110.685,174.72
X$26815 380 642 381 644 645 cell_1rw
* cell instance $26816 r0 *1 110.685,171.99
X$26816 380 641 381 644 645 cell_1rw
* cell instance $26817 r0 *1 110.685,174.72
X$26817 380 643 381 644 645 cell_1rw
* cell instance $26818 m0 *1 111.39,90.09
X$26818 382 581 383 644 645 cell_1rw
* cell instance $26819 r0 *1 111.39,90.09
X$26819 382 580 383 644 645 cell_1rw
* cell instance $26820 m0 *1 111.39,92.82
X$26820 382 583 383 644 645 cell_1rw
* cell instance $26821 m0 *1 111.39,95.55
X$26821 382 584 383 644 645 cell_1rw
* cell instance $26822 r0 *1 111.39,92.82
X$26822 382 582 383 644 645 cell_1rw
* cell instance $26823 r0 *1 111.39,95.55
X$26823 382 585 383 644 645 cell_1rw
* cell instance $26824 m0 *1 111.39,98.28
X$26824 382 586 383 644 645 cell_1rw
* cell instance $26825 m0 *1 111.39,101.01
X$26825 382 588 383 644 645 cell_1rw
* cell instance $26826 r0 *1 111.39,98.28
X$26826 382 587 383 644 645 cell_1rw
* cell instance $26827 r0 *1 111.39,101.01
X$26827 382 589 383 644 645 cell_1rw
* cell instance $26828 m0 *1 111.39,103.74
X$26828 382 590 383 644 645 cell_1rw
* cell instance $26829 r0 *1 111.39,103.74
X$26829 382 591 383 644 645 cell_1rw
* cell instance $26830 m0 *1 111.39,106.47
X$26830 382 593 383 644 645 cell_1rw
* cell instance $26831 r0 *1 111.39,106.47
X$26831 382 592 383 644 645 cell_1rw
* cell instance $26832 m0 *1 111.39,109.2
X$26832 382 594 383 644 645 cell_1rw
* cell instance $26833 r0 *1 111.39,109.2
X$26833 382 595 383 644 645 cell_1rw
* cell instance $26834 m0 *1 111.39,111.93
X$26834 382 597 383 644 645 cell_1rw
* cell instance $26835 r0 *1 111.39,111.93
X$26835 382 596 383 644 645 cell_1rw
* cell instance $26836 m0 *1 111.39,114.66
X$26836 382 598 383 644 645 cell_1rw
* cell instance $26837 r0 *1 111.39,114.66
X$26837 382 599 383 644 645 cell_1rw
* cell instance $26838 m0 *1 111.39,117.39
X$26838 382 600 383 644 645 cell_1rw
* cell instance $26839 m0 *1 111.39,120.12
X$26839 382 602 383 644 645 cell_1rw
* cell instance $26840 r0 *1 111.39,117.39
X$26840 382 601 383 644 645 cell_1rw
* cell instance $26841 r0 *1 111.39,120.12
X$26841 382 603 383 644 645 cell_1rw
* cell instance $26842 m0 *1 111.39,122.85
X$26842 382 604 383 644 645 cell_1rw
* cell instance $26843 r0 *1 111.39,122.85
X$26843 382 605 383 644 645 cell_1rw
* cell instance $26844 m0 *1 111.39,125.58
X$26844 382 606 383 644 645 cell_1rw
* cell instance $26845 r0 *1 111.39,125.58
X$26845 382 607 383 644 645 cell_1rw
* cell instance $26846 m0 *1 111.39,128.31
X$26846 382 609 383 644 645 cell_1rw
* cell instance $26847 r0 *1 111.39,128.31
X$26847 382 608 383 644 645 cell_1rw
* cell instance $26848 m0 *1 111.39,131.04
X$26848 382 610 383 644 645 cell_1rw
* cell instance $26849 r0 *1 111.39,131.04
X$26849 382 611 383 644 645 cell_1rw
* cell instance $26850 m0 *1 111.39,133.77
X$26850 382 612 383 644 645 cell_1rw
* cell instance $26851 m0 *1 111.39,136.5
X$26851 382 615 383 644 645 cell_1rw
* cell instance $26852 r0 *1 111.39,133.77
X$26852 382 613 383 644 645 cell_1rw
* cell instance $26853 r0 *1 111.39,136.5
X$26853 382 614 383 644 645 cell_1rw
* cell instance $26854 m0 *1 111.39,139.23
X$26854 382 617 383 644 645 cell_1rw
* cell instance $26855 r0 *1 111.39,139.23
X$26855 382 616 383 644 645 cell_1rw
* cell instance $26856 m0 *1 111.39,141.96
X$26856 382 618 383 644 645 cell_1rw
* cell instance $26857 r0 *1 111.39,141.96
X$26857 382 619 383 644 645 cell_1rw
* cell instance $26858 m0 *1 111.39,144.69
X$26858 382 620 383 644 645 cell_1rw
* cell instance $26859 r0 *1 111.39,144.69
X$26859 382 621 383 644 645 cell_1rw
* cell instance $26860 m0 *1 111.39,147.42
X$26860 382 622 383 644 645 cell_1rw
* cell instance $26861 r0 *1 111.39,147.42
X$26861 382 623 383 644 645 cell_1rw
* cell instance $26862 m0 *1 111.39,150.15
X$26862 382 624 383 644 645 cell_1rw
* cell instance $26863 m0 *1 111.39,152.88
X$26863 382 626 383 644 645 cell_1rw
* cell instance $26864 r0 *1 111.39,150.15
X$26864 382 625 383 644 645 cell_1rw
* cell instance $26865 r0 *1 111.39,152.88
X$26865 382 627 383 644 645 cell_1rw
* cell instance $26866 m0 *1 111.39,155.61
X$26866 382 628 383 644 645 cell_1rw
* cell instance $26867 r0 *1 111.39,155.61
X$26867 382 629 383 644 645 cell_1rw
* cell instance $26868 m0 *1 111.39,158.34
X$26868 382 630 383 644 645 cell_1rw
* cell instance $26869 r0 *1 111.39,158.34
X$26869 382 631 383 644 645 cell_1rw
* cell instance $26870 m0 *1 111.39,161.07
X$26870 382 632 383 644 645 cell_1rw
* cell instance $26871 m0 *1 111.39,163.8
X$26871 382 634 383 644 645 cell_1rw
* cell instance $26872 r0 *1 111.39,161.07
X$26872 382 633 383 644 645 cell_1rw
* cell instance $26873 m0 *1 111.39,166.53
X$26873 382 637 383 644 645 cell_1rw
* cell instance $26874 r0 *1 111.39,163.8
X$26874 382 635 383 644 645 cell_1rw
* cell instance $26875 r0 *1 111.39,166.53
X$26875 382 636 383 644 645 cell_1rw
* cell instance $26876 m0 *1 111.39,169.26
X$26876 382 639 383 644 645 cell_1rw
* cell instance $26877 r0 *1 111.39,169.26
X$26877 382 638 383 644 645 cell_1rw
* cell instance $26878 m0 *1 111.39,171.99
X$26878 382 640 383 644 645 cell_1rw
* cell instance $26879 m0 *1 111.39,174.72
X$26879 382 642 383 644 645 cell_1rw
* cell instance $26880 r0 *1 111.39,171.99
X$26880 382 641 383 644 645 cell_1rw
* cell instance $26881 r0 *1 111.39,174.72
X$26881 382 643 383 644 645 cell_1rw
* cell instance $26882 m0 *1 112.095,90.09
X$26882 384 581 385 644 645 cell_1rw
* cell instance $26883 r0 *1 112.095,90.09
X$26883 384 580 385 644 645 cell_1rw
* cell instance $26884 m0 *1 112.095,92.82
X$26884 384 583 385 644 645 cell_1rw
* cell instance $26885 r0 *1 112.095,92.82
X$26885 384 582 385 644 645 cell_1rw
* cell instance $26886 m0 *1 112.095,95.55
X$26886 384 584 385 644 645 cell_1rw
* cell instance $26887 m0 *1 112.095,98.28
X$26887 384 586 385 644 645 cell_1rw
* cell instance $26888 r0 *1 112.095,95.55
X$26888 384 585 385 644 645 cell_1rw
* cell instance $26889 r0 *1 112.095,98.28
X$26889 384 587 385 644 645 cell_1rw
* cell instance $26890 m0 *1 112.095,101.01
X$26890 384 588 385 644 645 cell_1rw
* cell instance $26891 r0 *1 112.095,101.01
X$26891 384 589 385 644 645 cell_1rw
* cell instance $26892 m0 *1 112.095,103.74
X$26892 384 590 385 644 645 cell_1rw
* cell instance $26893 r0 *1 112.095,103.74
X$26893 384 591 385 644 645 cell_1rw
* cell instance $26894 m0 *1 112.095,106.47
X$26894 384 593 385 644 645 cell_1rw
* cell instance $26895 m0 *1 112.095,109.2
X$26895 384 594 385 644 645 cell_1rw
* cell instance $26896 r0 *1 112.095,106.47
X$26896 384 592 385 644 645 cell_1rw
* cell instance $26897 m0 *1 112.095,111.93
X$26897 384 597 385 644 645 cell_1rw
* cell instance $26898 r0 *1 112.095,109.2
X$26898 384 595 385 644 645 cell_1rw
* cell instance $26899 r0 *1 112.095,111.93
X$26899 384 596 385 644 645 cell_1rw
* cell instance $26900 m0 *1 112.095,114.66
X$26900 384 598 385 644 645 cell_1rw
* cell instance $26901 r0 *1 112.095,114.66
X$26901 384 599 385 644 645 cell_1rw
* cell instance $26902 m0 *1 112.095,117.39
X$26902 384 600 385 644 645 cell_1rw
* cell instance $26903 r0 *1 112.095,117.39
X$26903 384 601 385 644 645 cell_1rw
* cell instance $26904 m0 *1 112.095,120.12
X$26904 384 602 385 644 645 cell_1rw
* cell instance $26905 m0 *1 112.095,122.85
X$26905 384 604 385 644 645 cell_1rw
* cell instance $26906 r0 *1 112.095,120.12
X$26906 384 603 385 644 645 cell_1rw
* cell instance $26907 r0 *1 112.095,122.85
X$26907 384 605 385 644 645 cell_1rw
* cell instance $26908 m0 *1 112.095,125.58
X$26908 384 606 385 644 645 cell_1rw
* cell instance $26909 m0 *1 112.095,128.31
X$26909 384 609 385 644 645 cell_1rw
* cell instance $26910 r0 *1 112.095,125.58
X$26910 384 607 385 644 645 cell_1rw
* cell instance $26911 r0 *1 112.095,128.31
X$26911 384 608 385 644 645 cell_1rw
* cell instance $26912 m0 *1 112.095,131.04
X$26912 384 610 385 644 645 cell_1rw
* cell instance $26913 r0 *1 112.095,131.04
X$26913 384 611 385 644 645 cell_1rw
* cell instance $26914 m0 *1 112.095,133.77
X$26914 384 612 385 644 645 cell_1rw
* cell instance $26915 r0 *1 112.095,133.77
X$26915 384 613 385 644 645 cell_1rw
* cell instance $26916 m0 *1 112.095,136.5
X$26916 384 615 385 644 645 cell_1rw
* cell instance $26917 r0 *1 112.095,136.5
X$26917 384 614 385 644 645 cell_1rw
* cell instance $26918 m0 *1 112.095,139.23
X$26918 384 617 385 644 645 cell_1rw
* cell instance $26919 r0 *1 112.095,139.23
X$26919 384 616 385 644 645 cell_1rw
* cell instance $26920 m0 *1 112.095,141.96
X$26920 384 618 385 644 645 cell_1rw
* cell instance $26921 r0 *1 112.095,141.96
X$26921 384 619 385 644 645 cell_1rw
* cell instance $26922 m0 *1 112.095,144.69
X$26922 384 620 385 644 645 cell_1rw
* cell instance $26923 r0 *1 112.095,144.69
X$26923 384 621 385 644 645 cell_1rw
* cell instance $26924 m0 *1 112.095,147.42
X$26924 384 622 385 644 645 cell_1rw
* cell instance $26925 r0 *1 112.095,147.42
X$26925 384 623 385 644 645 cell_1rw
* cell instance $26926 m0 *1 112.095,150.15
X$26926 384 624 385 644 645 cell_1rw
* cell instance $26927 r0 *1 112.095,150.15
X$26927 384 625 385 644 645 cell_1rw
* cell instance $26928 m0 *1 112.095,152.88
X$26928 384 626 385 644 645 cell_1rw
* cell instance $26929 r0 *1 112.095,152.88
X$26929 384 627 385 644 645 cell_1rw
* cell instance $26930 m0 *1 112.095,155.61
X$26930 384 628 385 644 645 cell_1rw
* cell instance $26931 r0 *1 112.095,155.61
X$26931 384 629 385 644 645 cell_1rw
* cell instance $26932 m0 *1 112.095,158.34
X$26932 384 630 385 644 645 cell_1rw
* cell instance $26933 m0 *1 112.095,161.07
X$26933 384 632 385 644 645 cell_1rw
* cell instance $26934 r0 *1 112.095,158.34
X$26934 384 631 385 644 645 cell_1rw
* cell instance $26935 r0 *1 112.095,161.07
X$26935 384 633 385 644 645 cell_1rw
* cell instance $26936 m0 *1 112.095,163.8
X$26936 384 634 385 644 645 cell_1rw
* cell instance $26937 r0 *1 112.095,163.8
X$26937 384 635 385 644 645 cell_1rw
* cell instance $26938 m0 *1 112.095,166.53
X$26938 384 637 385 644 645 cell_1rw
* cell instance $26939 r0 *1 112.095,166.53
X$26939 384 636 385 644 645 cell_1rw
* cell instance $26940 m0 *1 112.095,169.26
X$26940 384 639 385 644 645 cell_1rw
* cell instance $26941 r0 *1 112.095,169.26
X$26941 384 638 385 644 645 cell_1rw
* cell instance $26942 m0 *1 112.095,171.99
X$26942 384 640 385 644 645 cell_1rw
* cell instance $26943 r0 *1 112.095,171.99
X$26943 384 641 385 644 645 cell_1rw
* cell instance $26944 m0 *1 112.095,174.72
X$26944 384 642 385 644 645 cell_1rw
* cell instance $26945 r0 *1 112.095,174.72
X$26945 384 643 385 644 645 cell_1rw
* cell instance $26946 m0 *1 112.8,90.09
X$26946 386 581 387 644 645 cell_1rw
* cell instance $26947 r0 *1 112.8,90.09
X$26947 386 580 387 644 645 cell_1rw
* cell instance $26948 m0 *1 112.8,92.82
X$26948 386 583 387 644 645 cell_1rw
* cell instance $26949 r0 *1 112.8,92.82
X$26949 386 582 387 644 645 cell_1rw
* cell instance $26950 m0 *1 112.8,95.55
X$26950 386 584 387 644 645 cell_1rw
* cell instance $26951 r0 *1 112.8,95.55
X$26951 386 585 387 644 645 cell_1rw
* cell instance $26952 m0 *1 112.8,98.28
X$26952 386 586 387 644 645 cell_1rw
* cell instance $26953 r0 *1 112.8,98.28
X$26953 386 587 387 644 645 cell_1rw
* cell instance $26954 m0 *1 112.8,101.01
X$26954 386 588 387 644 645 cell_1rw
* cell instance $26955 r0 *1 112.8,101.01
X$26955 386 589 387 644 645 cell_1rw
* cell instance $26956 m0 *1 112.8,103.74
X$26956 386 590 387 644 645 cell_1rw
* cell instance $26957 r0 *1 112.8,103.74
X$26957 386 591 387 644 645 cell_1rw
* cell instance $26958 m0 *1 112.8,106.47
X$26958 386 593 387 644 645 cell_1rw
* cell instance $26959 r0 *1 112.8,106.47
X$26959 386 592 387 644 645 cell_1rw
* cell instance $26960 m0 *1 112.8,109.2
X$26960 386 594 387 644 645 cell_1rw
* cell instance $26961 m0 *1 112.8,111.93
X$26961 386 597 387 644 645 cell_1rw
* cell instance $26962 r0 *1 112.8,109.2
X$26962 386 595 387 644 645 cell_1rw
* cell instance $26963 r0 *1 112.8,111.93
X$26963 386 596 387 644 645 cell_1rw
* cell instance $26964 m0 *1 112.8,114.66
X$26964 386 598 387 644 645 cell_1rw
* cell instance $26965 m0 *1 112.8,117.39
X$26965 386 600 387 644 645 cell_1rw
* cell instance $26966 r0 *1 112.8,114.66
X$26966 386 599 387 644 645 cell_1rw
* cell instance $26967 m0 *1 112.8,120.12
X$26967 386 602 387 644 645 cell_1rw
* cell instance $26968 r0 *1 112.8,117.39
X$26968 386 601 387 644 645 cell_1rw
* cell instance $26969 r0 *1 112.8,120.12
X$26969 386 603 387 644 645 cell_1rw
* cell instance $26970 m0 *1 112.8,122.85
X$26970 386 604 387 644 645 cell_1rw
* cell instance $26971 m0 *1 112.8,125.58
X$26971 386 606 387 644 645 cell_1rw
* cell instance $26972 r0 *1 112.8,122.85
X$26972 386 605 387 644 645 cell_1rw
* cell instance $26973 r0 *1 112.8,125.58
X$26973 386 607 387 644 645 cell_1rw
* cell instance $26974 m0 *1 112.8,128.31
X$26974 386 609 387 644 645 cell_1rw
* cell instance $26975 r0 *1 112.8,128.31
X$26975 386 608 387 644 645 cell_1rw
* cell instance $26976 m0 *1 112.8,131.04
X$26976 386 610 387 644 645 cell_1rw
* cell instance $26977 r0 *1 112.8,131.04
X$26977 386 611 387 644 645 cell_1rw
* cell instance $26978 m0 *1 112.8,133.77
X$26978 386 612 387 644 645 cell_1rw
* cell instance $26979 r0 *1 112.8,133.77
X$26979 386 613 387 644 645 cell_1rw
* cell instance $26980 m0 *1 112.8,136.5
X$26980 386 615 387 644 645 cell_1rw
* cell instance $26981 m0 *1 112.8,139.23
X$26981 386 617 387 644 645 cell_1rw
* cell instance $26982 r0 *1 112.8,136.5
X$26982 386 614 387 644 645 cell_1rw
* cell instance $26983 r0 *1 112.8,139.23
X$26983 386 616 387 644 645 cell_1rw
* cell instance $26984 m0 *1 112.8,141.96
X$26984 386 618 387 644 645 cell_1rw
* cell instance $26985 r0 *1 112.8,141.96
X$26985 386 619 387 644 645 cell_1rw
* cell instance $26986 m0 *1 112.8,144.69
X$26986 386 620 387 644 645 cell_1rw
* cell instance $26987 r0 *1 112.8,144.69
X$26987 386 621 387 644 645 cell_1rw
* cell instance $26988 m0 *1 112.8,147.42
X$26988 386 622 387 644 645 cell_1rw
* cell instance $26989 m0 *1 112.8,150.15
X$26989 386 624 387 644 645 cell_1rw
* cell instance $26990 r0 *1 112.8,147.42
X$26990 386 623 387 644 645 cell_1rw
* cell instance $26991 r0 *1 112.8,150.15
X$26991 386 625 387 644 645 cell_1rw
* cell instance $26992 m0 *1 112.8,152.88
X$26992 386 626 387 644 645 cell_1rw
* cell instance $26993 r0 *1 112.8,152.88
X$26993 386 627 387 644 645 cell_1rw
* cell instance $26994 m0 *1 112.8,155.61
X$26994 386 628 387 644 645 cell_1rw
* cell instance $26995 r0 *1 112.8,155.61
X$26995 386 629 387 644 645 cell_1rw
* cell instance $26996 m0 *1 112.8,158.34
X$26996 386 630 387 644 645 cell_1rw
* cell instance $26997 r0 *1 112.8,158.34
X$26997 386 631 387 644 645 cell_1rw
* cell instance $26998 m0 *1 112.8,161.07
X$26998 386 632 387 644 645 cell_1rw
* cell instance $26999 r0 *1 112.8,161.07
X$26999 386 633 387 644 645 cell_1rw
* cell instance $27000 m0 *1 112.8,163.8
X$27000 386 634 387 644 645 cell_1rw
* cell instance $27001 r0 *1 112.8,163.8
X$27001 386 635 387 644 645 cell_1rw
* cell instance $27002 m0 *1 112.8,166.53
X$27002 386 637 387 644 645 cell_1rw
* cell instance $27003 r0 *1 112.8,166.53
X$27003 386 636 387 644 645 cell_1rw
* cell instance $27004 m0 *1 112.8,169.26
X$27004 386 639 387 644 645 cell_1rw
* cell instance $27005 r0 *1 112.8,169.26
X$27005 386 638 387 644 645 cell_1rw
* cell instance $27006 m0 *1 112.8,171.99
X$27006 386 640 387 644 645 cell_1rw
* cell instance $27007 r0 *1 112.8,171.99
X$27007 386 641 387 644 645 cell_1rw
* cell instance $27008 m0 *1 112.8,174.72
X$27008 386 642 387 644 645 cell_1rw
* cell instance $27009 r0 *1 112.8,174.72
X$27009 386 643 387 644 645 cell_1rw
* cell instance $27010 m0 *1 113.505,90.09
X$27010 388 581 389 644 645 cell_1rw
* cell instance $27011 r0 *1 113.505,90.09
X$27011 388 580 389 644 645 cell_1rw
* cell instance $27012 m0 *1 113.505,92.82
X$27012 388 583 389 644 645 cell_1rw
* cell instance $27013 m0 *1 113.505,95.55
X$27013 388 584 389 644 645 cell_1rw
* cell instance $27014 r0 *1 113.505,92.82
X$27014 388 582 389 644 645 cell_1rw
* cell instance $27015 r0 *1 113.505,95.55
X$27015 388 585 389 644 645 cell_1rw
* cell instance $27016 m0 *1 113.505,98.28
X$27016 388 586 389 644 645 cell_1rw
* cell instance $27017 r0 *1 113.505,98.28
X$27017 388 587 389 644 645 cell_1rw
* cell instance $27018 m0 *1 113.505,101.01
X$27018 388 588 389 644 645 cell_1rw
* cell instance $27019 r0 *1 113.505,101.01
X$27019 388 589 389 644 645 cell_1rw
* cell instance $27020 m0 *1 113.505,103.74
X$27020 388 590 389 644 645 cell_1rw
* cell instance $27021 r0 *1 113.505,103.74
X$27021 388 591 389 644 645 cell_1rw
* cell instance $27022 m0 *1 113.505,106.47
X$27022 388 593 389 644 645 cell_1rw
* cell instance $27023 m0 *1 113.505,109.2
X$27023 388 594 389 644 645 cell_1rw
* cell instance $27024 r0 *1 113.505,106.47
X$27024 388 592 389 644 645 cell_1rw
* cell instance $27025 r0 *1 113.505,109.2
X$27025 388 595 389 644 645 cell_1rw
* cell instance $27026 m0 *1 113.505,111.93
X$27026 388 597 389 644 645 cell_1rw
* cell instance $27027 r0 *1 113.505,111.93
X$27027 388 596 389 644 645 cell_1rw
* cell instance $27028 m0 *1 113.505,114.66
X$27028 388 598 389 644 645 cell_1rw
* cell instance $27029 m0 *1 113.505,117.39
X$27029 388 600 389 644 645 cell_1rw
* cell instance $27030 r0 *1 113.505,114.66
X$27030 388 599 389 644 645 cell_1rw
* cell instance $27031 r0 *1 113.505,117.39
X$27031 388 601 389 644 645 cell_1rw
* cell instance $27032 m0 *1 113.505,120.12
X$27032 388 602 389 644 645 cell_1rw
* cell instance $27033 r0 *1 113.505,120.12
X$27033 388 603 389 644 645 cell_1rw
* cell instance $27034 m0 *1 113.505,122.85
X$27034 388 604 389 644 645 cell_1rw
* cell instance $27035 r0 *1 113.505,122.85
X$27035 388 605 389 644 645 cell_1rw
* cell instance $27036 m0 *1 113.505,125.58
X$27036 388 606 389 644 645 cell_1rw
* cell instance $27037 r0 *1 113.505,125.58
X$27037 388 607 389 644 645 cell_1rw
* cell instance $27038 m0 *1 113.505,128.31
X$27038 388 609 389 644 645 cell_1rw
* cell instance $27039 r0 *1 113.505,128.31
X$27039 388 608 389 644 645 cell_1rw
* cell instance $27040 m0 *1 113.505,131.04
X$27040 388 610 389 644 645 cell_1rw
* cell instance $27041 r0 *1 113.505,131.04
X$27041 388 611 389 644 645 cell_1rw
* cell instance $27042 m0 *1 113.505,133.77
X$27042 388 612 389 644 645 cell_1rw
* cell instance $27043 m0 *1 113.505,136.5
X$27043 388 615 389 644 645 cell_1rw
* cell instance $27044 r0 *1 113.505,133.77
X$27044 388 613 389 644 645 cell_1rw
* cell instance $27045 r0 *1 113.505,136.5
X$27045 388 614 389 644 645 cell_1rw
* cell instance $27046 m0 *1 113.505,139.23
X$27046 388 617 389 644 645 cell_1rw
* cell instance $27047 r0 *1 113.505,139.23
X$27047 388 616 389 644 645 cell_1rw
* cell instance $27048 m0 *1 113.505,141.96
X$27048 388 618 389 644 645 cell_1rw
* cell instance $27049 r0 *1 113.505,141.96
X$27049 388 619 389 644 645 cell_1rw
* cell instance $27050 m0 *1 113.505,144.69
X$27050 388 620 389 644 645 cell_1rw
* cell instance $27051 m0 *1 113.505,147.42
X$27051 388 622 389 644 645 cell_1rw
* cell instance $27052 r0 *1 113.505,144.69
X$27052 388 621 389 644 645 cell_1rw
* cell instance $27053 r0 *1 113.505,147.42
X$27053 388 623 389 644 645 cell_1rw
* cell instance $27054 m0 *1 113.505,150.15
X$27054 388 624 389 644 645 cell_1rw
* cell instance $27055 r0 *1 113.505,150.15
X$27055 388 625 389 644 645 cell_1rw
* cell instance $27056 m0 *1 113.505,152.88
X$27056 388 626 389 644 645 cell_1rw
* cell instance $27057 m0 *1 113.505,155.61
X$27057 388 628 389 644 645 cell_1rw
* cell instance $27058 r0 *1 113.505,152.88
X$27058 388 627 389 644 645 cell_1rw
* cell instance $27059 r0 *1 113.505,155.61
X$27059 388 629 389 644 645 cell_1rw
* cell instance $27060 m0 *1 113.505,158.34
X$27060 388 630 389 644 645 cell_1rw
* cell instance $27061 r0 *1 113.505,158.34
X$27061 388 631 389 644 645 cell_1rw
* cell instance $27062 m0 *1 113.505,161.07
X$27062 388 632 389 644 645 cell_1rw
* cell instance $27063 r0 *1 113.505,161.07
X$27063 388 633 389 644 645 cell_1rw
* cell instance $27064 m0 *1 113.505,163.8
X$27064 388 634 389 644 645 cell_1rw
* cell instance $27065 m0 *1 113.505,166.53
X$27065 388 637 389 644 645 cell_1rw
* cell instance $27066 r0 *1 113.505,163.8
X$27066 388 635 389 644 645 cell_1rw
* cell instance $27067 m0 *1 113.505,169.26
X$27067 388 639 389 644 645 cell_1rw
* cell instance $27068 r0 *1 113.505,166.53
X$27068 388 636 389 644 645 cell_1rw
* cell instance $27069 r0 *1 113.505,169.26
X$27069 388 638 389 644 645 cell_1rw
* cell instance $27070 m0 *1 113.505,171.99
X$27070 388 640 389 644 645 cell_1rw
* cell instance $27071 r0 *1 113.505,171.99
X$27071 388 641 389 644 645 cell_1rw
* cell instance $27072 m0 *1 113.505,174.72
X$27072 388 642 389 644 645 cell_1rw
* cell instance $27073 r0 *1 113.505,174.72
X$27073 388 643 389 644 645 cell_1rw
* cell instance $27074 m0 *1 114.21,90.09
X$27074 390 581 391 644 645 cell_1rw
* cell instance $27075 r0 *1 114.21,90.09
X$27075 390 580 391 644 645 cell_1rw
* cell instance $27076 m0 *1 114.21,92.82
X$27076 390 583 391 644 645 cell_1rw
* cell instance $27077 m0 *1 114.21,95.55
X$27077 390 584 391 644 645 cell_1rw
* cell instance $27078 r0 *1 114.21,92.82
X$27078 390 582 391 644 645 cell_1rw
* cell instance $27079 m0 *1 114.21,98.28
X$27079 390 586 391 644 645 cell_1rw
* cell instance $27080 r0 *1 114.21,95.55
X$27080 390 585 391 644 645 cell_1rw
* cell instance $27081 r0 *1 114.21,98.28
X$27081 390 587 391 644 645 cell_1rw
* cell instance $27082 m0 *1 114.21,101.01
X$27082 390 588 391 644 645 cell_1rw
* cell instance $27083 r0 *1 114.21,101.01
X$27083 390 589 391 644 645 cell_1rw
* cell instance $27084 m0 *1 114.21,103.74
X$27084 390 590 391 644 645 cell_1rw
* cell instance $27085 r0 *1 114.21,103.74
X$27085 390 591 391 644 645 cell_1rw
* cell instance $27086 m0 *1 114.21,106.47
X$27086 390 593 391 644 645 cell_1rw
* cell instance $27087 r0 *1 114.21,106.47
X$27087 390 592 391 644 645 cell_1rw
* cell instance $27088 m0 *1 114.21,109.2
X$27088 390 594 391 644 645 cell_1rw
* cell instance $27089 r0 *1 114.21,109.2
X$27089 390 595 391 644 645 cell_1rw
* cell instance $27090 m0 *1 114.21,111.93
X$27090 390 597 391 644 645 cell_1rw
* cell instance $27091 r0 *1 114.21,111.93
X$27091 390 596 391 644 645 cell_1rw
* cell instance $27092 m0 *1 114.21,114.66
X$27092 390 598 391 644 645 cell_1rw
* cell instance $27093 r0 *1 114.21,114.66
X$27093 390 599 391 644 645 cell_1rw
* cell instance $27094 m0 *1 114.21,117.39
X$27094 390 600 391 644 645 cell_1rw
* cell instance $27095 r0 *1 114.21,117.39
X$27095 390 601 391 644 645 cell_1rw
* cell instance $27096 m0 *1 114.21,120.12
X$27096 390 602 391 644 645 cell_1rw
* cell instance $27097 r0 *1 114.21,120.12
X$27097 390 603 391 644 645 cell_1rw
* cell instance $27098 m0 *1 114.21,122.85
X$27098 390 604 391 644 645 cell_1rw
* cell instance $27099 r0 *1 114.21,122.85
X$27099 390 605 391 644 645 cell_1rw
* cell instance $27100 m0 *1 114.21,125.58
X$27100 390 606 391 644 645 cell_1rw
* cell instance $27101 r0 *1 114.21,125.58
X$27101 390 607 391 644 645 cell_1rw
* cell instance $27102 m0 *1 114.21,128.31
X$27102 390 609 391 644 645 cell_1rw
* cell instance $27103 r0 *1 114.21,128.31
X$27103 390 608 391 644 645 cell_1rw
* cell instance $27104 m0 *1 114.21,131.04
X$27104 390 610 391 644 645 cell_1rw
* cell instance $27105 r0 *1 114.21,131.04
X$27105 390 611 391 644 645 cell_1rw
* cell instance $27106 m0 *1 114.21,133.77
X$27106 390 612 391 644 645 cell_1rw
* cell instance $27107 r0 *1 114.21,133.77
X$27107 390 613 391 644 645 cell_1rw
* cell instance $27108 m0 *1 114.21,136.5
X$27108 390 615 391 644 645 cell_1rw
* cell instance $27109 r0 *1 114.21,136.5
X$27109 390 614 391 644 645 cell_1rw
* cell instance $27110 m0 *1 114.21,139.23
X$27110 390 617 391 644 645 cell_1rw
* cell instance $27111 r0 *1 114.21,139.23
X$27111 390 616 391 644 645 cell_1rw
* cell instance $27112 m0 *1 114.21,141.96
X$27112 390 618 391 644 645 cell_1rw
* cell instance $27113 r0 *1 114.21,141.96
X$27113 390 619 391 644 645 cell_1rw
* cell instance $27114 m0 *1 114.21,144.69
X$27114 390 620 391 644 645 cell_1rw
* cell instance $27115 m0 *1 114.21,147.42
X$27115 390 622 391 644 645 cell_1rw
* cell instance $27116 r0 *1 114.21,144.69
X$27116 390 621 391 644 645 cell_1rw
* cell instance $27117 r0 *1 114.21,147.42
X$27117 390 623 391 644 645 cell_1rw
* cell instance $27118 m0 *1 114.21,150.15
X$27118 390 624 391 644 645 cell_1rw
* cell instance $27119 m0 *1 114.21,152.88
X$27119 390 626 391 644 645 cell_1rw
* cell instance $27120 r0 *1 114.21,150.15
X$27120 390 625 391 644 645 cell_1rw
* cell instance $27121 r0 *1 114.21,152.88
X$27121 390 627 391 644 645 cell_1rw
* cell instance $27122 m0 *1 114.21,155.61
X$27122 390 628 391 644 645 cell_1rw
* cell instance $27123 m0 *1 114.21,158.34
X$27123 390 630 391 644 645 cell_1rw
* cell instance $27124 r0 *1 114.21,155.61
X$27124 390 629 391 644 645 cell_1rw
* cell instance $27125 m0 *1 114.21,161.07
X$27125 390 632 391 644 645 cell_1rw
* cell instance $27126 r0 *1 114.21,158.34
X$27126 390 631 391 644 645 cell_1rw
* cell instance $27127 r0 *1 114.21,161.07
X$27127 390 633 391 644 645 cell_1rw
* cell instance $27128 m0 *1 114.21,163.8
X$27128 390 634 391 644 645 cell_1rw
* cell instance $27129 r0 *1 114.21,163.8
X$27129 390 635 391 644 645 cell_1rw
* cell instance $27130 m0 *1 114.21,166.53
X$27130 390 637 391 644 645 cell_1rw
* cell instance $27131 r0 *1 114.21,166.53
X$27131 390 636 391 644 645 cell_1rw
* cell instance $27132 m0 *1 114.21,169.26
X$27132 390 639 391 644 645 cell_1rw
* cell instance $27133 r0 *1 114.21,169.26
X$27133 390 638 391 644 645 cell_1rw
* cell instance $27134 m0 *1 114.21,171.99
X$27134 390 640 391 644 645 cell_1rw
* cell instance $27135 m0 *1 114.21,174.72
X$27135 390 642 391 644 645 cell_1rw
* cell instance $27136 r0 *1 114.21,171.99
X$27136 390 641 391 644 645 cell_1rw
* cell instance $27137 r0 *1 114.21,174.72
X$27137 390 643 391 644 645 cell_1rw
* cell instance $27138 m0 *1 114.915,90.09
X$27138 392 581 393 644 645 cell_1rw
* cell instance $27139 r0 *1 114.915,90.09
X$27139 392 580 393 644 645 cell_1rw
* cell instance $27140 m0 *1 114.915,92.82
X$27140 392 583 393 644 645 cell_1rw
* cell instance $27141 r0 *1 114.915,92.82
X$27141 392 582 393 644 645 cell_1rw
* cell instance $27142 m0 *1 114.915,95.55
X$27142 392 584 393 644 645 cell_1rw
* cell instance $27143 m0 *1 114.915,98.28
X$27143 392 586 393 644 645 cell_1rw
* cell instance $27144 r0 *1 114.915,95.55
X$27144 392 585 393 644 645 cell_1rw
* cell instance $27145 m0 *1 114.915,101.01
X$27145 392 588 393 644 645 cell_1rw
* cell instance $27146 r0 *1 114.915,98.28
X$27146 392 587 393 644 645 cell_1rw
* cell instance $27147 r0 *1 114.915,101.01
X$27147 392 589 393 644 645 cell_1rw
* cell instance $27148 m0 *1 114.915,103.74
X$27148 392 590 393 644 645 cell_1rw
* cell instance $27149 r0 *1 114.915,103.74
X$27149 392 591 393 644 645 cell_1rw
* cell instance $27150 m0 *1 114.915,106.47
X$27150 392 593 393 644 645 cell_1rw
* cell instance $27151 r0 *1 114.915,106.47
X$27151 392 592 393 644 645 cell_1rw
* cell instance $27152 m0 *1 114.915,109.2
X$27152 392 594 393 644 645 cell_1rw
* cell instance $27153 m0 *1 114.915,111.93
X$27153 392 597 393 644 645 cell_1rw
* cell instance $27154 r0 *1 114.915,109.2
X$27154 392 595 393 644 645 cell_1rw
* cell instance $27155 r0 *1 114.915,111.93
X$27155 392 596 393 644 645 cell_1rw
* cell instance $27156 m0 *1 114.915,114.66
X$27156 392 598 393 644 645 cell_1rw
* cell instance $27157 r0 *1 114.915,114.66
X$27157 392 599 393 644 645 cell_1rw
* cell instance $27158 m0 *1 114.915,117.39
X$27158 392 600 393 644 645 cell_1rw
* cell instance $27159 r0 *1 114.915,117.39
X$27159 392 601 393 644 645 cell_1rw
* cell instance $27160 m0 *1 114.915,120.12
X$27160 392 602 393 644 645 cell_1rw
* cell instance $27161 r0 *1 114.915,120.12
X$27161 392 603 393 644 645 cell_1rw
* cell instance $27162 m0 *1 114.915,122.85
X$27162 392 604 393 644 645 cell_1rw
* cell instance $27163 r0 *1 114.915,122.85
X$27163 392 605 393 644 645 cell_1rw
* cell instance $27164 m0 *1 114.915,125.58
X$27164 392 606 393 644 645 cell_1rw
* cell instance $27165 r0 *1 114.915,125.58
X$27165 392 607 393 644 645 cell_1rw
* cell instance $27166 m0 *1 114.915,128.31
X$27166 392 609 393 644 645 cell_1rw
* cell instance $27167 r0 *1 114.915,128.31
X$27167 392 608 393 644 645 cell_1rw
* cell instance $27168 m0 *1 114.915,131.04
X$27168 392 610 393 644 645 cell_1rw
* cell instance $27169 r0 *1 114.915,131.04
X$27169 392 611 393 644 645 cell_1rw
* cell instance $27170 m0 *1 114.915,133.77
X$27170 392 612 393 644 645 cell_1rw
* cell instance $27171 r0 *1 114.915,133.77
X$27171 392 613 393 644 645 cell_1rw
* cell instance $27172 m0 *1 114.915,136.5
X$27172 392 615 393 644 645 cell_1rw
* cell instance $27173 r0 *1 114.915,136.5
X$27173 392 614 393 644 645 cell_1rw
* cell instance $27174 m0 *1 114.915,139.23
X$27174 392 617 393 644 645 cell_1rw
* cell instance $27175 m0 *1 114.915,141.96
X$27175 392 618 393 644 645 cell_1rw
* cell instance $27176 r0 *1 114.915,139.23
X$27176 392 616 393 644 645 cell_1rw
* cell instance $27177 m0 *1 114.915,144.69
X$27177 392 620 393 644 645 cell_1rw
* cell instance $27178 r0 *1 114.915,141.96
X$27178 392 619 393 644 645 cell_1rw
* cell instance $27179 r0 *1 114.915,144.69
X$27179 392 621 393 644 645 cell_1rw
* cell instance $27180 m0 *1 114.915,147.42
X$27180 392 622 393 644 645 cell_1rw
* cell instance $27181 r0 *1 114.915,147.42
X$27181 392 623 393 644 645 cell_1rw
* cell instance $27182 m0 *1 114.915,150.15
X$27182 392 624 393 644 645 cell_1rw
* cell instance $27183 r0 *1 114.915,150.15
X$27183 392 625 393 644 645 cell_1rw
* cell instance $27184 m0 *1 114.915,152.88
X$27184 392 626 393 644 645 cell_1rw
* cell instance $27185 r0 *1 114.915,152.88
X$27185 392 627 393 644 645 cell_1rw
* cell instance $27186 m0 *1 114.915,155.61
X$27186 392 628 393 644 645 cell_1rw
* cell instance $27187 r0 *1 114.915,155.61
X$27187 392 629 393 644 645 cell_1rw
* cell instance $27188 m0 *1 114.915,158.34
X$27188 392 630 393 644 645 cell_1rw
* cell instance $27189 r0 *1 114.915,158.34
X$27189 392 631 393 644 645 cell_1rw
* cell instance $27190 m0 *1 114.915,161.07
X$27190 392 632 393 644 645 cell_1rw
* cell instance $27191 r0 *1 114.915,161.07
X$27191 392 633 393 644 645 cell_1rw
* cell instance $27192 m0 *1 114.915,163.8
X$27192 392 634 393 644 645 cell_1rw
* cell instance $27193 m0 *1 114.915,166.53
X$27193 392 637 393 644 645 cell_1rw
* cell instance $27194 r0 *1 114.915,163.8
X$27194 392 635 393 644 645 cell_1rw
* cell instance $27195 r0 *1 114.915,166.53
X$27195 392 636 393 644 645 cell_1rw
* cell instance $27196 m0 *1 114.915,169.26
X$27196 392 639 393 644 645 cell_1rw
* cell instance $27197 r0 *1 114.915,169.26
X$27197 392 638 393 644 645 cell_1rw
* cell instance $27198 m0 *1 114.915,171.99
X$27198 392 640 393 644 645 cell_1rw
* cell instance $27199 r0 *1 114.915,171.99
X$27199 392 641 393 644 645 cell_1rw
* cell instance $27200 m0 *1 114.915,174.72
X$27200 392 642 393 644 645 cell_1rw
* cell instance $27201 r0 *1 114.915,174.72
X$27201 392 643 393 644 645 cell_1rw
* cell instance $27202 m0 *1 115.62,90.09
X$27202 394 581 395 644 645 cell_1rw
* cell instance $27203 r0 *1 115.62,90.09
X$27203 394 580 395 644 645 cell_1rw
* cell instance $27204 m0 *1 115.62,92.82
X$27204 394 583 395 644 645 cell_1rw
* cell instance $27205 m0 *1 115.62,95.55
X$27205 394 584 395 644 645 cell_1rw
* cell instance $27206 r0 *1 115.62,92.82
X$27206 394 582 395 644 645 cell_1rw
* cell instance $27207 r0 *1 115.62,95.55
X$27207 394 585 395 644 645 cell_1rw
* cell instance $27208 m0 *1 115.62,98.28
X$27208 394 586 395 644 645 cell_1rw
* cell instance $27209 r0 *1 115.62,98.28
X$27209 394 587 395 644 645 cell_1rw
* cell instance $27210 m0 *1 115.62,101.01
X$27210 394 588 395 644 645 cell_1rw
* cell instance $27211 r0 *1 115.62,101.01
X$27211 394 589 395 644 645 cell_1rw
* cell instance $27212 m0 *1 115.62,103.74
X$27212 394 590 395 644 645 cell_1rw
* cell instance $27213 r0 *1 115.62,103.74
X$27213 394 591 395 644 645 cell_1rw
* cell instance $27214 m0 *1 115.62,106.47
X$27214 394 593 395 644 645 cell_1rw
* cell instance $27215 r0 *1 115.62,106.47
X$27215 394 592 395 644 645 cell_1rw
* cell instance $27216 m0 *1 115.62,109.2
X$27216 394 594 395 644 645 cell_1rw
* cell instance $27217 m0 *1 115.62,111.93
X$27217 394 597 395 644 645 cell_1rw
* cell instance $27218 r0 *1 115.62,109.2
X$27218 394 595 395 644 645 cell_1rw
* cell instance $27219 r0 *1 115.62,111.93
X$27219 394 596 395 644 645 cell_1rw
* cell instance $27220 m0 *1 115.62,114.66
X$27220 394 598 395 644 645 cell_1rw
* cell instance $27221 r0 *1 115.62,114.66
X$27221 394 599 395 644 645 cell_1rw
* cell instance $27222 m0 *1 115.62,117.39
X$27222 394 600 395 644 645 cell_1rw
* cell instance $27223 r0 *1 115.62,117.39
X$27223 394 601 395 644 645 cell_1rw
* cell instance $27224 m0 *1 115.62,120.12
X$27224 394 602 395 644 645 cell_1rw
* cell instance $27225 r0 *1 115.62,120.12
X$27225 394 603 395 644 645 cell_1rw
* cell instance $27226 m0 *1 115.62,122.85
X$27226 394 604 395 644 645 cell_1rw
* cell instance $27227 r0 *1 115.62,122.85
X$27227 394 605 395 644 645 cell_1rw
* cell instance $27228 m0 *1 115.62,125.58
X$27228 394 606 395 644 645 cell_1rw
* cell instance $27229 r0 *1 115.62,125.58
X$27229 394 607 395 644 645 cell_1rw
* cell instance $27230 m0 *1 115.62,128.31
X$27230 394 609 395 644 645 cell_1rw
* cell instance $27231 r0 *1 115.62,128.31
X$27231 394 608 395 644 645 cell_1rw
* cell instance $27232 m0 *1 115.62,131.04
X$27232 394 610 395 644 645 cell_1rw
* cell instance $27233 r0 *1 115.62,131.04
X$27233 394 611 395 644 645 cell_1rw
* cell instance $27234 m0 *1 115.62,133.77
X$27234 394 612 395 644 645 cell_1rw
* cell instance $27235 r0 *1 115.62,133.77
X$27235 394 613 395 644 645 cell_1rw
* cell instance $27236 m0 *1 115.62,136.5
X$27236 394 615 395 644 645 cell_1rw
* cell instance $27237 r0 *1 115.62,136.5
X$27237 394 614 395 644 645 cell_1rw
* cell instance $27238 m0 *1 115.62,139.23
X$27238 394 617 395 644 645 cell_1rw
* cell instance $27239 r0 *1 115.62,139.23
X$27239 394 616 395 644 645 cell_1rw
* cell instance $27240 m0 *1 115.62,141.96
X$27240 394 618 395 644 645 cell_1rw
* cell instance $27241 r0 *1 115.62,141.96
X$27241 394 619 395 644 645 cell_1rw
* cell instance $27242 m0 *1 115.62,144.69
X$27242 394 620 395 644 645 cell_1rw
* cell instance $27243 r0 *1 115.62,144.69
X$27243 394 621 395 644 645 cell_1rw
* cell instance $27244 m0 *1 115.62,147.42
X$27244 394 622 395 644 645 cell_1rw
* cell instance $27245 r0 *1 115.62,147.42
X$27245 394 623 395 644 645 cell_1rw
* cell instance $27246 m0 *1 115.62,150.15
X$27246 394 624 395 644 645 cell_1rw
* cell instance $27247 m0 *1 115.62,152.88
X$27247 394 626 395 644 645 cell_1rw
* cell instance $27248 r0 *1 115.62,150.15
X$27248 394 625 395 644 645 cell_1rw
* cell instance $27249 m0 *1 115.62,155.61
X$27249 394 628 395 644 645 cell_1rw
* cell instance $27250 r0 *1 115.62,152.88
X$27250 394 627 395 644 645 cell_1rw
* cell instance $27251 m0 *1 115.62,158.34
X$27251 394 630 395 644 645 cell_1rw
* cell instance $27252 r0 *1 115.62,155.61
X$27252 394 629 395 644 645 cell_1rw
* cell instance $27253 r0 *1 115.62,158.34
X$27253 394 631 395 644 645 cell_1rw
* cell instance $27254 m0 *1 115.62,161.07
X$27254 394 632 395 644 645 cell_1rw
* cell instance $27255 r0 *1 115.62,161.07
X$27255 394 633 395 644 645 cell_1rw
* cell instance $27256 m0 *1 115.62,163.8
X$27256 394 634 395 644 645 cell_1rw
* cell instance $27257 r0 *1 115.62,163.8
X$27257 394 635 395 644 645 cell_1rw
* cell instance $27258 m0 *1 115.62,166.53
X$27258 394 637 395 644 645 cell_1rw
* cell instance $27259 r0 *1 115.62,166.53
X$27259 394 636 395 644 645 cell_1rw
* cell instance $27260 m0 *1 115.62,169.26
X$27260 394 639 395 644 645 cell_1rw
* cell instance $27261 r0 *1 115.62,169.26
X$27261 394 638 395 644 645 cell_1rw
* cell instance $27262 m0 *1 115.62,171.99
X$27262 394 640 395 644 645 cell_1rw
* cell instance $27263 r0 *1 115.62,171.99
X$27263 394 641 395 644 645 cell_1rw
* cell instance $27264 m0 *1 115.62,174.72
X$27264 394 642 395 644 645 cell_1rw
* cell instance $27265 r0 *1 115.62,174.72
X$27265 394 643 395 644 645 cell_1rw
* cell instance $27266 m0 *1 116.325,90.09
X$27266 396 581 397 644 645 cell_1rw
* cell instance $27267 r0 *1 116.325,90.09
X$27267 396 580 397 644 645 cell_1rw
* cell instance $27268 m0 *1 116.325,92.82
X$27268 396 583 397 644 645 cell_1rw
* cell instance $27269 r0 *1 116.325,92.82
X$27269 396 582 397 644 645 cell_1rw
* cell instance $27270 m0 *1 116.325,95.55
X$27270 396 584 397 644 645 cell_1rw
* cell instance $27271 r0 *1 116.325,95.55
X$27271 396 585 397 644 645 cell_1rw
* cell instance $27272 m0 *1 116.325,98.28
X$27272 396 586 397 644 645 cell_1rw
* cell instance $27273 r0 *1 116.325,98.28
X$27273 396 587 397 644 645 cell_1rw
* cell instance $27274 m0 *1 116.325,101.01
X$27274 396 588 397 644 645 cell_1rw
* cell instance $27275 r0 *1 116.325,101.01
X$27275 396 589 397 644 645 cell_1rw
* cell instance $27276 m0 *1 116.325,103.74
X$27276 396 590 397 644 645 cell_1rw
* cell instance $27277 r0 *1 116.325,103.74
X$27277 396 591 397 644 645 cell_1rw
* cell instance $27278 m0 *1 116.325,106.47
X$27278 396 593 397 644 645 cell_1rw
* cell instance $27279 r0 *1 116.325,106.47
X$27279 396 592 397 644 645 cell_1rw
* cell instance $27280 m0 *1 116.325,109.2
X$27280 396 594 397 644 645 cell_1rw
* cell instance $27281 r0 *1 116.325,109.2
X$27281 396 595 397 644 645 cell_1rw
* cell instance $27282 m0 *1 116.325,111.93
X$27282 396 597 397 644 645 cell_1rw
* cell instance $27283 r0 *1 116.325,111.93
X$27283 396 596 397 644 645 cell_1rw
* cell instance $27284 m0 *1 116.325,114.66
X$27284 396 598 397 644 645 cell_1rw
* cell instance $27285 r0 *1 116.325,114.66
X$27285 396 599 397 644 645 cell_1rw
* cell instance $27286 m0 *1 116.325,117.39
X$27286 396 600 397 644 645 cell_1rw
* cell instance $27287 r0 *1 116.325,117.39
X$27287 396 601 397 644 645 cell_1rw
* cell instance $27288 m0 *1 116.325,120.12
X$27288 396 602 397 644 645 cell_1rw
* cell instance $27289 r0 *1 116.325,120.12
X$27289 396 603 397 644 645 cell_1rw
* cell instance $27290 m0 *1 116.325,122.85
X$27290 396 604 397 644 645 cell_1rw
* cell instance $27291 m0 *1 116.325,125.58
X$27291 396 606 397 644 645 cell_1rw
* cell instance $27292 r0 *1 116.325,122.85
X$27292 396 605 397 644 645 cell_1rw
* cell instance $27293 r0 *1 116.325,125.58
X$27293 396 607 397 644 645 cell_1rw
* cell instance $27294 m0 *1 116.325,128.31
X$27294 396 609 397 644 645 cell_1rw
* cell instance $27295 r0 *1 116.325,128.31
X$27295 396 608 397 644 645 cell_1rw
* cell instance $27296 m0 *1 116.325,131.04
X$27296 396 610 397 644 645 cell_1rw
* cell instance $27297 r0 *1 116.325,131.04
X$27297 396 611 397 644 645 cell_1rw
* cell instance $27298 m0 *1 116.325,133.77
X$27298 396 612 397 644 645 cell_1rw
* cell instance $27299 m0 *1 116.325,136.5
X$27299 396 615 397 644 645 cell_1rw
* cell instance $27300 r0 *1 116.325,133.77
X$27300 396 613 397 644 645 cell_1rw
* cell instance $27301 r0 *1 116.325,136.5
X$27301 396 614 397 644 645 cell_1rw
* cell instance $27302 m0 *1 116.325,139.23
X$27302 396 617 397 644 645 cell_1rw
* cell instance $27303 r0 *1 116.325,139.23
X$27303 396 616 397 644 645 cell_1rw
* cell instance $27304 m0 *1 116.325,141.96
X$27304 396 618 397 644 645 cell_1rw
* cell instance $27305 r0 *1 116.325,141.96
X$27305 396 619 397 644 645 cell_1rw
* cell instance $27306 m0 *1 116.325,144.69
X$27306 396 620 397 644 645 cell_1rw
* cell instance $27307 r0 *1 116.325,144.69
X$27307 396 621 397 644 645 cell_1rw
* cell instance $27308 m0 *1 116.325,147.42
X$27308 396 622 397 644 645 cell_1rw
* cell instance $27309 r0 *1 116.325,147.42
X$27309 396 623 397 644 645 cell_1rw
* cell instance $27310 m0 *1 116.325,150.15
X$27310 396 624 397 644 645 cell_1rw
* cell instance $27311 r0 *1 116.325,150.15
X$27311 396 625 397 644 645 cell_1rw
* cell instance $27312 m0 *1 116.325,152.88
X$27312 396 626 397 644 645 cell_1rw
* cell instance $27313 r0 *1 116.325,152.88
X$27313 396 627 397 644 645 cell_1rw
* cell instance $27314 m0 *1 116.325,155.61
X$27314 396 628 397 644 645 cell_1rw
* cell instance $27315 r0 *1 116.325,155.61
X$27315 396 629 397 644 645 cell_1rw
* cell instance $27316 m0 *1 116.325,158.34
X$27316 396 630 397 644 645 cell_1rw
* cell instance $27317 r0 *1 116.325,158.34
X$27317 396 631 397 644 645 cell_1rw
* cell instance $27318 m0 *1 116.325,161.07
X$27318 396 632 397 644 645 cell_1rw
* cell instance $27319 r0 *1 116.325,161.07
X$27319 396 633 397 644 645 cell_1rw
* cell instance $27320 m0 *1 116.325,163.8
X$27320 396 634 397 644 645 cell_1rw
* cell instance $27321 r0 *1 116.325,163.8
X$27321 396 635 397 644 645 cell_1rw
* cell instance $27322 m0 *1 116.325,166.53
X$27322 396 637 397 644 645 cell_1rw
* cell instance $27323 r0 *1 116.325,166.53
X$27323 396 636 397 644 645 cell_1rw
* cell instance $27324 m0 *1 116.325,169.26
X$27324 396 639 397 644 645 cell_1rw
* cell instance $27325 r0 *1 116.325,169.26
X$27325 396 638 397 644 645 cell_1rw
* cell instance $27326 m0 *1 116.325,171.99
X$27326 396 640 397 644 645 cell_1rw
* cell instance $27327 r0 *1 116.325,171.99
X$27327 396 641 397 644 645 cell_1rw
* cell instance $27328 m0 *1 116.325,174.72
X$27328 396 642 397 644 645 cell_1rw
* cell instance $27329 r0 *1 116.325,174.72
X$27329 396 643 397 644 645 cell_1rw
* cell instance $27330 m0 *1 117.03,90.09
X$27330 398 581 399 644 645 cell_1rw
* cell instance $27331 r0 *1 117.03,90.09
X$27331 398 580 399 644 645 cell_1rw
* cell instance $27332 m0 *1 117.03,92.82
X$27332 398 583 399 644 645 cell_1rw
* cell instance $27333 r0 *1 117.03,92.82
X$27333 398 582 399 644 645 cell_1rw
* cell instance $27334 m0 *1 117.03,95.55
X$27334 398 584 399 644 645 cell_1rw
* cell instance $27335 m0 *1 117.03,98.28
X$27335 398 586 399 644 645 cell_1rw
* cell instance $27336 r0 *1 117.03,95.55
X$27336 398 585 399 644 645 cell_1rw
* cell instance $27337 m0 *1 117.03,101.01
X$27337 398 588 399 644 645 cell_1rw
* cell instance $27338 r0 *1 117.03,98.28
X$27338 398 587 399 644 645 cell_1rw
* cell instance $27339 r0 *1 117.03,101.01
X$27339 398 589 399 644 645 cell_1rw
* cell instance $27340 m0 *1 117.03,103.74
X$27340 398 590 399 644 645 cell_1rw
* cell instance $27341 r0 *1 117.03,103.74
X$27341 398 591 399 644 645 cell_1rw
* cell instance $27342 m0 *1 117.03,106.47
X$27342 398 593 399 644 645 cell_1rw
* cell instance $27343 r0 *1 117.03,106.47
X$27343 398 592 399 644 645 cell_1rw
* cell instance $27344 m0 *1 117.03,109.2
X$27344 398 594 399 644 645 cell_1rw
* cell instance $27345 r0 *1 117.03,109.2
X$27345 398 595 399 644 645 cell_1rw
* cell instance $27346 m0 *1 117.03,111.93
X$27346 398 597 399 644 645 cell_1rw
* cell instance $27347 r0 *1 117.03,111.93
X$27347 398 596 399 644 645 cell_1rw
* cell instance $27348 m0 *1 117.03,114.66
X$27348 398 598 399 644 645 cell_1rw
* cell instance $27349 r0 *1 117.03,114.66
X$27349 398 599 399 644 645 cell_1rw
* cell instance $27350 m0 *1 117.03,117.39
X$27350 398 600 399 644 645 cell_1rw
* cell instance $27351 r0 *1 117.03,117.39
X$27351 398 601 399 644 645 cell_1rw
* cell instance $27352 m0 *1 117.03,120.12
X$27352 398 602 399 644 645 cell_1rw
* cell instance $27353 r0 *1 117.03,120.12
X$27353 398 603 399 644 645 cell_1rw
* cell instance $27354 m0 *1 117.03,122.85
X$27354 398 604 399 644 645 cell_1rw
* cell instance $27355 r0 *1 117.03,122.85
X$27355 398 605 399 644 645 cell_1rw
* cell instance $27356 m0 *1 117.03,125.58
X$27356 398 606 399 644 645 cell_1rw
* cell instance $27357 r0 *1 117.03,125.58
X$27357 398 607 399 644 645 cell_1rw
* cell instance $27358 m0 *1 117.03,128.31
X$27358 398 609 399 644 645 cell_1rw
* cell instance $27359 r0 *1 117.03,128.31
X$27359 398 608 399 644 645 cell_1rw
* cell instance $27360 m0 *1 117.03,131.04
X$27360 398 610 399 644 645 cell_1rw
* cell instance $27361 r0 *1 117.03,131.04
X$27361 398 611 399 644 645 cell_1rw
* cell instance $27362 m0 *1 117.03,133.77
X$27362 398 612 399 644 645 cell_1rw
* cell instance $27363 m0 *1 117.03,136.5
X$27363 398 615 399 644 645 cell_1rw
* cell instance $27364 r0 *1 117.03,133.77
X$27364 398 613 399 644 645 cell_1rw
* cell instance $27365 m0 *1 117.03,139.23
X$27365 398 617 399 644 645 cell_1rw
* cell instance $27366 r0 *1 117.03,136.5
X$27366 398 614 399 644 645 cell_1rw
* cell instance $27367 r0 *1 117.03,139.23
X$27367 398 616 399 644 645 cell_1rw
* cell instance $27368 m0 *1 117.03,141.96
X$27368 398 618 399 644 645 cell_1rw
* cell instance $27369 r0 *1 117.03,141.96
X$27369 398 619 399 644 645 cell_1rw
* cell instance $27370 m0 *1 117.03,144.69
X$27370 398 620 399 644 645 cell_1rw
* cell instance $27371 r0 *1 117.03,144.69
X$27371 398 621 399 644 645 cell_1rw
* cell instance $27372 m0 *1 117.03,147.42
X$27372 398 622 399 644 645 cell_1rw
* cell instance $27373 r0 *1 117.03,147.42
X$27373 398 623 399 644 645 cell_1rw
* cell instance $27374 m0 *1 117.03,150.15
X$27374 398 624 399 644 645 cell_1rw
* cell instance $27375 r0 *1 117.03,150.15
X$27375 398 625 399 644 645 cell_1rw
* cell instance $27376 m0 *1 117.03,152.88
X$27376 398 626 399 644 645 cell_1rw
* cell instance $27377 m0 *1 117.03,155.61
X$27377 398 628 399 644 645 cell_1rw
* cell instance $27378 r0 *1 117.03,152.88
X$27378 398 627 399 644 645 cell_1rw
* cell instance $27379 r0 *1 117.03,155.61
X$27379 398 629 399 644 645 cell_1rw
* cell instance $27380 m0 *1 117.03,158.34
X$27380 398 630 399 644 645 cell_1rw
* cell instance $27381 r0 *1 117.03,158.34
X$27381 398 631 399 644 645 cell_1rw
* cell instance $27382 m0 *1 117.03,161.07
X$27382 398 632 399 644 645 cell_1rw
* cell instance $27383 r0 *1 117.03,161.07
X$27383 398 633 399 644 645 cell_1rw
* cell instance $27384 m0 *1 117.03,163.8
X$27384 398 634 399 644 645 cell_1rw
* cell instance $27385 r0 *1 117.03,163.8
X$27385 398 635 399 644 645 cell_1rw
* cell instance $27386 m0 *1 117.03,166.53
X$27386 398 637 399 644 645 cell_1rw
* cell instance $27387 r0 *1 117.03,166.53
X$27387 398 636 399 644 645 cell_1rw
* cell instance $27388 m0 *1 117.03,169.26
X$27388 398 639 399 644 645 cell_1rw
* cell instance $27389 r0 *1 117.03,169.26
X$27389 398 638 399 644 645 cell_1rw
* cell instance $27390 m0 *1 117.03,171.99
X$27390 398 640 399 644 645 cell_1rw
* cell instance $27391 r0 *1 117.03,171.99
X$27391 398 641 399 644 645 cell_1rw
* cell instance $27392 m0 *1 117.03,174.72
X$27392 398 642 399 644 645 cell_1rw
* cell instance $27393 r0 *1 117.03,174.72
X$27393 398 643 399 644 645 cell_1rw
* cell instance $27394 m0 *1 117.735,90.09
X$27394 400 581 401 644 645 cell_1rw
* cell instance $27395 r0 *1 117.735,90.09
X$27395 400 580 401 644 645 cell_1rw
* cell instance $27396 m0 *1 117.735,92.82
X$27396 400 583 401 644 645 cell_1rw
* cell instance $27397 m0 *1 117.735,95.55
X$27397 400 584 401 644 645 cell_1rw
* cell instance $27398 r0 *1 117.735,92.82
X$27398 400 582 401 644 645 cell_1rw
* cell instance $27399 r0 *1 117.735,95.55
X$27399 400 585 401 644 645 cell_1rw
* cell instance $27400 m0 *1 117.735,98.28
X$27400 400 586 401 644 645 cell_1rw
* cell instance $27401 m0 *1 117.735,101.01
X$27401 400 588 401 644 645 cell_1rw
* cell instance $27402 r0 *1 117.735,98.28
X$27402 400 587 401 644 645 cell_1rw
* cell instance $27403 m0 *1 117.735,103.74
X$27403 400 590 401 644 645 cell_1rw
* cell instance $27404 r0 *1 117.735,101.01
X$27404 400 589 401 644 645 cell_1rw
* cell instance $27405 r0 *1 117.735,103.74
X$27405 400 591 401 644 645 cell_1rw
* cell instance $27406 m0 *1 117.735,106.47
X$27406 400 593 401 644 645 cell_1rw
* cell instance $27407 m0 *1 117.735,109.2
X$27407 400 594 401 644 645 cell_1rw
* cell instance $27408 r0 *1 117.735,106.47
X$27408 400 592 401 644 645 cell_1rw
* cell instance $27409 m0 *1 117.735,111.93
X$27409 400 597 401 644 645 cell_1rw
* cell instance $27410 r0 *1 117.735,109.2
X$27410 400 595 401 644 645 cell_1rw
* cell instance $27411 r0 *1 117.735,111.93
X$27411 400 596 401 644 645 cell_1rw
* cell instance $27412 m0 *1 117.735,114.66
X$27412 400 598 401 644 645 cell_1rw
* cell instance $27413 r0 *1 117.735,114.66
X$27413 400 599 401 644 645 cell_1rw
* cell instance $27414 m0 *1 117.735,117.39
X$27414 400 600 401 644 645 cell_1rw
* cell instance $27415 m0 *1 117.735,120.12
X$27415 400 602 401 644 645 cell_1rw
* cell instance $27416 r0 *1 117.735,117.39
X$27416 400 601 401 644 645 cell_1rw
* cell instance $27417 r0 *1 117.735,120.12
X$27417 400 603 401 644 645 cell_1rw
* cell instance $27418 m0 *1 117.735,122.85
X$27418 400 604 401 644 645 cell_1rw
* cell instance $27419 r0 *1 117.735,122.85
X$27419 400 605 401 644 645 cell_1rw
* cell instance $27420 m0 *1 117.735,125.58
X$27420 400 606 401 644 645 cell_1rw
* cell instance $27421 r0 *1 117.735,125.58
X$27421 400 607 401 644 645 cell_1rw
* cell instance $27422 m0 *1 117.735,128.31
X$27422 400 609 401 644 645 cell_1rw
* cell instance $27423 r0 *1 117.735,128.31
X$27423 400 608 401 644 645 cell_1rw
* cell instance $27424 m0 *1 117.735,131.04
X$27424 400 610 401 644 645 cell_1rw
* cell instance $27425 r0 *1 117.735,131.04
X$27425 400 611 401 644 645 cell_1rw
* cell instance $27426 m0 *1 117.735,133.77
X$27426 400 612 401 644 645 cell_1rw
* cell instance $27427 m0 *1 117.735,136.5
X$27427 400 615 401 644 645 cell_1rw
* cell instance $27428 r0 *1 117.735,133.77
X$27428 400 613 401 644 645 cell_1rw
* cell instance $27429 r0 *1 117.735,136.5
X$27429 400 614 401 644 645 cell_1rw
* cell instance $27430 m0 *1 117.735,139.23
X$27430 400 617 401 644 645 cell_1rw
* cell instance $27431 r0 *1 117.735,139.23
X$27431 400 616 401 644 645 cell_1rw
* cell instance $27432 m0 *1 117.735,141.96
X$27432 400 618 401 644 645 cell_1rw
* cell instance $27433 m0 *1 117.735,144.69
X$27433 400 620 401 644 645 cell_1rw
* cell instance $27434 r0 *1 117.735,141.96
X$27434 400 619 401 644 645 cell_1rw
* cell instance $27435 r0 *1 117.735,144.69
X$27435 400 621 401 644 645 cell_1rw
* cell instance $27436 m0 *1 117.735,147.42
X$27436 400 622 401 644 645 cell_1rw
* cell instance $27437 m0 *1 117.735,150.15
X$27437 400 624 401 644 645 cell_1rw
* cell instance $27438 r0 *1 117.735,147.42
X$27438 400 623 401 644 645 cell_1rw
* cell instance $27439 r0 *1 117.735,150.15
X$27439 400 625 401 644 645 cell_1rw
* cell instance $27440 m0 *1 117.735,152.88
X$27440 400 626 401 644 645 cell_1rw
* cell instance $27441 m0 *1 117.735,155.61
X$27441 400 628 401 644 645 cell_1rw
* cell instance $27442 r0 *1 117.735,152.88
X$27442 400 627 401 644 645 cell_1rw
* cell instance $27443 r0 *1 117.735,155.61
X$27443 400 629 401 644 645 cell_1rw
* cell instance $27444 m0 *1 117.735,158.34
X$27444 400 630 401 644 645 cell_1rw
* cell instance $27445 r0 *1 117.735,158.34
X$27445 400 631 401 644 645 cell_1rw
* cell instance $27446 m0 *1 117.735,161.07
X$27446 400 632 401 644 645 cell_1rw
* cell instance $27447 r0 *1 117.735,161.07
X$27447 400 633 401 644 645 cell_1rw
* cell instance $27448 m0 *1 117.735,163.8
X$27448 400 634 401 644 645 cell_1rw
* cell instance $27449 r0 *1 117.735,163.8
X$27449 400 635 401 644 645 cell_1rw
* cell instance $27450 m0 *1 117.735,166.53
X$27450 400 637 401 644 645 cell_1rw
* cell instance $27451 r0 *1 117.735,166.53
X$27451 400 636 401 644 645 cell_1rw
* cell instance $27452 m0 *1 117.735,169.26
X$27452 400 639 401 644 645 cell_1rw
* cell instance $27453 r0 *1 117.735,169.26
X$27453 400 638 401 644 645 cell_1rw
* cell instance $27454 m0 *1 117.735,171.99
X$27454 400 640 401 644 645 cell_1rw
* cell instance $27455 r0 *1 117.735,171.99
X$27455 400 641 401 644 645 cell_1rw
* cell instance $27456 m0 *1 117.735,174.72
X$27456 400 642 401 644 645 cell_1rw
* cell instance $27457 r0 *1 117.735,174.72
X$27457 400 643 401 644 645 cell_1rw
* cell instance $27458 m0 *1 118.44,90.09
X$27458 402 581 403 644 645 cell_1rw
* cell instance $27459 r0 *1 118.44,90.09
X$27459 402 580 403 644 645 cell_1rw
* cell instance $27460 m0 *1 118.44,92.82
X$27460 402 583 403 644 645 cell_1rw
* cell instance $27461 r0 *1 118.44,92.82
X$27461 402 582 403 644 645 cell_1rw
* cell instance $27462 m0 *1 118.44,95.55
X$27462 402 584 403 644 645 cell_1rw
* cell instance $27463 r0 *1 118.44,95.55
X$27463 402 585 403 644 645 cell_1rw
* cell instance $27464 m0 *1 118.44,98.28
X$27464 402 586 403 644 645 cell_1rw
* cell instance $27465 r0 *1 118.44,98.28
X$27465 402 587 403 644 645 cell_1rw
* cell instance $27466 m0 *1 118.44,101.01
X$27466 402 588 403 644 645 cell_1rw
* cell instance $27467 r0 *1 118.44,101.01
X$27467 402 589 403 644 645 cell_1rw
* cell instance $27468 m0 *1 118.44,103.74
X$27468 402 590 403 644 645 cell_1rw
* cell instance $27469 r0 *1 118.44,103.74
X$27469 402 591 403 644 645 cell_1rw
* cell instance $27470 m0 *1 118.44,106.47
X$27470 402 593 403 644 645 cell_1rw
* cell instance $27471 m0 *1 118.44,109.2
X$27471 402 594 403 644 645 cell_1rw
* cell instance $27472 r0 *1 118.44,106.47
X$27472 402 592 403 644 645 cell_1rw
* cell instance $27473 m0 *1 118.44,111.93
X$27473 402 597 403 644 645 cell_1rw
* cell instance $27474 r0 *1 118.44,109.2
X$27474 402 595 403 644 645 cell_1rw
* cell instance $27475 r0 *1 118.44,111.93
X$27475 402 596 403 644 645 cell_1rw
* cell instance $27476 m0 *1 118.44,114.66
X$27476 402 598 403 644 645 cell_1rw
* cell instance $27477 r0 *1 118.44,114.66
X$27477 402 599 403 644 645 cell_1rw
* cell instance $27478 m0 *1 118.44,117.39
X$27478 402 600 403 644 645 cell_1rw
* cell instance $27479 r0 *1 118.44,117.39
X$27479 402 601 403 644 645 cell_1rw
* cell instance $27480 m0 *1 118.44,120.12
X$27480 402 602 403 644 645 cell_1rw
* cell instance $27481 r0 *1 118.44,120.12
X$27481 402 603 403 644 645 cell_1rw
* cell instance $27482 m0 *1 118.44,122.85
X$27482 402 604 403 644 645 cell_1rw
* cell instance $27483 r0 *1 118.44,122.85
X$27483 402 605 403 644 645 cell_1rw
* cell instance $27484 m0 *1 118.44,125.58
X$27484 402 606 403 644 645 cell_1rw
* cell instance $27485 r0 *1 118.44,125.58
X$27485 402 607 403 644 645 cell_1rw
* cell instance $27486 m0 *1 118.44,128.31
X$27486 402 609 403 644 645 cell_1rw
* cell instance $27487 r0 *1 118.44,128.31
X$27487 402 608 403 644 645 cell_1rw
* cell instance $27488 m0 *1 118.44,131.04
X$27488 402 610 403 644 645 cell_1rw
* cell instance $27489 r0 *1 118.44,131.04
X$27489 402 611 403 644 645 cell_1rw
* cell instance $27490 m0 *1 118.44,133.77
X$27490 402 612 403 644 645 cell_1rw
* cell instance $27491 m0 *1 118.44,136.5
X$27491 402 615 403 644 645 cell_1rw
* cell instance $27492 r0 *1 118.44,133.77
X$27492 402 613 403 644 645 cell_1rw
* cell instance $27493 r0 *1 118.44,136.5
X$27493 402 614 403 644 645 cell_1rw
* cell instance $27494 m0 *1 118.44,139.23
X$27494 402 617 403 644 645 cell_1rw
* cell instance $27495 m0 *1 118.44,141.96
X$27495 402 618 403 644 645 cell_1rw
* cell instance $27496 r0 *1 118.44,139.23
X$27496 402 616 403 644 645 cell_1rw
* cell instance $27497 m0 *1 118.44,144.69
X$27497 402 620 403 644 645 cell_1rw
* cell instance $27498 r0 *1 118.44,141.96
X$27498 402 619 403 644 645 cell_1rw
* cell instance $27499 r0 *1 118.44,144.69
X$27499 402 621 403 644 645 cell_1rw
* cell instance $27500 m0 *1 118.44,147.42
X$27500 402 622 403 644 645 cell_1rw
* cell instance $27501 r0 *1 118.44,147.42
X$27501 402 623 403 644 645 cell_1rw
* cell instance $27502 m0 *1 118.44,150.15
X$27502 402 624 403 644 645 cell_1rw
* cell instance $27503 r0 *1 118.44,150.15
X$27503 402 625 403 644 645 cell_1rw
* cell instance $27504 m0 *1 118.44,152.88
X$27504 402 626 403 644 645 cell_1rw
* cell instance $27505 r0 *1 118.44,152.88
X$27505 402 627 403 644 645 cell_1rw
* cell instance $27506 m0 *1 118.44,155.61
X$27506 402 628 403 644 645 cell_1rw
* cell instance $27507 r0 *1 118.44,155.61
X$27507 402 629 403 644 645 cell_1rw
* cell instance $27508 m0 *1 118.44,158.34
X$27508 402 630 403 644 645 cell_1rw
* cell instance $27509 m0 *1 118.44,161.07
X$27509 402 632 403 644 645 cell_1rw
* cell instance $27510 r0 *1 118.44,158.34
X$27510 402 631 403 644 645 cell_1rw
* cell instance $27511 r0 *1 118.44,161.07
X$27511 402 633 403 644 645 cell_1rw
* cell instance $27512 m0 *1 118.44,163.8
X$27512 402 634 403 644 645 cell_1rw
* cell instance $27513 r0 *1 118.44,163.8
X$27513 402 635 403 644 645 cell_1rw
* cell instance $27514 m0 *1 118.44,166.53
X$27514 402 637 403 644 645 cell_1rw
* cell instance $27515 r0 *1 118.44,166.53
X$27515 402 636 403 644 645 cell_1rw
* cell instance $27516 m0 *1 118.44,169.26
X$27516 402 639 403 644 645 cell_1rw
* cell instance $27517 r0 *1 118.44,169.26
X$27517 402 638 403 644 645 cell_1rw
* cell instance $27518 m0 *1 118.44,171.99
X$27518 402 640 403 644 645 cell_1rw
* cell instance $27519 r0 *1 118.44,171.99
X$27519 402 641 403 644 645 cell_1rw
* cell instance $27520 m0 *1 118.44,174.72
X$27520 402 642 403 644 645 cell_1rw
* cell instance $27521 r0 *1 118.44,174.72
X$27521 402 643 403 644 645 cell_1rw
* cell instance $27522 m0 *1 119.145,90.09
X$27522 404 581 405 644 645 cell_1rw
* cell instance $27523 r0 *1 119.145,90.09
X$27523 404 580 405 644 645 cell_1rw
* cell instance $27524 m0 *1 119.145,92.82
X$27524 404 583 405 644 645 cell_1rw
* cell instance $27525 r0 *1 119.145,92.82
X$27525 404 582 405 644 645 cell_1rw
* cell instance $27526 m0 *1 119.145,95.55
X$27526 404 584 405 644 645 cell_1rw
* cell instance $27527 r0 *1 119.145,95.55
X$27527 404 585 405 644 645 cell_1rw
* cell instance $27528 m0 *1 119.145,98.28
X$27528 404 586 405 644 645 cell_1rw
* cell instance $27529 r0 *1 119.145,98.28
X$27529 404 587 405 644 645 cell_1rw
* cell instance $27530 m0 *1 119.145,101.01
X$27530 404 588 405 644 645 cell_1rw
* cell instance $27531 r0 *1 119.145,101.01
X$27531 404 589 405 644 645 cell_1rw
* cell instance $27532 m0 *1 119.145,103.74
X$27532 404 590 405 644 645 cell_1rw
* cell instance $27533 m0 *1 119.145,106.47
X$27533 404 593 405 644 645 cell_1rw
* cell instance $27534 r0 *1 119.145,103.74
X$27534 404 591 405 644 645 cell_1rw
* cell instance $27535 r0 *1 119.145,106.47
X$27535 404 592 405 644 645 cell_1rw
* cell instance $27536 m0 *1 119.145,109.2
X$27536 404 594 405 644 645 cell_1rw
* cell instance $27537 m0 *1 119.145,111.93
X$27537 404 597 405 644 645 cell_1rw
* cell instance $27538 r0 *1 119.145,109.2
X$27538 404 595 405 644 645 cell_1rw
* cell instance $27539 r0 *1 119.145,111.93
X$27539 404 596 405 644 645 cell_1rw
* cell instance $27540 m0 *1 119.145,114.66
X$27540 404 598 405 644 645 cell_1rw
* cell instance $27541 r0 *1 119.145,114.66
X$27541 404 599 405 644 645 cell_1rw
* cell instance $27542 m0 *1 119.145,117.39
X$27542 404 600 405 644 645 cell_1rw
* cell instance $27543 r0 *1 119.145,117.39
X$27543 404 601 405 644 645 cell_1rw
* cell instance $27544 m0 *1 119.145,120.12
X$27544 404 602 405 644 645 cell_1rw
* cell instance $27545 r0 *1 119.145,120.12
X$27545 404 603 405 644 645 cell_1rw
* cell instance $27546 m0 *1 119.145,122.85
X$27546 404 604 405 644 645 cell_1rw
* cell instance $27547 r0 *1 119.145,122.85
X$27547 404 605 405 644 645 cell_1rw
* cell instance $27548 m0 *1 119.145,125.58
X$27548 404 606 405 644 645 cell_1rw
* cell instance $27549 r0 *1 119.145,125.58
X$27549 404 607 405 644 645 cell_1rw
* cell instance $27550 m0 *1 119.145,128.31
X$27550 404 609 405 644 645 cell_1rw
* cell instance $27551 r0 *1 119.145,128.31
X$27551 404 608 405 644 645 cell_1rw
* cell instance $27552 m0 *1 119.145,131.04
X$27552 404 610 405 644 645 cell_1rw
* cell instance $27553 r0 *1 119.145,131.04
X$27553 404 611 405 644 645 cell_1rw
* cell instance $27554 m0 *1 119.145,133.77
X$27554 404 612 405 644 645 cell_1rw
* cell instance $27555 m0 *1 119.145,136.5
X$27555 404 615 405 644 645 cell_1rw
* cell instance $27556 r0 *1 119.145,133.77
X$27556 404 613 405 644 645 cell_1rw
* cell instance $27557 m0 *1 119.145,139.23
X$27557 404 617 405 644 645 cell_1rw
* cell instance $27558 r0 *1 119.145,136.5
X$27558 404 614 405 644 645 cell_1rw
* cell instance $27559 r0 *1 119.145,139.23
X$27559 404 616 405 644 645 cell_1rw
* cell instance $27560 m0 *1 119.145,141.96
X$27560 404 618 405 644 645 cell_1rw
* cell instance $27561 r0 *1 119.145,141.96
X$27561 404 619 405 644 645 cell_1rw
* cell instance $27562 m0 *1 119.145,144.69
X$27562 404 620 405 644 645 cell_1rw
* cell instance $27563 r0 *1 119.145,144.69
X$27563 404 621 405 644 645 cell_1rw
* cell instance $27564 m0 *1 119.145,147.42
X$27564 404 622 405 644 645 cell_1rw
* cell instance $27565 r0 *1 119.145,147.42
X$27565 404 623 405 644 645 cell_1rw
* cell instance $27566 m0 *1 119.145,150.15
X$27566 404 624 405 644 645 cell_1rw
* cell instance $27567 r0 *1 119.145,150.15
X$27567 404 625 405 644 645 cell_1rw
* cell instance $27568 m0 *1 119.145,152.88
X$27568 404 626 405 644 645 cell_1rw
* cell instance $27569 r0 *1 119.145,152.88
X$27569 404 627 405 644 645 cell_1rw
* cell instance $27570 m0 *1 119.145,155.61
X$27570 404 628 405 644 645 cell_1rw
* cell instance $27571 r0 *1 119.145,155.61
X$27571 404 629 405 644 645 cell_1rw
* cell instance $27572 m0 *1 119.145,158.34
X$27572 404 630 405 644 645 cell_1rw
* cell instance $27573 m0 *1 119.145,161.07
X$27573 404 632 405 644 645 cell_1rw
* cell instance $27574 r0 *1 119.145,158.34
X$27574 404 631 405 644 645 cell_1rw
* cell instance $27575 r0 *1 119.145,161.07
X$27575 404 633 405 644 645 cell_1rw
* cell instance $27576 m0 *1 119.145,163.8
X$27576 404 634 405 644 645 cell_1rw
* cell instance $27577 r0 *1 119.145,163.8
X$27577 404 635 405 644 645 cell_1rw
* cell instance $27578 m0 *1 119.145,166.53
X$27578 404 637 405 644 645 cell_1rw
* cell instance $27579 r0 *1 119.145,166.53
X$27579 404 636 405 644 645 cell_1rw
* cell instance $27580 m0 *1 119.145,169.26
X$27580 404 639 405 644 645 cell_1rw
* cell instance $27581 r0 *1 119.145,169.26
X$27581 404 638 405 644 645 cell_1rw
* cell instance $27582 m0 *1 119.145,171.99
X$27582 404 640 405 644 645 cell_1rw
* cell instance $27583 r0 *1 119.145,171.99
X$27583 404 641 405 644 645 cell_1rw
* cell instance $27584 m0 *1 119.145,174.72
X$27584 404 642 405 644 645 cell_1rw
* cell instance $27585 r0 *1 119.145,174.72
X$27585 404 643 405 644 645 cell_1rw
* cell instance $27586 m0 *1 119.85,90.09
X$27586 406 581 407 644 645 cell_1rw
* cell instance $27587 r0 *1 119.85,90.09
X$27587 406 580 407 644 645 cell_1rw
* cell instance $27588 m0 *1 119.85,92.82
X$27588 406 583 407 644 645 cell_1rw
* cell instance $27589 m0 *1 119.85,95.55
X$27589 406 584 407 644 645 cell_1rw
* cell instance $27590 r0 *1 119.85,92.82
X$27590 406 582 407 644 645 cell_1rw
* cell instance $27591 r0 *1 119.85,95.55
X$27591 406 585 407 644 645 cell_1rw
* cell instance $27592 m0 *1 119.85,98.28
X$27592 406 586 407 644 645 cell_1rw
* cell instance $27593 r0 *1 119.85,98.28
X$27593 406 587 407 644 645 cell_1rw
* cell instance $27594 m0 *1 119.85,101.01
X$27594 406 588 407 644 645 cell_1rw
* cell instance $27595 r0 *1 119.85,101.01
X$27595 406 589 407 644 645 cell_1rw
* cell instance $27596 m0 *1 119.85,103.74
X$27596 406 590 407 644 645 cell_1rw
* cell instance $27597 r0 *1 119.85,103.74
X$27597 406 591 407 644 645 cell_1rw
* cell instance $27598 m0 *1 119.85,106.47
X$27598 406 593 407 644 645 cell_1rw
* cell instance $27599 r0 *1 119.85,106.47
X$27599 406 592 407 644 645 cell_1rw
* cell instance $27600 m0 *1 119.85,109.2
X$27600 406 594 407 644 645 cell_1rw
* cell instance $27601 r0 *1 119.85,109.2
X$27601 406 595 407 644 645 cell_1rw
* cell instance $27602 m0 *1 119.85,111.93
X$27602 406 597 407 644 645 cell_1rw
* cell instance $27603 r0 *1 119.85,111.93
X$27603 406 596 407 644 645 cell_1rw
* cell instance $27604 m0 *1 119.85,114.66
X$27604 406 598 407 644 645 cell_1rw
* cell instance $27605 r0 *1 119.85,114.66
X$27605 406 599 407 644 645 cell_1rw
* cell instance $27606 m0 *1 119.85,117.39
X$27606 406 600 407 644 645 cell_1rw
* cell instance $27607 r0 *1 119.85,117.39
X$27607 406 601 407 644 645 cell_1rw
* cell instance $27608 m0 *1 119.85,120.12
X$27608 406 602 407 644 645 cell_1rw
* cell instance $27609 r0 *1 119.85,120.12
X$27609 406 603 407 644 645 cell_1rw
* cell instance $27610 m0 *1 119.85,122.85
X$27610 406 604 407 644 645 cell_1rw
* cell instance $27611 r0 *1 119.85,122.85
X$27611 406 605 407 644 645 cell_1rw
* cell instance $27612 m0 *1 119.85,125.58
X$27612 406 606 407 644 645 cell_1rw
* cell instance $27613 r0 *1 119.85,125.58
X$27613 406 607 407 644 645 cell_1rw
* cell instance $27614 m0 *1 119.85,128.31
X$27614 406 609 407 644 645 cell_1rw
* cell instance $27615 r0 *1 119.85,128.31
X$27615 406 608 407 644 645 cell_1rw
* cell instance $27616 m0 *1 119.85,131.04
X$27616 406 610 407 644 645 cell_1rw
* cell instance $27617 r0 *1 119.85,131.04
X$27617 406 611 407 644 645 cell_1rw
* cell instance $27618 m0 *1 119.85,133.77
X$27618 406 612 407 644 645 cell_1rw
* cell instance $27619 r0 *1 119.85,133.77
X$27619 406 613 407 644 645 cell_1rw
* cell instance $27620 m0 *1 119.85,136.5
X$27620 406 615 407 644 645 cell_1rw
* cell instance $27621 r0 *1 119.85,136.5
X$27621 406 614 407 644 645 cell_1rw
* cell instance $27622 m0 *1 119.85,139.23
X$27622 406 617 407 644 645 cell_1rw
* cell instance $27623 r0 *1 119.85,139.23
X$27623 406 616 407 644 645 cell_1rw
* cell instance $27624 m0 *1 119.85,141.96
X$27624 406 618 407 644 645 cell_1rw
* cell instance $27625 r0 *1 119.85,141.96
X$27625 406 619 407 644 645 cell_1rw
* cell instance $27626 m0 *1 119.85,144.69
X$27626 406 620 407 644 645 cell_1rw
* cell instance $27627 r0 *1 119.85,144.69
X$27627 406 621 407 644 645 cell_1rw
* cell instance $27628 m0 *1 119.85,147.42
X$27628 406 622 407 644 645 cell_1rw
* cell instance $27629 m0 *1 119.85,150.15
X$27629 406 624 407 644 645 cell_1rw
* cell instance $27630 r0 *1 119.85,147.42
X$27630 406 623 407 644 645 cell_1rw
* cell instance $27631 m0 *1 119.85,152.88
X$27631 406 626 407 644 645 cell_1rw
* cell instance $27632 r0 *1 119.85,150.15
X$27632 406 625 407 644 645 cell_1rw
* cell instance $27633 r0 *1 119.85,152.88
X$27633 406 627 407 644 645 cell_1rw
* cell instance $27634 m0 *1 119.85,155.61
X$27634 406 628 407 644 645 cell_1rw
* cell instance $27635 m0 *1 119.85,158.34
X$27635 406 630 407 644 645 cell_1rw
* cell instance $27636 r0 *1 119.85,155.61
X$27636 406 629 407 644 645 cell_1rw
* cell instance $27637 r0 *1 119.85,158.34
X$27637 406 631 407 644 645 cell_1rw
* cell instance $27638 m0 *1 119.85,161.07
X$27638 406 632 407 644 645 cell_1rw
* cell instance $27639 r0 *1 119.85,161.07
X$27639 406 633 407 644 645 cell_1rw
* cell instance $27640 m0 *1 119.85,163.8
X$27640 406 634 407 644 645 cell_1rw
* cell instance $27641 r0 *1 119.85,163.8
X$27641 406 635 407 644 645 cell_1rw
* cell instance $27642 m0 *1 119.85,166.53
X$27642 406 637 407 644 645 cell_1rw
* cell instance $27643 m0 *1 119.85,169.26
X$27643 406 639 407 644 645 cell_1rw
* cell instance $27644 r0 *1 119.85,166.53
X$27644 406 636 407 644 645 cell_1rw
* cell instance $27645 r0 *1 119.85,169.26
X$27645 406 638 407 644 645 cell_1rw
* cell instance $27646 m0 *1 119.85,171.99
X$27646 406 640 407 644 645 cell_1rw
* cell instance $27647 r0 *1 119.85,171.99
X$27647 406 641 407 644 645 cell_1rw
* cell instance $27648 m0 *1 119.85,174.72
X$27648 406 642 407 644 645 cell_1rw
* cell instance $27649 r0 *1 119.85,174.72
X$27649 406 643 407 644 645 cell_1rw
* cell instance $27650 m0 *1 120.555,90.09
X$27650 408 581 409 644 645 cell_1rw
* cell instance $27651 m0 *1 120.555,92.82
X$27651 408 583 409 644 645 cell_1rw
* cell instance $27652 r0 *1 120.555,90.09
X$27652 408 580 409 644 645 cell_1rw
* cell instance $27653 r0 *1 120.555,92.82
X$27653 408 582 409 644 645 cell_1rw
* cell instance $27654 m0 *1 120.555,95.55
X$27654 408 584 409 644 645 cell_1rw
* cell instance $27655 r0 *1 120.555,95.55
X$27655 408 585 409 644 645 cell_1rw
* cell instance $27656 m0 *1 120.555,98.28
X$27656 408 586 409 644 645 cell_1rw
* cell instance $27657 r0 *1 120.555,98.28
X$27657 408 587 409 644 645 cell_1rw
* cell instance $27658 m0 *1 120.555,101.01
X$27658 408 588 409 644 645 cell_1rw
* cell instance $27659 r0 *1 120.555,101.01
X$27659 408 589 409 644 645 cell_1rw
* cell instance $27660 m0 *1 120.555,103.74
X$27660 408 590 409 644 645 cell_1rw
* cell instance $27661 r0 *1 120.555,103.74
X$27661 408 591 409 644 645 cell_1rw
* cell instance $27662 m0 *1 120.555,106.47
X$27662 408 593 409 644 645 cell_1rw
* cell instance $27663 m0 *1 120.555,109.2
X$27663 408 594 409 644 645 cell_1rw
* cell instance $27664 r0 *1 120.555,106.47
X$27664 408 592 409 644 645 cell_1rw
* cell instance $27665 r0 *1 120.555,109.2
X$27665 408 595 409 644 645 cell_1rw
* cell instance $27666 m0 *1 120.555,111.93
X$27666 408 597 409 644 645 cell_1rw
* cell instance $27667 m0 *1 120.555,114.66
X$27667 408 598 409 644 645 cell_1rw
* cell instance $27668 r0 *1 120.555,111.93
X$27668 408 596 409 644 645 cell_1rw
* cell instance $27669 r0 *1 120.555,114.66
X$27669 408 599 409 644 645 cell_1rw
* cell instance $27670 m0 *1 120.555,117.39
X$27670 408 600 409 644 645 cell_1rw
* cell instance $27671 m0 *1 120.555,120.12
X$27671 408 602 409 644 645 cell_1rw
* cell instance $27672 r0 *1 120.555,117.39
X$27672 408 601 409 644 645 cell_1rw
* cell instance $27673 r0 *1 120.555,120.12
X$27673 408 603 409 644 645 cell_1rw
* cell instance $27674 m0 *1 120.555,122.85
X$27674 408 604 409 644 645 cell_1rw
* cell instance $27675 r0 *1 120.555,122.85
X$27675 408 605 409 644 645 cell_1rw
* cell instance $27676 m0 *1 120.555,125.58
X$27676 408 606 409 644 645 cell_1rw
* cell instance $27677 m0 *1 120.555,128.31
X$27677 408 609 409 644 645 cell_1rw
* cell instance $27678 r0 *1 120.555,125.58
X$27678 408 607 409 644 645 cell_1rw
* cell instance $27679 m0 *1 120.555,131.04
X$27679 408 610 409 644 645 cell_1rw
* cell instance $27680 r0 *1 120.555,128.31
X$27680 408 608 409 644 645 cell_1rw
* cell instance $27681 r0 *1 120.555,131.04
X$27681 408 611 409 644 645 cell_1rw
* cell instance $27682 m0 *1 120.555,133.77
X$27682 408 612 409 644 645 cell_1rw
* cell instance $27683 r0 *1 120.555,133.77
X$27683 408 613 409 644 645 cell_1rw
* cell instance $27684 m0 *1 120.555,136.5
X$27684 408 615 409 644 645 cell_1rw
* cell instance $27685 m0 *1 120.555,139.23
X$27685 408 617 409 644 645 cell_1rw
* cell instance $27686 r0 *1 120.555,136.5
X$27686 408 614 409 644 645 cell_1rw
* cell instance $27687 r0 *1 120.555,139.23
X$27687 408 616 409 644 645 cell_1rw
* cell instance $27688 m0 *1 120.555,141.96
X$27688 408 618 409 644 645 cell_1rw
* cell instance $27689 r0 *1 120.555,141.96
X$27689 408 619 409 644 645 cell_1rw
* cell instance $27690 m0 *1 120.555,144.69
X$27690 408 620 409 644 645 cell_1rw
* cell instance $27691 r0 *1 120.555,144.69
X$27691 408 621 409 644 645 cell_1rw
* cell instance $27692 m0 *1 120.555,147.42
X$27692 408 622 409 644 645 cell_1rw
* cell instance $27693 r0 *1 120.555,147.42
X$27693 408 623 409 644 645 cell_1rw
* cell instance $27694 m0 *1 120.555,150.15
X$27694 408 624 409 644 645 cell_1rw
* cell instance $27695 r0 *1 120.555,150.15
X$27695 408 625 409 644 645 cell_1rw
* cell instance $27696 m0 *1 120.555,152.88
X$27696 408 626 409 644 645 cell_1rw
* cell instance $27697 r0 *1 120.555,152.88
X$27697 408 627 409 644 645 cell_1rw
* cell instance $27698 m0 *1 120.555,155.61
X$27698 408 628 409 644 645 cell_1rw
* cell instance $27699 r0 *1 120.555,155.61
X$27699 408 629 409 644 645 cell_1rw
* cell instance $27700 m0 *1 120.555,158.34
X$27700 408 630 409 644 645 cell_1rw
* cell instance $27701 r0 *1 120.555,158.34
X$27701 408 631 409 644 645 cell_1rw
* cell instance $27702 m0 *1 120.555,161.07
X$27702 408 632 409 644 645 cell_1rw
* cell instance $27703 r0 *1 120.555,161.07
X$27703 408 633 409 644 645 cell_1rw
* cell instance $27704 m0 *1 120.555,163.8
X$27704 408 634 409 644 645 cell_1rw
* cell instance $27705 m0 *1 120.555,166.53
X$27705 408 637 409 644 645 cell_1rw
* cell instance $27706 r0 *1 120.555,163.8
X$27706 408 635 409 644 645 cell_1rw
* cell instance $27707 r0 *1 120.555,166.53
X$27707 408 636 409 644 645 cell_1rw
* cell instance $27708 m0 *1 120.555,169.26
X$27708 408 639 409 644 645 cell_1rw
* cell instance $27709 m0 *1 120.555,171.99
X$27709 408 640 409 644 645 cell_1rw
* cell instance $27710 r0 *1 120.555,169.26
X$27710 408 638 409 644 645 cell_1rw
* cell instance $27711 r0 *1 120.555,171.99
X$27711 408 641 409 644 645 cell_1rw
* cell instance $27712 m0 *1 120.555,174.72
X$27712 408 642 409 644 645 cell_1rw
* cell instance $27713 r0 *1 120.555,174.72
X$27713 408 643 409 644 645 cell_1rw
* cell instance $27714 m0 *1 121.26,90.09
X$27714 410 581 411 644 645 cell_1rw
* cell instance $27715 r0 *1 121.26,90.09
X$27715 410 580 411 644 645 cell_1rw
* cell instance $27716 m0 *1 121.26,92.82
X$27716 410 583 411 644 645 cell_1rw
* cell instance $27717 r0 *1 121.26,92.82
X$27717 410 582 411 644 645 cell_1rw
* cell instance $27718 m0 *1 121.26,95.55
X$27718 410 584 411 644 645 cell_1rw
* cell instance $27719 r0 *1 121.26,95.55
X$27719 410 585 411 644 645 cell_1rw
* cell instance $27720 m0 *1 121.26,98.28
X$27720 410 586 411 644 645 cell_1rw
* cell instance $27721 r0 *1 121.26,98.28
X$27721 410 587 411 644 645 cell_1rw
* cell instance $27722 m0 *1 121.26,101.01
X$27722 410 588 411 644 645 cell_1rw
* cell instance $27723 r0 *1 121.26,101.01
X$27723 410 589 411 644 645 cell_1rw
* cell instance $27724 m0 *1 121.26,103.74
X$27724 410 590 411 644 645 cell_1rw
* cell instance $27725 r0 *1 121.26,103.74
X$27725 410 591 411 644 645 cell_1rw
* cell instance $27726 m0 *1 121.26,106.47
X$27726 410 593 411 644 645 cell_1rw
* cell instance $27727 m0 *1 121.26,109.2
X$27727 410 594 411 644 645 cell_1rw
* cell instance $27728 r0 *1 121.26,106.47
X$27728 410 592 411 644 645 cell_1rw
* cell instance $27729 r0 *1 121.26,109.2
X$27729 410 595 411 644 645 cell_1rw
* cell instance $27730 m0 *1 121.26,111.93
X$27730 410 597 411 644 645 cell_1rw
* cell instance $27731 r0 *1 121.26,111.93
X$27731 410 596 411 644 645 cell_1rw
* cell instance $27732 m0 *1 121.26,114.66
X$27732 410 598 411 644 645 cell_1rw
* cell instance $27733 r0 *1 121.26,114.66
X$27733 410 599 411 644 645 cell_1rw
* cell instance $27734 m0 *1 121.26,117.39
X$27734 410 600 411 644 645 cell_1rw
* cell instance $27735 r0 *1 121.26,117.39
X$27735 410 601 411 644 645 cell_1rw
* cell instance $27736 m0 *1 121.26,120.12
X$27736 410 602 411 644 645 cell_1rw
* cell instance $27737 r0 *1 121.26,120.12
X$27737 410 603 411 644 645 cell_1rw
* cell instance $27738 m0 *1 121.26,122.85
X$27738 410 604 411 644 645 cell_1rw
* cell instance $27739 r0 *1 121.26,122.85
X$27739 410 605 411 644 645 cell_1rw
* cell instance $27740 m0 *1 121.26,125.58
X$27740 410 606 411 644 645 cell_1rw
* cell instance $27741 r0 *1 121.26,125.58
X$27741 410 607 411 644 645 cell_1rw
* cell instance $27742 m0 *1 121.26,128.31
X$27742 410 609 411 644 645 cell_1rw
* cell instance $27743 r0 *1 121.26,128.31
X$27743 410 608 411 644 645 cell_1rw
* cell instance $27744 m0 *1 121.26,131.04
X$27744 410 610 411 644 645 cell_1rw
* cell instance $27745 r0 *1 121.26,131.04
X$27745 410 611 411 644 645 cell_1rw
* cell instance $27746 m0 *1 121.26,133.77
X$27746 410 612 411 644 645 cell_1rw
* cell instance $27747 r0 *1 121.26,133.77
X$27747 410 613 411 644 645 cell_1rw
* cell instance $27748 m0 *1 121.26,136.5
X$27748 410 615 411 644 645 cell_1rw
* cell instance $27749 m0 *1 121.26,139.23
X$27749 410 617 411 644 645 cell_1rw
* cell instance $27750 r0 *1 121.26,136.5
X$27750 410 614 411 644 645 cell_1rw
* cell instance $27751 r0 *1 121.26,139.23
X$27751 410 616 411 644 645 cell_1rw
* cell instance $27752 m0 *1 121.26,141.96
X$27752 410 618 411 644 645 cell_1rw
* cell instance $27753 r0 *1 121.26,141.96
X$27753 410 619 411 644 645 cell_1rw
* cell instance $27754 m0 *1 121.26,144.69
X$27754 410 620 411 644 645 cell_1rw
* cell instance $27755 r0 *1 121.26,144.69
X$27755 410 621 411 644 645 cell_1rw
* cell instance $27756 m0 *1 121.26,147.42
X$27756 410 622 411 644 645 cell_1rw
* cell instance $27757 m0 *1 121.26,150.15
X$27757 410 624 411 644 645 cell_1rw
* cell instance $27758 r0 *1 121.26,147.42
X$27758 410 623 411 644 645 cell_1rw
* cell instance $27759 m0 *1 121.26,152.88
X$27759 410 626 411 644 645 cell_1rw
* cell instance $27760 r0 *1 121.26,150.15
X$27760 410 625 411 644 645 cell_1rw
* cell instance $27761 r0 *1 121.26,152.88
X$27761 410 627 411 644 645 cell_1rw
* cell instance $27762 m0 *1 121.26,155.61
X$27762 410 628 411 644 645 cell_1rw
* cell instance $27763 r0 *1 121.26,155.61
X$27763 410 629 411 644 645 cell_1rw
* cell instance $27764 m0 *1 121.26,158.34
X$27764 410 630 411 644 645 cell_1rw
* cell instance $27765 r0 *1 121.26,158.34
X$27765 410 631 411 644 645 cell_1rw
* cell instance $27766 m0 *1 121.26,161.07
X$27766 410 632 411 644 645 cell_1rw
* cell instance $27767 r0 *1 121.26,161.07
X$27767 410 633 411 644 645 cell_1rw
* cell instance $27768 m0 *1 121.26,163.8
X$27768 410 634 411 644 645 cell_1rw
* cell instance $27769 r0 *1 121.26,163.8
X$27769 410 635 411 644 645 cell_1rw
* cell instance $27770 m0 *1 121.26,166.53
X$27770 410 637 411 644 645 cell_1rw
* cell instance $27771 r0 *1 121.26,166.53
X$27771 410 636 411 644 645 cell_1rw
* cell instance $27772 m0 *1 121.26,169.26
X$27772 410 639 411 644 645 cell_1rw
* cell instance $27773 m0 *1 121.26,171.99
X$27773 410 640 411 644 645 cell_1rw
* cell instance $27774 r0 *1 121.26,169.26
X$27774 410 638 411 644 645 cell_1rw
* cell instance $27775 r0 *1 121.26,171.99
X$27775 410 641 411 644 645 cell_1rw
* cell instance $27776 m0 *1 121.26,174.72
X$27776 410 642 411 644 645 cell_1rw
* cell instance $27777 r0 *1 121.26,174.72
X$27777 410 643 411 644 645 cell_1rw
* cell instance $27778 m0 *1 121.965,90.09
X$27778 412 581 413 644 645 cell_1rw
* cell instance $27779 r0 *1 121.965,90.09
X$27779 412 580 413 644 645 cell_1rw
* cell instance $27780 m0 *1 121.965,92.82
X$27780 412 583 413 644 645 cell_1rw
* cell instance $27781 r0 *1 121.965,92.82
X$27781 412 582 413 644 645 cell_1rw
* cell instance $27782 m0 *1 121.965,95.55
X$27782 412 584 413 644 645 cell_1rw
* cell instance $27783 m0 *1 121.965,98.28
X$27783 412 586 413 644 645 cell_1rw
* cell instance $27784 r0 *1 121.965,95.55
X$27784 412 585 413 644 645 cell_1rw
* cell instance $27785 r0 *1 121.965,98.28
X$27785 412 587 413 644 645 cell_1rw
* cell instance $27786 m0 *1 121.965,101.01
X$27786 412 588 413 644 645 cell_1rw
* cell instance $27787 r0 *1 121.965,101.01
X$27787 412 589 413 644 645 cell_1rw
* cell instance $27788 m0 *1 121.965,103.74
X$27788 412 590 413 644 645 cell_1rw
* cell instance $27789 r0 *1 121.965,103.74
X$27789 412 591 413 644 645 cell_1rw
* cell instance $27790 m0 *1 121.965,106.47
X$27790 412 593 413 644 645 cell_1rw
* cell instance $27791 r0 *1 121.965,106.47
X$27791 412 592 413 644 645 cell_1rw
* cell instance $27792 m0 *1 121.965,109.2
X$27792 412 594 413 644 645 cell_1rw
* cell instance $27793 r0 *1 121.965,109.2
X$27793 412 595 413 644 645 cell_1rw
* cell instance $27794 m0 *1 121.965,111.93
X$27794 412 597 413 644 645 cell_1rw
* cell instance $27795 r0 *1 121.965,111.93
X$27795 412 596 413 644 645 cell_1rw
* cell instance $27796 m0 *1 121.965,114.66
X$27796 412 598 413 644 645 cell_1rw
* cell instance $27797 r0 *1 121.965,114.66
X$27797 412 599 413 644 645 cell_1rw
* cell instance $27798 m0 *1 121.965,117.39
X$27798 412 600 413 644 645 cell_1rw
* cell instance $27799 m0 *1 121.965,120.12
X$27799 412 602 413 644 645 cell_1rw
* cell instance $27800 r0 *1 121.965,117.39
X$27800 412 601 413 644 645 cell_1rw
* cell instance $27801 r0 *1 121.965,120.12
X$27801 412 603 413 644 645 cell_1rw
* cell instance $27802 m0 *1 121.965,122.85
X$27802 412 604 413 644 645 cell_1rw
* cell instance $27803 r0 *1 121.965,122.85
X$27803 412 605 413 644 645 cell_1rw
* cell instance $27804 m0 *1 121.965,125.58
X$27804 412 606 413 644 645 cell_1rw
* cell instance $27805 r0 *1 121.965,125.58
X$27805 412 607 413 644 645 cell_1rw
* cell instance $27806 m0 *1 121.965,128.31
X$27806 412 609 413 644 645 cell_1rw
* cell instance $27807 m0 *1 121.965,131.04
X$27807 412 610 413 644 645 cell_1rw
* cell instance $27808 r0 *1 121.965,128.31
X$27808 412 608 413 644 645 cell_1rw
* cell instance $27809 r0 *1 121.965,131.04
X$27809 412 611 413 644 645 cell_1rw
* cell instance $27810 m0 *1 121.965,133.77
X$27810 412 612 413 644 645 cell_1rw
* cell instance $27811 r0 *1 121.965,133.77
X$27811 412 613 413 644 645 cell_1rw
* cell instance $27812 m0 *1 121.965,136.5
X$27812 412 615 413 644 645 cell_1rw
* cell instance $27813 r0 *1 121.965,136.5
X$27813 412 614 413 644 645 cell_1rw
* cell instance $27814 m0 *1 121.965,139.23
X$27814 412 617 413 644 645 cell_1rw
* cell instance $27815 r0 *1 121.965,139.23
X$27815 412 616 413 644 645 cell_1rw
* cell instance $27816 m0 *1 121.965,141.96
X$27816 412 618 413 644 645 cell_1rw
* cell instance $27817 r0 *1 121.965,141.96
X$27817 412 619 413 644 645 cell_1rw
* cell instance $27818 m0 *1 121.965,144.69
X$27818 412 620 413 644 645 cell_1rw
* cell instance $27819 r0 *1 121.965,144.69
X$27819 412 621 413 644 645 cell_1rw
* cell instance $27820 m0 *1 121.965,147.42
X$27820 412 622 413 644 645 cell_1rw
* cell instance $27821 r0 *1 121.965,147.42
X$27821 412 623 413 644 645 cell_1rw
* cell instance $27822 m0 *1 121.965,150.15
X$27822 412 624 413 644 645 cell_1rw
* cell instance $27823 r0 *1 121.965,150.15
X$27823 412 625 413 644 645 cell_1rw
* cell instance $27824 m0 *1 121.965,152.88
X$27824 412 626 413 644 645 cell_1rw
* cell instance $27825 m0 *1 121.965,155.61
X$27825 412 628 413 644 645 cell_1rw
* cell instance $27826 r0 *1 121.965,152.88
X$27826 412 627 413 644 645 cell_1rw
* cell instance $27827 m0 *1 121.965,158.34
X$27827 412 630 413 644 645 cell_1rw
* cell instance $27828 r0 *1 121.965,155.61
X$27828 412 629 413 644 645 cell_1rw
* cell instance $27829 r0 *1 121.965,158.34
X$27829 412 631 413 644 645 cell_1rw
* cell instance $27830 m0 *1 121.965,161.07
X$27830 412 632 413 644 645 cell_1rw
* cell instance $27831 r0 *1 121.965,161.07
X$27831 412 633 413 644 645 cell_1rw
* cell instance $27832 m0 *1 121.965,163.8
X$27832 412 634 413 644 645 cell_1rw
* cell instance $27833 m0 *1 121.965,166.53
X$27833 412 637 413 644 645 cell_1rw
* cell instance $27834 r0 *1 121.965,163.8
X$27834 412 635 413 644 645 cell_1rw
* cell instance $27835 r0 *1 121.965,166.53
X$27835 412 636 413 644 645 cell_1rw
* cell instance $27836 m0 *1 121.965,169.26
X$27836 412 639 413 644 645 cell_1rw
* cell instance $27837 r0 *1 121.965,169.26
X$27837 412 638 413 644 645 cell_1rw
* cell instance $27838 m0 *1 121.965,171.99
X$27838 412 640 413 644 645 cell_1rw
* cell instance $27839 r0 *1 121.965,171.99
X$27839 412 641 413 644 645 cell_1rw
* cell instance $27840 m0 *1 121.965,174.72
X$27840 412 642 413 644 645 cell_1rw
* cell instance $27841 r0 *1 121.965,174.72
X$27841 412 643 413 644 645 cell_1rw
* cell instance $27842 m0 *1 122.67,90.09
X$27842 414 581 415 644 645 cell_1rw
* cell instance $27843 r0 *1 122.67,90.09
X$27843 414 580 415 644 645 cell_1rw
* cell instance $27844 m0 *1 122.67,92.82
X$27844 414 583 415 644 645 cell_1rw
* cell instance $27845 r0 *1 122.67,92.82
X$27845 414 582 415 644 645 cell_1rw
* cell instance $27846 m0 *1 122.67,95.55
X$27846 414 584 415 644 645 cell_1rw
* cell instance $27847 r0 *1 122.67,95.55
X$27847 414 585 415 644 645 cell_1rw
* cell instance $27848 m0 *1 122.67,98.28
X$27848 414 586 415 644 645 cell_1rw
* cell instance $27849 r0 *1 122.67,98.28
X$27849 414 587 415 644 645 cell_1rw
* cell instance $27850 m0 *1 122.67,101.01
X$27850 414 588 415 644 645 cell_1rw
* cell instance $27851 r0 *1 122.67,101.01
X$27851 414 589 415 644 645 cell_1rw
* cell instance $27852 m0 *1 122.67,103.74
X$27852 414 590 415 644 645 cell_1rw
* cell instance $27853 r0 *1 122.67,103.74
X$27853 414 591 415 644 645 cell_1rw
* cell instance $27854 m0 *1 122.67,106.47
X$27854 414 593 415 644 645 cell_1rw
* cell instance $27855 r0 *1 122.67,106.47
X$27855 414 592 415 644 645 cell_1rw
* cell instance $27856 m0 *1 122.67,109.2
X$27856 414 594 415 644 645 cell_1rw
* cell instance $27857 r0 *1 122.67,109.2
X$27857 414 595 415 644 645 cell_1rw
* cell instance $27858 m0 *1 122.67,111.93
X$27858 414 597 415 644 645 cell_1rw
* cell instance $27859 r0 *1 122.67,111.93
X$27859 414 596 415 644 645 cell_1rw
* cell instance $27860 m0 *1 122.67,114.66
X$27860 414 598 415 644 645 cell_1rw
* cell instance $27861 r0 *1 122.67,114.66
X$27861 414 599 415 644 645 cell_1rw
* cell instance $27862 m0 *1 122.67,117.39
X$27862 414 600 415 644 645 cell_1rw
* cell instance $27863 m0 *1 122.67,120.12
X$27863 414 602 415 644 645 cell_1rw
* cell instance $27864 r0 *1 122.67,117.39
X$27864 414 601 415 644 645 cell_1rw
* cell instance $27865 r0 *1 122.67,120.12
X$27865 414 603 415 644 645 cell_1rw
* cell instance $27866 m0 *1 122.67,122.85
X$27866 414 604 415 644 645 cell_1rw
* cell instance $27867 r0 *1 122.67,122.85
X$27867 414 605 415 644 645 cell_1rw
* cell instance $27868 m0 *1 122.67,125.58
X$27868 414 606 415 644 645 cell_1rw
* cell instance $27869 r0 *1 122.67,125.58
X$27869 414 607 415 644 645 cell_1rw
* cell instance $27870 m0 *1 122.67,128.31
X$27870 414 609 415 644 645 cell_1rw
* cell instance $27871 r0 *1 122.67,128.31
X$27871 414 608 415 644 645 cell_1rw
* cell instance $27872 m0 *1 122.67,131.04
X$27872 414 610 415 644 645 cell_1rw
* cell instance $27873 r0 *1 122.67,131.04
X$27873 414 611 415 644 645 cell_1rw
* cell instance $27874 m0 *1 122.67,133.77
X$27874 414 612 415 644 645 cell_1rw
* cell instance $27875 m0 *1 122.67,136.5
X$27875 414 615 415 644 645 cell_1rw
* cell instance $27876 r0 *1 122.67,133.77
X$27876 414 613 415 644 645 cell_1rw
* cell instance $27877 r0 *1 122.67,136.5
X$27877 414 614 415 644 645 cell_1rw
* cell instance $27878 m0 *1 122.67,139.23
X$27878 414 617 415 644 645 cell_1rw
* cell instance $27879 r0 *1 122.67,139.23
X$27879 414 616 415 644 645 cell_1rw
* cell instance $27880 m0 *1 122.67,141.96
X$27880 414 618 415 644 645 cell_1rw
* cell instance $27881 r0 *1 122.67,141.96
X$27881 414 619 415 644 645 cell_1rw
* cell instance $27882 m0 *1 122.67,144.69
X$27882 414 620 415 644 645 cell_1rw
* cell instance $27883 r0 *1 122.67,144.69
X$27883 414 621 415 644 645 cell_1rw
* cell instance $27884 m0 *1 122.67,147.42
X$27884 414 622 415 644 645 cell_1rw
* cell instance $27885 r0 *1 122.67,147.42
X$27885 414 623 415 644 645 cell_1rw
* cell instance $27886 m0 *1 122.67,150.15
X$27886 414 624 415 644 645 cell_1rw
* cell instance $27887 r0 *1 122.67,150.15
X$27887 414 625 415 644 645 cell_1rw
* cell instance $27888 m0 *1 122.67,152.88
X$27888 414 626 415 644 645 cell_1rw
* cell instance $27889 m0 *1 122.67,155.61
X$27889 414 628 415 644 645 cell_1rw
* cell instance $27890 r0 *1 122.67,152.88
X$27890 414 627 415 644 645 cell_1rw
* cell instance $27891 r0 *1 122.67,155.61
X$27891 414 629 415 644 645 cell_1rw
* cell instance $27892 m0 *1 122.67,158.34
X$27892 414 630 415 644 645 cell_1rw
* cell instance $27893 r0 *1 122.67,158.34
X$27893 414 631 415 644 645 cell_1rw
* cell instance $27894 m0 *1 122.67,161.07
X$27894 414 632 415 644 645 cell_1rw
* cell instance $27895 r0 *1 122.67,161.07
X$27895 414 633 415 644 645 cell_1rw
* cell instance $27896 m0 *1 122.67,163.8
X$27896 414 634 415 644 645 cell_1rw
* cell instance $27897 m0 *1 122.67,166.53
X$27897 414 637 415 644 645 cell_1rw
* cell instance $27898 r0 *1 122.67,163.8
X$27898 414 635 415 644 645 cell_1rw
* cell instance $27899 r0 *1 122.67,166.53
X$27899 414 636 415 644 645 cell_1rw
* cell instance $27900 m0 *1 122.67,169.26
X$27900 414 639 415 644 645 cell_1rw
* cell instance $27901 r0 *1 122.67,169.26
X$27901 414 638 415 644 645 cell_1rw
* cell instance $27902 m0 *1 122.67,171.99
X$27902 414 640 415 644 645 cell_1rw
* cell instance $27903 m0 *1 122.67,174.72
X$27903 414 642 415 644 645 cell_1rw
* cell instance $27904 r0 *1 122.67,171.99
X$27904 414 641 415 644 645 cell_1rw
* cell instance $27905 r0 *1 122.67,174.72
X$27905 414 643 415 644 645 cell_1rw
* cell instance $27906 m0 *1 123.375,90.09
X$27906 416 581 417 644 645 cell_1rw
* cell instance $27907 r0 *1 123.375,90.09
X$27907 416 580 417 644 645 cell_1rw
* cell instance $27908 m0 *1 123.375,92.82
X$27908 416 583 417 644 645 cell_1rw
* cell instance $27909 r0 *1 123.375,92.82
X$27909 416 582 417 644 645 cell_1rw
* cell instance $27910 m0 *1 123.375,95.55
X$27910 416 584 417 644 645 cell_1rw
* cell instance $27911 r0 *1 123.375,95.55
X$27911 416 585 417 644 645 cell_1rw
* cell instance $27912 m0 *1 123.375,98.28
X$27912 416 586 417 644 645 cell_1rw
* cell instance $27913 r0 *1 123.375,98.28
X$27913 416 587 417 644 645 cell_1rw
* cell instance $27914 m0 *1 123.375,101.01
X$27914 416 588 417 644 645 cell_1rw
* cell instance $27915 r0 *1 123.375,101.01
X$27915 416 589 417 644 645 cell_1rw
* cell instance $27916 m0 *1 123.375,103.74
X$27916 416 590 417 644 645 cell_1rw
* cell instance $27917 r0 *1 123.375,103.74
X$27917 416 591 417 644 645 cell_1rw
* cell instance $27918 m0 *1 123.375,106.47
X$27918 416 593 417 644 645 cell_1rw
* cell instance $27919 r0 *1 123.375,106.47
X$27919 416 592 417 644 645 cell_1rw
* cell instance $27920 m0 *1 123.375,109.2
X$27920 416 594 417 644 645 cell_1rw
* cell instance $27921 r0 *1 123.375,109.2
X$27921 416 595 417 644 645 cell_1rw
* cell instance $27922 m0 *1 123.375,111.93
X$27922 416 597 417 644 645 cell_1rw
* cell instance $27923 r0 *1 123.375,111.93
X$27923 416 596 417 644 645 cell_1rw
* cell instance $27924 m0 *1 123.375,114.66
X$27924 416 598 417 644 645 cell_1rw
* cell instance $27925 r0 *1 123.375,114.66
X$27925 416 599 417 644 645 cell_1rw
* cell instance $27926 m0 *1 123.375,117.39
X$27926 416 600 417 644 645 cell_1rw
* cell instance $27927 r0 *1 123.375,117.39
X$27927 416 601 417 644 645 cell_1rw
* cell instance $27928 m0 *1 123.375,120.12
X$27928 416 602 417 644 645 cell_1rw
* cell instance $27929 m0 *1 123.375,122.85
X$27929 416 604 417 644 645 cell_1rw
* cell instance $27930 r0 *1 123.375,120.12
X$27930 416 603 417 644 645 cell_1rw
* cell instance $27931 r0 *1 123.375,122.85
X$27931 416 605 417 644 645 cell_1rw
* cell instance $27932 m0 *1 123.375,125.58
X$27932 416 606 417 644 645 cell_1rw
* cell instance $27933 r0 *1 123.375,125.58
X$27933 416 607 417 644 645 cell_1rw
* cell instance $27934 m0 *1 123.375,128.31
X$27934 416 609 417 644 645 cell_1rw
* cell instance $27935 r0 *1 123.375,128.31
X$27935 416 608 417 644 645 cell_1rw
* cell instance $27936 m0 *1 123.375,131.04
X$27936 416 610 417 644 645 cell_1rw
* cell instance $27937 r0 *1 123.375,131.04
X$27937 416 611 417 644 645 cell_1rw
* cell instance $27938 m0 *1 123.375,133.77
X$27938 416 612 417 644 645 cell_1rw
* cell instance $27939 r0 *1 123.375,133.77
X$27939 416 613 417 644 645 cell_1rw
* cell instance $27940 m0 *1 123.375,136.5
X$27940 416 615 417 644 645 cell_1rw
* cell instance $27941 r0 *1 123.375,136.5
X$27941 416 614 417 644 645 cell_1rw
* cell instance $27942 m0 *1 123.375,139.23
X$27942 416 617 417 644 645 cell_1rw
* cell instance $27943 r0 *1 123.375,139.23
X$27943 416 616 417 644 645 cell_1rw
* cell instance $27944 m0 *1 123.375,141.96
X$27944 416 618 417 644 645 cell_1rw
* cell instance $27945 r0 *1 123.375,141.96
X$27945 416 619 417 644 645 cell_1rw
* cell instance $27946 m0 *1 123.375,144.69
X$27946 416 620 417 644 645 cell_1rw
* cell instance $27947 m0 *1 123.375,147.42
X$27947 416 622 417 644 645 cell_1rw
* cell instance $27948 r0 *1 123.375,144.69
X$27948 416 621 417 644 645 cell_1rw
* cell instance $27949 r0 *1 123.375,147.42
X$27949 416 623 417 644 645 cell_1rw
* cell instance $27950 m0 *1 123.375,150.15
X$27950 416 624 417 644 645 cell_1rw
* cell instance $27951 r0 *1 123.375,150.15
X$27951 416 625 417 644 645 cell_1rw
* cell instance $27952 m0 *1 123.375,152.88
X$27952 416 626 417 644 645 cell_1rw
* cell instance $27953 r0 *1 123.375,152.88
X$27953 416 627 417 644 645 cell_1rw
* cell instance $27954 m0 *1 123.375,155.61
X$27954 416 628 417 644 645 cell_1rw
* cell instance $27955 r0 *1 123.375,155.61
X$27955 416 629 417 644 645 cell_1rw
* cell instance $27956 m0 *1 123.375,158.34
X$27956 416 630 417 644 645 cell_1rw
* cell instance $27957 r0 *1 123.375,158.34
X$27957 416 631 417 644 645 cell_1rw
* cell instance $27958 m0 *1 123.375,161.07
X$27958 416 632 417 644 645 cell_1rw
* cell instance $27959 r0 *1 123.375,161.07
X$27959 416 633 417 644 645 cell_1rw
* cell instance $27960 m0 *1 123.375,163.8
X$27960 416 634 417 644 645 cell_1rw
* cell instance $27961 m0 *1 123.375,166.53
X$27961 416 637 417 644 645 cell_1rw
* cell instance $27962 r0 *1 123.375,163.8
X$27962 416 635 417 644 645 cell_1rw
* cell instance $27963 m0 *1 123.375,169.26
X$27963 416 639 417 644 645 cell_1rw
* cell instance $27964 r0 *1 123.375,166.53
X$27964 416 636 417 644 645 cell_1rw
* cell instance $27965 r0 *1 123.375,169.26
X$27965 416 638 417 644 645 cell_1rw
* cell instance $27966 m0 *1 123.375,171.99
X$27966 416 640 417 644 645 cell_1rw
* cell instance $27967 r0 *1 123.375,171.99
X$27967 416 641 417 644 645 cell_1rw
* cell instance $27968 m0 *1 123.375,174.72
X$27968 416 642 417 644 645 cell_1rw
* cell instance $27969 r0 *1 123.375,174.72
X$27969 416 643 417 644 645 cell_1rw
* cell instance $27970 m0 *1 124.08,90.09
X$27970 418 581 419 644 645 cell_1rw
* cell instance $27971 m0 *1 124.08,92.82
X$27971 418 583 419 644 645 cell_1rw
* cell instance $27972 r0 *1 124.08,90.09
X$27972 418 580 419 644 645 cell_1rw
* cell instance $27973 r0 *1 124.08,92.82
X$27973 418 582 419 644 645 cell_1rw
* cell instance $27974 m0 *1 124.08,95.55
X$27974 418 584 419 644 645 cell_1rw
* cell instance $27975 r0 *1 124.08,95.55
X$27975 418 585 419 644 645 cell_1rw
* cell instance $27976 m0 *1 124.08,98.28
X$27976 418 586 419 644 645 cell_1rw
* cell instance $27977 r0 *1 124.08,98.28
X$27977 418 587 419 644 645 cell_1rw
* cell instance $27978 m0 *1 124.08,101.01
X$27978 418 588 419 644 645 cell_1rw
* cell instance $27979 r0 *1 124.08,101.01
X$27979 418 589 419 644 645 cell_1rw
* cell instance $27980 m0 *1 124.08,103.74
X$27980 418 590 419 644 645 cell_1rw
* cell instance $27981 r0 *1 124.08,103.74
X$27981 418 591 419 644 645 cell_1rw
* cell instance $27982 m0 *1 124.08,106.47
X$27982 418 593 419 644 645 cell_1rw
* cell instance $27983 m0 *1 124.08,109.2
X$27983 418 594 419 644 645 cell_1rw
* cell instance $27984 r0 *1 124.08,106.47
X$27984 418 592 419 644 645 cell_1rw
* cell instance $27985 r0 *1 124.08,109.2
X$27985 418 595 419 644 645 cell_1rw
* cell instance $27986 m0 *1 124.08,111.93
X$27986 418 597 419 644 645 cell_1rw
* cell instance $27987 r0 *1 124.08,111.93
X$27987 418 596 419 644 645 cell_1rw
* cell instance $27988 m0 *1 124.08,114.66
X$27988 418 598 419 644 645 cell_1rw
* cell instance $27989 r0 *1 124.08,114.66
X$27989 418 599 419 644 645 cell_1rw
* cell instance $27990 m0 *1 124.08,117.39
X$27990 418 600 419 644 645 cell_1rw
* cell instance $27991 r0 *1 124.08,117.39
X$27991 418 601 419 644 645 cell_1rw
* cell instance $27992 m0 *1 124.08,120.12
X$27992 418 602 419 644 645 cell_1rw
* cell instance $27993 r0 *1 124.08,120.12
X$27993 418 603 419 644 645 cell_1rw
* cell instance $27994 m0 *1 124.08,122.85
X$27994 418 604 419 644 645 cell_1rw
* cell instance $27995 r0 *1 124.08,122.85
X$27995 418 605 419 644 645 cell_1rw
* cell instance $27996 m0 *1 124.08,125.58
X$27996 418 606 419 644 645 cell_1rw
* cell instance $27997 r0 *1 124.08,125.58
X$27997 418 607 419 644 645 cell_1rw
* cell instance $27998 m0 *1 124.08,128.31
X$27998 418 609 419 644 645 cell_1rw
* cell instance $27999 m0 *1 124.08,131.04
X$27999 418 610 419 644 645 cell_1rw
* cell instance $28000 r0 *1 124.08,128.31
X$28000 418 608 419 644 645 cell_1rw
* cell instance $28001 r0 *1 124.08,131.04
X$28001 418 611 419 644 645 cell_1rw
* cell instance $28002 m0 *1 124.08,133.77
X$28002 418 612 419 644 645 cell_1rw
* cell instance $28003 r0 *1 124.08,133.77
X$28003 418 613 419 644 645 cell_1rw
* cell instance $28004 m0 *1 124.08,136.5
X$28004 418 615 419 644 645 cell_1rw
* cell instance $28005 r0 *1 124.08,136.5
X$28005 418 614 419 644 645 cell_1rw
* cell instance $28006 m0 *1 124.08,139.23
X$28006 418 617 419 644 645 cell_1rw
* cell instance $28007 m0 *1 124.08,141.96
X$28007 418 618 419 644 645 cell_1rw
* cell instance $28008 r0 *1 124.08,139.23
X$28008 418 616 419 644 645 cell_1rw
* cell instance $28009 r0 *1 124.08,141.96
X$28009 418 619 419 644 645 cell_1rw
* cell instance $28010 m0 *1 124.08,144.69
X$28010 418 620 419 644 645 cell_1rw
* cell instance $28011 r0 *1 124.08,144.69
X$28011 418 621 419 644 645 cell_1rw
* cell instance $28012 m0 *1 124.08,147.42
X$28012 418 622 419 644 645 cell_1rw
* cell instance $28013 r0 *1 124.08,147.42
X$28013 418 623 419 644 645 cell_1rw
* cell instance $28014 m0 *1 124.08,150.15
X$28014 418 624 419 644 645 cell_1rw
* cell instance $28015 r0 *1 124.08,150.15
X$28015 418 625 419 644 645 cell_1rw
* cell instance $28016 m0 *1 124.08,152.88
X$28016 418 626 419 644 645 cell_1rw
* cell instance $28017 r0 *1 124.08,152.88
X$28017 418 627 419 644 645 cell_1rw
* cell instance $28018 m0 *1 124.08,155.61
X$28018 418 628 419 644 645 cell_1rw
* cell instance $28019 r0 *1 124.08,155.61
X$28019 418 629 419 644 645 cell_1rw
* cell instance $28020 m0 *1 124.08,158.34
X$28020 418 630 419 644 645 cell_1rw
* cell instance $28021 r0 *1 124.08,158.34
X$28021 418 631 419 644 645 cell_1rw
* cell instance $28022 m0 *1 124.08,161.07
X$28022 418 632 419 644 645 cell_1rw
* cell instance $28023 r0 *1 124.08,161.07
X$28023 418 633 419 644 645 cell_1rw
* cell instance $28024 m0 *1 124.08,163.8
X$28024 418 634 419 644 645 cell_1rw
* cell instance $28025 m0 *1 124.08,166.53
X$28025 418 637 419 644 645 cell_1rw
* cell instance $28026 r0 *1 124.08,163.8
X$28026 418 635 419 644 645 cell_1rw
* cell instance $28027 r0 *1 124.08,166.53
X$28027 418 636 419 644 645 cell_1rw
* cell instance $28028 m0 *1 124.08,169.26
X$28028 418 639 419 644 645 cell_1rw
* cell instance $28029 r0 *1 124.08,169.26
X$28029 418 638 419 644 645 cell_1rw
* cell instance $28030 m0 *1 124.08,171.99
X$28030 418 640 419 644 645 cell_1rw
* cell instance $28031 m0 *1 124.08,174.72
X$28031 418 642 419 644 645 cell_1rw
* cell instance $28032 r0 *1 124.08,171.99
X$28032 418 641 419 644 645 cell_1rw
* cell instance $28033 r0 *1 124.08,174.72
X$28033 418 643 419 644 645 cell_1rw
* cell instance $28034 m0 *1 124.785,90.09
X$28034 420 581 421 644 645 cell_1rw
* cell instance $28035 r0 *1 124.785,90.09
X$28035 420 580 421 644 645 cell_1rw
* cell instance $28036 m0 *1 124.785,92.82
X$28036 420 583 421 644 645 cell_1rw
* cell instance $28037 r0 *1 124.785,92.82
X$28037 420 582 421 644 645 cell_1rw
* cell instance $28038 m0 *1 124.785,95.55
X$28038 420 584 421 644 645 cell_1rw
* cell instance $28039 r0 *1 124.785,95.55
X$28039 420 585 421 644 645 cell_1rw
* cell instance $28040 m0 *1 124.785,98.28
X$28040 420 586 421 644 645 cell_1rw
* cell instance $28041 m0 *1 124.785,101.01
X$28041 420 588 421 644 645 cell_1rw
* cell instance $28042 r0 *1 124.785,98.28
X$28042 420 587 421 644 645 cell_1rw
* cell instance $28043 r0 *1 124.785,101.01
X$28043 420 589 421 644 645 cell_1rw
* cell instance $28044 m0 *1 124.785,103.74
X$28044 420 590 421 644 645 cell_1rw
* cell instance $28045 r0 *1 124.785,103.74
X$28045 420 591 421 644 645 cell_1rw
* cell instance $28046 m0 *1 124.785,106.47
X$28046 420 593 421 644 645 cell_1rw
* cell instance $28047 r0 *1 124.785,106.47
X$28047 420 592 421 644 645 cell_1rw
* cell instance $28048 m0 *1 124.785,109.2
X$28048 420 594 421 644 645 cell_1rw
* cell instance $28049 r0 *1 124.785,109.2
X$28049 420 595 421 644 645 cell_1rw
* cell instance $28050 m0 *1 124.785,111.93
X$28050 420 597 421 644 645 cell_1rw
* cell instance $28051 r0 *1 124.785,111.93
X$28051 420 596 421 644 645 cell_1rw
* cell instance $28052 m0 *1 124.785,114.66
X$28052 420 598 421 644 645 cell_1rw
* cell instance $28053 r0 *1 124.785,114.66
X$28053 420 599 421 644 645 cell_1rw
* cell instance $28054 m0 *1 124.785,117.39
X$28054 420 600 421 644 645 cell_1rw
* cell instance $28055 r0 *1 124.785,117.39
X$28055 420 601 421 644 645 cell_1rw
* cell instance $28056 m0 *1 124.785,120.12
X$28056 420 602 421 644 645 cell_1rw
* cell instance $28057 r0 *1 124.785,120.12
X$28057 420 603 421 644 645 cell_1rw
* cell instance $28058 m0 *1 124.785,122.85
X$28058 420 604 421 644 645 cell_1rw
* cell instance $28059 m0 *1 124.785,125.58
X$28059 420 606 421 644 645 cell_1rw
* cell instance $28060 r0 *1 124.785,122.85
X$28060 420 605 421 644 645 cell_1rw
* cell instance $28061 m0 *1 124.785,128.31
X$28061 420 609 421 644 645 cell_1rw
* cell instance $28062 r0 *1 124.785,125.58
X$28062 420 607 421 644 645 cell_1rw
* cell instance $28063 r0 *1 124.785,128.31
X$28063 420 608 421 644 645 cell_1rw
* cell instance $28064 m0 *1 124.785,131.04
X$28064 420 610 421 644 645 cell_1rw
* cell instance $28065 r0 *1 124.785,131.04
X$28065 420 611 421 644 645 cell_1rw
* cell instance $28066 m0 *1 124.785,133.77
X$28066 420 612 421 644 645 cell_1rw
* cell instance $28067 m0 *1 124.785,136.5
X$28067 420 615 421 644 645 cell_1rw
* cell instance $28068 r0 *1 124.785,133.77
X$28068 420 613 421 644 645 cell_1rw
* cell instance $28069 m0 *1 124.785,139.23
X$28069 420 617 421 644 645 cell_1rw
* cell instance $28070 r0 *1 124.785,136.5
X$28070 420 614 421 644 645 cell_1rw
* cell instance $28071 r0 *1 124.785,139.23
X$28071 420 616 421 644 645 cell_1rw
* cell instance $28072 m0 *1 124.785,141.96
X$28072 420 618 421 644 645 cell_1rw
* cell instance $28073 r0 *1 124.785,141.96
X$28073 420 619 421 644 645 cell_1rw
* cell instance $28074 m0 *1 124.785,144.69
X$28074 420 620 421 644 645 cell_1rw
* cell instance $28075 r0 *1 124.785,144.69
X$28075 420 621 421 644 645 cell_1rw
* cell instance $28076 m0 *1 124.785,147.42
X$28076 420 622 421 644 645 cell_1rw
* cell instance $28077 r0 *1 124.785,147.42
X$28077 420 623 421 644 645 cell_1rw
* cell instance $28078 m0 *1 124.785,150.15
X$28078 420 624 421 644 645 cell_1rw
* cell instance $28079 r0 *1 124.785,150.15
X$28079 420 625 421 644 645 cell_1rw
* cell instance $28080 m0 *1 124.785,152.88
X$28080 420 626 421 644 645 cell_1rw
* cell instance $28081 r0 *1 124.785,152.88
X$28081 420 627 421 644 645 cell_1rw
* cell instance $28082 m0 *1 124.785,155.61
X$28082 420 628 421 644 645 cell_1rw
* cell instance $28083 r0 *1 124.785,155.61
X$28083 420 629 421 644 645 cell_1rw
* cell instance $28084 m0 *1 124.785,158.34
X$28084 420 630 421 644 645 cell_1rw
* cell instance $28085 r0 *1 124.785,158.34
X$28085 420 631 421 644 645 cell_1rw
* cell instance $28086 m0 *1 124.785,161.07
X$28086 420 632 421 644 645 cell_1rw
* cell instance $28087 r0 *1 124.785,161.07
X$28087 420 633 421 644 645 cell_1rw
* cell instance $28088 m0 *1 124.785,163.8
X$28088 420 634 421 644 645 cell_1rw
* cell instance $28089 m0 *1 124.785,166.53
X$28089 420 637 421 644 645 cell_1rw
* cell instance $28090 r0 *1 124.785,163.8
X$28090 420 635 421 644 645 cell_1rw
* cell instance $28091 r0 *1 124.785,166.53
X$28091 420 636 421 644 645 cell_1rw
* cell instance $28092 m0 *1 124.785,169.26
X$28092 420 639 421 644 645 cell_1rw
* cell instance $28093 r0 *1 124.785,169.26
X$28093 420 638 421 644 645 cell_1rw
* cell instance $28094 m0 *1 124.785,171.99
X$28094 420 640 421 644 645 cell_1rw
* cell instance $28095 r0 *1 124.785,171.99
X$28095 420 641 421 644 645 cell_1rw
* cell instance $28096 m0 *1 124.785,174.72
X$28096 420 642 421 644 645 cell_1rw
* cell instance $28097 r0 *1 124.785,174.72
X$28097 420 643 421 644 645 cell_1rw
* cell instance $28098 m0 *1 125.49,90.09
X$28098 422 581 423 644 645 cell_1rw
* cell instance $28099 m0 *1 125.49,92.82
X$28099 422 583 423 644 645 cell_1rw
* cell instance $28100 r0 *1 125.49,90.09
X$28100 422 580 423 644 645 cell_1rw
* cell instance $28101 r0 *1 125.49,92.82
X$28101 422 582 423 644 645 cell_1rw
* cell instance $28102 m0 *1 125.49,95.55
X$28102 422 584 423 644 645 cell_1rw
* cell instance $28103 r0 *1 125.49,95.55
X$28103 422 585 423 644 645 cell_1rw
* cell instance $28104 m0 *1 125.49,98.28
X$28104 422 586 423 644 645 cell_1rw
* cell instance $28105 r0 *1 125.49,98.28
X$28105 422 587 423 644 645 cell_1rw
* cell instance $28106 m0 *1 125.49,101.01
X$28106 422 588 423 644 645 cell_1rw
* cell instance $28107 r0 *1 125.49,101.01
X$28107 422 589 423 644 645 cell_1rw
* cell instance $28108 m0 *1 125.49,103.74
X$28108 422 590 423 644 645 cell_1rw
* cell instance $28109 r0 *1 125.49,103.74
X$28109 422 591 423 644 645 cell_1rw
* cell instance $28110 m0 *1 125.49,106.47
X$28110 422 593 423 644 645 cell_1rw
* cell instance $28111 r0 *1 125.49,106.47
X$28111 422 592 423 644 645 cell_1rw
* cell instance $28112 m0 *1 125.49,109.2
X$28112 422 594 423 644 645 cell_1rw
* cell instance $28113 r0 *1 125.49,109.2
X$28113 422 595 423 644 645 cell_1rw
* cell instance $28114 m0 *1 125.49,111.93
X$28114 422 597 423 644 645 cell_1rw
* cell instance $28115 m0 *1 125.49,114.66
X$28115 422 598 423 644 645 cell_1rw
* cell instance $28116 r0 *1 125.49,111.93
X$28116 422 596 423 644 645 cell_1rw
* cell instance $28117 r0 *1 125.49,114.66
X$28117 422 599 423 644 645 cell_1rw
* cell instance $28118 m0 *1 125.49,117.39
X$28118 422 600 423 644 645 cell_1rw
* cell instance $28119 r0 *1 125.49,117.39
X$28119 422 601 423 644 645 cell_1rw
* cell instance $28120 m0 *1 125.49,120.12
X$28120 422 602 423 644 645 cell_1rw
* cell instance $28121 r0 *1 125.49,120.12
X$28121 422 603 423 644 645 cell_1rw
* cell instance $28122 m0 *1 125.49,122.85
X$28122 422 604 423 644 645 cell_1rw
* cell instance $28123 r0 *1 125.49,122.85
X$28123 422 605 423 644 645 cell_1rw
* cell instance $28124 m0 *1 125.49,125.58
X$28124 422 606 423 644 645 cell_1rw
* cell instance $28125 r0 *1 125.49,125.58
X$28125 422 607 423 644 645 cell_1rw
* cell instance $28126 m0 *1 125.49,128.31
X$28126 422 609 423 644 645 cell_1rw
* cell instance $28127 r0 *1 125.49,128.31
X$28127 422 608 423 644 645 cell_1rw
* cell instance $28128 m0 *1 125.49,131.04
X$28128 422 610 423 644 645 cell_1rw
* cell instance $28129 r0 *1 125.49,131.04
X$28129 422 611 423 644 645 cell_1rw
* cell instance $28130 m0 *1 125.49,133.77
X$28130 422 612 423 644 645 cell_1rw
* cell instance $28131 r0 *1 125.49,133.77
X$28131 422 613 423 644 645 cell_1rw
* cell instance $28132 m0 *1 125.49,136.5
X$28132 422 615 423 644 645 cell_1rw
* cell instance $28133 m0 *1 125.49,139.23
X$28133 422 617 423 644 645 cell_1rw
* cell instance $28134 r0 *1 125.49,136.5
X$28134 422 614 423 644 645 cell_1rw
* cell instance $28135 r0 *1 125.49,139.23
X$28135 422 616 423 644 645 cell_1rw
* cell instance $28136 m0 *1 125.49,141.96
X$28136 422 618 423 644 645 cell_1rw
* cell instance $28137 r0 *1 125.49,141.96
X$28137 422 619 423 644 645 cell_1rw
* cell instance $28138 m0 *1 125.49,144.69
X$28138 422 620 423 644 645 cell_1rw
* cell instance $28139 r0 *1 125.49,144.69
X$28139 422 621 423 644 645 cell_1rw
* cell instance $28140 m0 *1 125.49,147.42
X$28140 422 622 423 644 645 cell_1rw
* cell instance $28141 r0 *1 125.49,147.42
X$28141 422 623 423 644 645 cell_1rw
* cell instance $28142 m0 *1 125.49,150.15
X$28142 422 624 423 644 645 cell_1rw
* cell instance $28143 r0 *1 125.49,150.15
X$28143 422 625 423 644 645 cell_1rw
* cell instance $28144 m0 *1 125.49,152.88
X$28144 422 626 423 644 645 cell_1rw
* cell instance $28145 m0 *1 125.49,155.61
X$28145 422 628 423 644 645 cell_1rw
* cell instance $28146 r0 *1 125.49,152.88
X$28146 422 627 423 644 645 cell_1rw
* cell instance $28147 r0 *1 125.49,155.61
X$28147 422 629 423 644 645 cell_1rw
* cell instance $28148 m0 *1 125.49,158.34
X$28148 422 630 423 644 645 cell_1rw
* cell instance $28149 m0 *1 125.49,161.07
X$28149 422 632 423 644 645 cell_1rw
* cell instance $28150 r0 *1 125.49,158.34
X$28150 422 631 423 644 645 cell_1rw
* cell instance $28151 r0 *1 125.49,161.07
X$28151 422 633 423 644 645 cell_1rw
* cell instance $28152 m0 *1 125.49,163.8
X$28152 422 634 423 644 645 cell_1rw
* cell instance $28153 r0 *1 125.49,163.8
X$28153 422 635 423 644 645 cell_1rw
* cell instance $28154 m0 *1 125.49,166.53
X$28154 422 637 423 644 645 cell_1rw
* cell instance $28155 m0 *1 125.49,169.26
X$28155 422 639 423 644 645 cell_1rw
* cell instance $28156 r0 *1 125.49,166.53
X$28156 422 636 423 644 645 cell_1rw
* cell instance $28157 r0 *1 125.49,169.26
X$28157 422 638 423 644 645 cell_1rw
* cell instance $28158 m0 *1 125.49,171.99
X$28158 422 640 423 644 645 cell_1rw
* cell instance $28159 r0 *1 125.49,171.99
X$28159 422 641 423 644 645 cell_1rw
* cell instance $28160 m0 *1 125.49,174.72
X$28160 422 642 423 644 645 cell_1rw
* cell instance $28161 r0 *1 125.49,174.72
X$28161 422 643 423 644 645 cell_1rw
* cell instance $28162 m0 *1 126.195,90.09
X$28162 424 581 425 644 645 cell_1rw
* cell instance $28163 r0 *1 126.195,90.09
X$28163 424 580 425 644 645 cell_1rw
* cell instance $28164 m0 *1 126.195,92.82
X$28164 424 583 425 644 645 cell_1rw
* cell instance $28165 r0 *1 126.195,92.82
X$28165 424 582 425 644 645 cell_1rw
* cell instance $28166 m0 *1 126.195,95.55
X$28166 424 584 425 644 645 cell_1rw
* cell instance $28167 m0 *1 126.195,98.28
X$28167 424 586 425 644 645 cell_1rw
* cell instance $28168 r0 *1 126.195,95.55
X$28168 424 585 425 644 645 cell_1rw
* cell instance $28169 r0 *1 126.195,98.28
X$28169 424 587 425 644 645 cell_1rw
* cell instance $28170 m0 *1 126.195,101.01
X$28170 424 588 425 644 645 cell_1rw
* cell instance $28171 m0 *1 126.195,103.74
X$28171 424 590 425 644 645 cell_1rw
* cell instance $28172 r0 *1 126.195,101.01
X$28172 424 589 425 644 645 cell_1rw
* cell instance $28173 r0 *1 126.195,103.74
X$28173 424 591 425 644 645 cell_1rw
* cell instance $28174 m0 *1 126.195,106.47
X$28174 424 593 425 644 645 cell_1rw
* cell instance $28175 r0 *1 126.195,106.47
X$28175 424 592 425 644 645 cell_1rw
* cell instance $28176 m0 *1 126.195,109.2
X$28176 424 594 425 644 645 cell_1rw
* cell instance $28177 r0 *1 126.195,109.2
X$28177 424 595 425 644 645 cell_1rw
* cell instance $28178 m0 *1 126.195,111.93
X$28178 424 597 425 644 645 cell_1rw
* cell instance $28179 r0 *1 126.195,111.93
X$28179 424 596 425 644 645 cell_1rw
* cell instance $28180 m0 *1 126.195,114.66
X$28180 424 598 425 644 645 cell_1rw
* cell instance $28181 r0 *1 126.195,114.66
X$28181 424 599 425 644 645 cell_1rw
* cell instance $28182 m0 *1 126.195,117.39
X$28182 424 600 425 644 645 cell_1rw
* cell instance $28183 r0 *1 126.195,117.39
X$28183 424 601 425 644 645 cell_1rw
* cell instance $28184 m0 *1 126.195,120.12
X$28184 424 602 425 644 645 cell_1rw
* cell instance $28185 r0 *1 126.195,120.12
X$28185 424 603 425 644 645 cell_1rw
* cell instance $28186 m0 *1 126.195,122.85
X$28186 424 604 425 644 645 cell_1rw
* cell instance $28187 r0 *1 126.195,122.85
X$28187 424 605 425 644 645 cell_1rw
* cell instance $28188 m0 *1 126.195,125.58
X$28188 424 606 425 644 645 cell_1rw
* cell instance $28189 r0 *1 126.195,125.58
X$28189 424 607 425 644 645 cell_1rw
* cell instance $28190 m0 *1 126.195,128.31
X$28190 424 609 425 644 645 cell_1rw
* cell instance $28191 r0 *1 126.195,128.31
X$28191 424 608 425 644 645 cell_1rw
* cell instance $28192 m0 *1 126.195,131.04
X$28192 424 610 425 644 645 cell_1rw
* cell instance $28193 m0 *1 126.195,133.77
X$28193 424 612 425 644 645 cell_1rw
* cell instance $28194 r0 *1 126.195,131.04
X$28194 424 611 425 644 645 cell_1rw
* cell instance $28195 r0 *1 126.195,133.77
X$28195 424 613 425 644 645 cell_1rw
* cell instance $28196 m0 *1 126.195,136.5
X$28196 424 615 425 644 645 cell_1rw
* cell instance $28197 r0 *1 126.195,136.5
X$28197 424 614 425 644 645 cell_1rw
* cell instance $28198 m0 *1 126.195,139.23
X$28198 424 617 425 644 645 cell_1rw
* cell instance $28199 r0 *1 126.195,139.23
X$28199 424 616 425 644 645 cell_1rw
* cell instance $28200 m0 *1 126.195,141.96
X$28200 424 618 425 644 645 cell_1rw
* cell instance $28201 r0 *1 126.195,141.96
X$28201 424 619 425 644 645 cell_1rw
* cell instance $28202 m0 *1 126.195,144.69
X$28202 424 620 425 644 645 cell_1rw
* cell instance $28203 r0 *1 126.195,144.69
X$28203 424 621 425 644 645 cell_1rw
* cell instance $28204 m0 *1 126.195,147.42
X$28204 424 622 425 644 645 cell_1rw
* cell instance $28205 r0 *1 126.195,147.42
X$28205 424 623 425 644 645 cell_1rw
* cell instance $28206 m0 *1 126.195,150.15
X$28206 424 624 425 644 645 cell_1rw
* cell instance $28207 m0 *1 126.195,152.88
X$28207 424 626 425 644 645 cell_1rw
* cell instance $28208 r0 *1 126.195,150.15
X$28208 424 625 425 644 645 cell_1rw
* cell instance $28209 r0 *1 126.195,152.88
X$28209 424 627 425 644 645 cell_1rw
* cell instance $28210 m0 *1 126.195,155.61
X$28210 424 628 425 644 645 cell_1rw
* cell instance $28211 r0 *1 126.195,155.61
X$28211 424 629 425 644 645 cell_1rw
* cell instance $28212 m0 *1 126.195,158.34
X$28212 424 630 425 644 645 cell_1rw
* cell instance $28213 m0 *1 126.195,161.07
X$28213 424 632 425 644 645 cell_1rw
* cell instance $28214 r0 *1 126.195,158.34
X$28214 424 631 425 644 645 cell_1rw
* cell instance $28215 r0 *1 126.195,161.07
X$28215 424 633 425 644 645 cell_1rw
* cell instance $28216 m0 *1 126.195,163.8
X$28216 424 634 425 644 645 cell_1rw
* cell instance $28217 m0 *1 126.195,166.53
X$28217 424 637 425 644 645 cell_1rw
* cell instance $28218 r0 *1 126.195,163.8
X$28218 424 635 425 644 645 cell_1rw
* cell instance $28219 r0 *1 126.195,166.53
X$28219 424 636 425 644 645 cell_1rw
* cell instance $28220 m0 *1 126.195,169.26
X$28220 424 639 425 644 645 cell_1rw
* cell instance $28221 r0 *1 126.195,169.26
X$28221 424 638 425 644 645 cell_1rw
* cell instance $28222 m0 *1 126.195,171.99
X$28222 424 640 425 644 645 cell_1rw
* cell instance $28223 m0 *1 126.195,174.72
X$28223 424 642 425 644 645 cell_1rw
* cell instance $28224 r0 *1 126.195,171.99
X$28224 424 641 425 644 645 cell_1rw
* cell instance $28225 r0 *1 126.195,174.72
X$28225 424 643 425 644 645 cell_1rw
* cell instance $28226 m0 *1 126.9,90.09
X$28226 426 581 427 644 645 cell_1rw
* cell instance $28227 r0 *1 126.9,90.09
X$28227 426 580 427 644 645 cell_1rw
* cell instance $28228 m0 *1 126.9,92.82
X$28228 426 583 427 644 645 cell_1rw
* cell instance $28229 r0 *1 126.9,92.82
X$28229 426 582 427 644 645 cell_1rw
* cell instance $28230 m0 *1 126.9,95.55
X$28230 426 584 427 644 645 cell_1rw
* cell instance $28231 r0 *1 126.9,95.55
X$28231 426 585 427 644 645 cell_1rw
* cell instance $28232 m0 *1 126.9,98.28
X$28232 426 586 427 644 645 cell_1rw
* cell instance $28233 r0 *1 126.9,98.28
X$28233 426 587 427 644 645 cell_1rw
* cell instance $28234 m0 *1 126.9,101.01
X$28234 426 588 427 644 645 cell_1rw
* cell instance $28235 r0 *1 126.9,101.01
X$28235 426 589 427 644 645 cell_1rw
* cell instance $28236 m0 *1 126.9,103.74
X$28236 426 590 427 644 645 cell_1rw
* cell instance $28237 r0 *1 126.9,103.74
X$28237 426 591 427 644 645 cell_1rw
* cell instance $28238 m0 *1 126.9,106.47
X$28238 426 593 427 644 645 cell_1rw
* cell instance $28239 r0 *1 126.9,106.47
X$28239 426 592 427 644 645 cell_1rw
* cell instance $28240 m0 *1 126.9,109.2
X$28240 426 594 427 644 645 cell_1rw
* cell instance $28241 m0 *1 126.9,111.93
X$28241 426 597 427 644 645 cell_1rw
* cell instance $28242 r0 *1 126.9,109.2
X$28242 426 595 427 644 645 cell_1rw
* cell instance $28243 r0 *1 126.9,111.93
X$28243 426 596 427 644 645 cell_1rw
* cell instance $28244 m0 *1 126.9,114.66
X$28244 426 598 427 644 645 cell_1rw
* cell instance $28245 r0 *1 126.9,114.66
X$28245 426 599 427 644 645 cell_1rw
* cell instance $28246 m0 *1 126.9,117.39
X$28246 426 600 427 644 645 cell_1rw
* cell instance $28247 r0 *1 126.9,117.39
X$28247 426 601 427 644 645 cell_1rw
* cell instance $28248 m0 *1 126.9,120.12
X$28248 426 602 427 644 645 cell_1rw
* cell instance $28249 r0 *1 126.9,120.12
X$28249 426 603 427 644 645 cell_1rw
* cell instance $28250 m0 *1 126.9,122.85
X$28250 426 604 427 644 645 cell_1rw
* cell instance $28251 r0 *1 126.9,122.85
X$28251 426 605 427 644 645 cell_1rw
* cell instance $28252 m0 *1 126.9,125.58
X$28252 426 606 427 644 645 cell_1rw
* cell instance $28253 r0 *1 126.9,125.58
X$28253 426 607 427 644 645 cell_1rw
* cell instance $28254 m0 *1 126.9,128.31
X$28254 426 609 427 644 645 cell_1rw
* cell instance $28255 r0 *1 126.9,128.31
X$28255 426 608 427 644 645 cell_1rw
* cell instance $28256 m0 *1 126.9,131.04
X$28256 426 610 427 644 645 cell_1rw
* cell instance $28257 r0 *1 126.9,131.04
X$28257 426 611 427 644 645 cell_1rw
* cell instance $28258 m0 *1 126.9,133.77
X$28258 426 612 427 644 645 cell_1rw
* cell instance $28259 r0 *1 126.9,133.77
X$28259 426 613 427 644 645 cell_1rw
* cell instance $28260 m0 *1 126.9,136.5
X$28260 426 615 427 644 645 cell_1rw
* cell instance $28261 r0 *1 126.9,136.5
X$28261 426 614 427 644 645 cell_1rw
* cell instance $28262 m0 *1 126.9,139.23
X$28262 426 617 427 644 645 cell_1rw
* cell instance $28263 r0 *1 126.9,139.23
X$28263 426 616 427 644 645 cell_1rw
* cell instance $28264 m0 *1 126.9,141.96
X$28264 426 618 427 644 645 cell_1rw
* cell instance $28265 r0 *1 126.9,141.96
X$28265 426 619 427 644 645 cell_1rw
* cell instance $28266 m0 *1 126.9,144.69
X$28266 426 620 427 644 645 cell_1rw
* cell instance $28267 r0 *1 126.9,144.69
X$28267 426 621 427 644 645 cell_1rw
* cell instance $28268 m0 *1 126.9,147.42
X$28268 426 622 427 644 645 cell_1rw
* cell instance $28269 r0 *1 126.9,147.42
X$28269 426 623 427 644 645 cell_1rw
* cell instance $28270 m0 *1 126.9,150.15
X$28270 426 624 427 644 645 cell_1rw
* cell instance $28271 m0 *1 126.9,152.88
X$28271 426 626 427 644 645 cell_1rw
* cell instance $28272 r0 *1 126.9,150.15
X$28272 426 625 427 644 645 cell_1rw
* cell instance $28273 r0 *1 126.9,152.88
X$28273 426 627 427 644 645 cell_1rw
* cell instance $28274 m0 *1 126.9,155.61
X$28274 426 628 427 644 645 cell_1rw
* cell instance $28275 r0 *1 126.9,155.61
X$28275 426 629 427 644 645 cell_1rw
* cell instance $28276 m0 *1 126.9,158.34
X$28276 426 630 427 644 645 cell_1rw
* cell instance $28277 r0 *1 126.9,158.34
X$28277 426 631 427 644 645 cell_1rw
* cell instance $28278 m0 *1 126.9,161.07
X$28278 426 632 427 644 645 cell_1rw
* cell instance $28279 r0 *1 126.9,161.07
X$28279 426 633 427 644 645 cell_1rw
* cell instance $28280 m0 *1 126.9,163.8
X$28280 426 634 427 644 645 cell_1rw
* cell instance $28281 r0 *1 126.9,163.8
X$28281 426 635 427 644 645 cell_1rw
* cell instance $28282 m0 *1 126.9,166.53
X$28282 426 637 427 644 645 cell_1rw
* cell instance $28283 r0 *1 126.9,166.53
X$28283 426 636 427 644 645 cell_1rw
* cell instance $28284 m0 *1 126.9,169.26
X$28284 426 639 427 644 645 cell_1rw
* cell instance $28285 m0 *1 126.9,171.99
X$28285 426 640 427 644 645 cell_1rw
* cell instance $28286 r0 *1 126.9,169.26
X$28286 426 638 427 644 645 cell_1rw
* cell instance $28287 r0 *1 126.9,171.99
X$28287 426 641 427 644 645 cell_1rw
* cell instance $28288 m0 *1 126.9,174.72
X$28288 426 642 427 644 645 cell_1rw
* cell instance $28289 r0 *1 126.9,174.72
X$28289 426 643 427 644 645 cell_1rw
* cell instance $28290 m0 *1 127.605,90.09
X$28290 428 581 429 644 645 cell_1rw
* cell instance $28291 r0 *1 127.605,90.09
X$28291 428 580 429 644 645 cell_1rw
* cell instance $28292 m0 *1 127.605,92.82
X$28292 428 583 429 644 645 cell_1rw
* cell instance $28293 r0 *1 127.605,92.82
X$28293 428 582 429 644 645 cell_1rw
* cell instance $28294 m0 *1 127.605,95.55
X$28294 428 584 429 644 645 cell_1rw
* cell instance $28295 r0 *1 127.605,95.55
X$28295 428 585 429 644 645 cell_1rw
* cell instance $28296 m0 *1 127.605,98.28
X$28296 428 586 429 644 645 cell_1rw
* cell instance $28297 m0 *1 127.605,101.01
X$28297 428 588 429 644 645 cell_1rw
* cell instance $28298 r0 *1 127.605,98.28
X$28298 428 587 429 644 645 cell_1rw
* cell instance $28299 r0 *1 127.605,101.01
X$28299 428 589 429 644 645 cell_1rw
* cell instance $28300 m0 *1 127.605,103.74
X$28300 428 590 429 644 645 cell_1rw
* cell instance $28301 r0 *1 127.605,103.74
X$28301 428 591 429 644 645 cell_1rw
* cell instance $28302 m0 *1 127.605,106.47
X$28302 428 593 429 644 645 cell_1rw
* cell instance $28303 m0 *1 127.605,109.2
X$28303 428 594 429 644 645 cell_1rw
* cell instance $28304 r0 *1 127.605,106.47
X$28304 428 592 429 644 645 cell_1rw
* cell instance $28305 r0 *1 127.605,109.2
X$28305 428 595 429 644 645 cell_1rw
* cell instance $28306 m0 *1 127.605,111.93
X$28306 428 597 429 644 645 cell_1rw
* cell instance $28307 r0 *1 127.605,111.93
X$28307 428 596 429 644 645 cell_1rw
* cell instance $28308 m0 *1 127.605,114.66
X$28308 428 598 429 644 645 cell_1rw
* cell instance $28309 m0 *1 127.605,117.39
X$28309 428 600 429 644 645 cell_1rw
* cell instance $28310 r0 *1 127.605,114.66
X$28310 428 599 429 644 645 cell_1rw
* cell instance $28311 m0 *1 127.605,120.12
X$28311 428 602 429 644 645 cell_1rw
* cell instance $28312 r0 *1 127.605,117.39
X$28312 428 601 429 644 645 cell_1rw
* cell instance $28313 r0 *1 127.605,120.12
X$28313 428 603 429 644 645 cell_1rw
* cell instance $28314 m0 *1 127.605,122.85
X$28314 428 604 429 644 645 cell_1rw
* cell instance $28315 m0 *1 127.605,125.58
X$28315 428 606 429 644 645 cell_1rw
* cell instance $28316 r0 *1 127.605,122.85
X$28316 428 605 429 644 645 cell_1rw
* cell instance $28317 m0 *1 127.605,128.31
X$28317 428 609 429 644 645 cell_1rw
* cell instance $28318 r0 *1 127.605,125.58
X$28318 428 607 429 644 645 cell_1rw
* cell instance $28319 r0 *1 127.605,128.31
X$28319 428 608 429 644 645 cell_1rw
* cell instance $28320 m0 *1 127.605,131.04
X$28320 428 610 429 644 645 cell_1rw
* cell instance $28321 m0 *1 127.605,133.77
X$28321 428 612 429 644 645 cell_1rw
* cell instance $28322 r0 *1 127.605,131.04
X$28322 428 611 429 644 645 cell_1rw
* cell instance $28323 r0 *1 127.605,133.77
X$28323 428 613 429 644 645 cell_1rw
* cell instance $28324 m0 *1 127.605,136.5
X$28324 428 615 429 644 645 cell_1rw
* cell instance $28325 r0 *1 127.605,136.5
X$28325 428 614 429 644 645 cell_1rw
* cell instance $28326 m0 *1 127.605,139.23
X$28326 428 617 429 644 645 cell_1rw
* cell instance $28327 r0 *1 127.605,139.23
X$28327 428 616 429 644 645 cell_1rw
* cell instance $28328 m0 *1 127.605,141.96
X$28328 428 618 429 644 645 cell_1rw
* cell instance $28329 r0 *1 127.605,141.96
X$28329 428 619 429 644 645 cell_1rw
* cell instance $28330 m0 *1 127.605,144.69
X$28330 428 620 429 644 645 cell_1rw
* cell instance $28331 r0 *1 127.605,144.69
X$28331 428 621 429 644 645 cell_1rw
* cell instance $28332 m0 *1 127.605,147.42
X$28332 428 622 429 644 645 cell_1rw
* cell instance $28333 r0 *1 127.605,147.42
X$28333 428 623 429 644 645 cell_1rw
* cell instance $28334 m0 *1 127.605,150.15
X$28334 428 624 429 644 645 cell_1rw
* cell instance $28335 r0 *1 127.605,150.15
X$28335 428 625 429 644 645 cell_1rw
* cell instance $28336 m0 *1 127.605,152.88
X$28336 428 626 429 644 645 cell_1rw
* cell instance $28337 r0 *1 127.605,152.88
X$28337 428 627 429 644 645 cell_1rw
* cell instance $28338 m0 *1 127.605,155.61
X$28338 428 628 429 644 645 cell_1rw
* cell instance $28339 r0 *1 127.605,155.61
X$28339 428 629 429 644 645 cell_1rw
* cell instance $28340 m0 *1 127.605,158.34
X$28340 428 630 429 644 645 cell_1rw
* cell instance $28341 r0 *1 127.605,158.34
X$28341 428 631 429 644 645 cell_1rw
* cell instance $28342 m0 *1 127.605,161.07
X$28342 428 632 429 644 645 cell_1rw
* cell instance $28343 r0 *1 127.605,161.07
X$28343 428 633 429 644 645 cell_1rw
* cell instance $28344 m0 *1 127.605,163.8
X$28344 428 634 429 644 645 cell_1rw
* cell instance $28345 r0 *1 127.605,163.8
X$28345 428 635 429 644 645 cell_1rw
* cell instance $28346 m0 *1 127.605,166.53
X$28346 428 637 429 644 645 cell_1rw
* cell instance $28347 r0 *1 127.605,166.53
X$28347 428 636 429 644 645 cell_1rw
* cell instance $28348 m0 *1 127.605,169.26
X$28348 428 639 429 644 645 cell_1rw
* cell instance $28349 r0 *1 127.605,169.26
X$28349 428 638 429 644 645 cell_1rw
* cell instance $28350 m0 *1 127.605,171.99
X$28350 428 640 429 644 645 cell_1rw
* cell instance $28351 r0 *1 127.605,171.99
X$28351 428 641 429 644 645 cell_1rw
* cell instance $28352 m0 *1 127.605,174.72
X$28352 428 642 429 644 645 cell_1rw
* cell instance $28353 r0 *1 127.605,174.72
X$28353 428 643 429 644 645 cell_1rw
* cell instance $28354 m0 *1 128.31,90.09
X$28354 430 581 431 644 645 cell_1rw
* cell instance $28355 m0 *1 128.31,92.82
X$28355 430 583 431 644 645 cell_1rw
* cell instance $28356 r0 *1 128.31,90.09
X$28356 430 580 431 644 645 cell_1rw
* cell instance $28357 r0 *1 128.31,92.82
X$28357 430 582 431 644 645 cell_1rw
* cell instance $28358 m0 *1 128.31,95.55
X$28358 430 584 431 644 645 cell_1rw
* cell instance $28359 r0 *1 128.31,95.55
X$28359 430 585 431 644 645 cell_1rw
* cell instance $28360 m0 *1 128.31,98.28
X$28360 430 586 431 644 645 cell_1rw
* cell instance $28361 r0 *1 128.31,98.28
X$28361 430 587 431 644 645 cell_1rw
* cell instance $28362 m0 *1 128.31,101.01
X$28362 430 588 431 644 645 cell_1rw
* cell instance $28363 r0 *1 128.31,101.01
X$28363 430 589 431 644 645 cell_1rw
* cell instance $28364 m0 *1 128.31,103.74
X$28364 430 590 431 644 645 cell_1rw
* cell instance $28365 r0 *1 128.31,103.74
X$28365 430 591 431 644 645 cell_1rw
* cell instance $28366 m0 *1 128.31,106.47
X$28366 430 593 431 644 645 cell_1rw
* cell instance $28367 r0 *1 128.31,106.47
X$28367 430 592 431 644 645 cell_1rw
* cell instance $28368 m0 *1 128.31,109.2
X$28368 430 594 431 644 645 cell_1rw
* cell instance $28369 r0 *1 128.31,109.2
X$28369 430 595 431 644 645 cell_1rw
* cell instance $28370 m0 *1 128.31,111.93
X$28370 430 597 431 644 645 cell_1rw
* cell instance $28371 r0 *1 128.31,111.93
X$28371 430 596 431 644 645 cell_1rw
* cell instance $28372 m0 *1 128.31,114.66
X$28372 430 598 431 644 645 cell_1rw
* cell instance $28373 m0 *1 128.31,117.39
X$28373 430 600 431 644 645 cell_1rw
* cell instance $28374 r0 *1 128.31,114.66
X$28374 430 599 431 644 645 cell_1rw
* cell instance $28375 r0 *1 128.31,117.39
X$28375 430 601 431 644 645 cell_1rw
* cell instance $28376 m0 *1 128.31,120.12
X$28376 430 602 431 644 645 cell_1rw
* cell instance $28377 r0 *1 128.31,120.12
X$28377 430 603 431 644 645 cell_1rw
* cell instance $28378 m0 *1 128.31,122.85
X$28378 430 604 431 644 645 cell_1rw
* cell instance $28379 r0 *1 128.31,122.85
X$28379 430 605 431 644 645 cell_1rw
* cell instance $28380 m0 *1 128.31,125.58
X$28380 430 606 431 644 645 cell_1rw
* cell instance $28381 r0 *1 128.31,125.58
X$28381 430 607 431 644 645 cell_1rw
* cell instance $28382 m0 *1 128.31,128.31
X$28382 430 609 431 644 645 cell_1rw
* cell instance $28383 r0 *1 128.31,128.31
X$28383 430 608 431 644 645 cell_1rw
* cell instance $28384 m0 *1 128.31,131.04
X$28384 430 610 431 644 645 cell_1rw
* cell instance $28385 r0 *1 128.31,131.04
X$28385 430 611 431 644 645 cell_1rw
* cell instance $28386 m0 *1 128.31,133.77
X$28386 430 612 431 644 645 cell_1rw
* cell instance $28387 r0 *1 128.31,133.77
X$28387 430 613 431 644 645 cell_1rw
* cell instance $28388 m0 *1 128.31,136.5
X$28388 430 615 431 644 645 cell_1rw
* cell instance $28389 m0 *1 128.31,139.23
X$28389 430 617 431 644 645 cell_1rw
* cell instance $28390 r0 *1 128.31,136.5
X$28390 430 614 431 644 645 cell_1rw
* cell instance $28391 r0 *1 128.31,139.23
X$28391 430 616 431 644 645 cell_1rw
* cell instance $28392 m0 *1 128.31,141.96
X$28392 430 618 431 644 645 cell_1rw
* cell instance $28393 r0 *1 128.31,141.96
X$28393 430 619 431 644 645 cell_1rw
* cell instance $28394 m0 *1 128.31,144.69
X$28394 430 620 431 644 645 cell_1rw
* cell instance $28395 r0 *1 128.31,144.69
X$28395 430 621 431 644 645 cell_1rw
* cell instance $28396 m0 *1 128.31,147.42
X$28396 430 622 431 644 645 cell_1rw
* cell instance $28397 r0 *1 128.31,147.42
X$28397 430 623 431 644 645 cell_1rw
* cell instance $28398 m0 *1 128.31,150.15
X$28398 430 624 431 644 645 cell_1rw
* cell instance $28399 m0 *1 128.31,152.88
X$28399 430 626 431 644 645 cell_1rw
* cell instance $28400 r0 *1 128.31,150.15
X$28400 430 625 431 644 645 cell_1rw
* cell instance $28401 r0 *1 128.31,152.88
X$28401 430 627 431 644 645 cell_1rw
* cell instance $28402 m0 *1 128.31,155.61
X$28402 430 628 431 644 645 cell_1rw
* cell instance $28403 r0 *1 128.31,155.61
X$28403 430 629 431 644 645 cell_1rw
* cell instance $28404 m0 *1 128.31,158.34
X$28404 430 630 431 644 645 cell_1rw
* cell instance $28405 r0 *1 128.31,158.34
X$28405 430 631 431 644 645 cell_1rw
* cell instance $28406 m0 *1 128.31,161.07
X$28406 430 632 431 644 645 cell_1rw
* cell instance $28407 r0 *1 128.31,161.07
X$28407 430 633 431 644 645 cell_1rw
* cell instance $28408 m0 *1 128.31,163.8
X$28408 430 634 431 644 645 cell_1rw
* cell instance $28409 r0 *1 128.31,163.8
X$28409 430 635 431 644 645 cell_1rw
* cell instance $28410 m0 *1 128.31,166.53
X$28410 430 637 431 644 645 cell_1rw
* cell instance $28411 r0 *1 128.31,166.53
X$28411 430 636 431 644 645 cell_1rw
* cell instance $28412 m0 *1 128.31,169.26
X$28412 430 639 431 644 645 cell_1rw
* cell instance $28413 r0 *1 128.31,169.26
X$28413 430 638 431 644 645 cell_1rw
* cell instance $28414 m0 *1 128.31,171.99
X$28414 430 640 431 644 645 cell_1rw
* cell instance $28415 r0 *1 128.31,171.99
X$28415 430 641 431 644 645 cell_1rw
* cell instance $28416 m0 *1 128.31,174.72
X$28416 430 642 431 644 645 cell_1rw
* cell instance $28417 r0 *1 128.31,174.72
X$28417 430 643 431 644 645 cell_1rw
* cell instance $28418 m0 *1 129.015,90.09
X$28418 432 581 433 644 645 cell_1rw
* cell instance $28419 r0 *1 129.015,90.09
X$28419 432 580 433 644 645 cell_1rw
* cell instance $28420 m0 *1 129.015,92.82
X$28420 432 583 433 644 645 cell_1rw
* cell instance $28421 m0 *1 129.015,95.55
X$28421 432 584 433 644 645 cell_1rw
* cell instance $28422 r0 *1 129.015,92.82
X$28422 432 582 433 644 645 cell_1rw
* cell instance $28423 m0 *1 129.015,98.28
X$28423 432 586 433 644 645 cell_1rw
* cell instance $28424 r0 *1 129.015,95.55
X$28424 432 585 433 644 645 cell_1rw
* cell instance $28425 r0 *1 129.015,98.28
X$28425 432 587 433 644 645 cell_1rw
* cell instance $28426 m0 *1 129.015,101.01
X$28426 432 588 433 644 645 cell_1rw
* cell instance $28427 r0 *1 129.015,101.01
X$28427 432 589 433 644 645 cell_1rw
* cell instance $28428 m0 *1 129.015,103.74
X$28428 432 590 433 644 645 cell_1rw
* cell instance $28429 r0 *1 129.015,103.74
X$28429 432 591 433 644 645 cell_1rw
* cell instance $28430 m0 *1 129.015,106.47
X$28430 432 593 433 644 645 cell_1rw
* cell instance $28431 r0 *1 129.015,106.47
X$28431 432 592 433 644 645 cell_1rw
* cell instance $28432 m0 *1 129.015,109.2
X$28432 432 594 433 644 645 cell_1rw
* cell instance $28433 r0 *1 129.015,109.2
X$28433 432 595 433 644 645 cell_1rw
* cell instance $28434 m0 *1 129.015,111.93
X$28434 432 597 433 644 645 cell_1rw
* cell instance $28435 r0 *1 129.015,111.93
X$28435 432 596 433 644 645 cell_1rw
* cell instance $28436 m0 *1 129.015,114.66
X$28436 432 598 433 644 645 cell_1rw
* cell instance $28437 r0 *1 129.015,114.66
X$28437 432 599 433 644 645 cell_1rw
* cell instance $28438 m0 *1 129.015,117.39
X$28438 432 600 433 644 645 cell_1rw
* cell instance $28439 r0 *1 129.015,117.39
X$28439 432 601 433 644 645 cell_1rw
* cell instance $28440 m0 *1 129.015,120.12
X$28440 432 602 433 644 645 cell_1rw
* cell instance $28441 r0 *1 129.015,120.12
X$28441 432 603 433 644 645 cell_1rw
* cell instance $28442 m0 *1 129.015,122.85
X$28442 432 604 433 644 645 cell_1rw
* cell instance $28443 m0 *1 129.015,125.58
X$28443 432 606 433 644 645 cell_1rw
* cell instance $28444 r0 *1 129.015,122.85
X$28444 432 605 433 644 645 cell_1rw
* cell instance $28445 r0 *1 129.015,125.58
X$28445 432 607 433 644 645 cell_1rw
* cell instance $28446 m0 *1 129.015,128.31
X$28446 432 609 433 644 645 cell_1rw
* cell instance $28447 r0 *1 129.015,128.31
X$28447 432 608 433 644 645 cell_1rw
* cell instance $28448 m0 *1 129.015,131.04
X$28448 432 610 433 644 645 cell_1rw
* cell instance $28449 r0 *1 129.015,131.04
X$28449 432 611 433 644 645 cell_1rw
* cell instance $28450 m0 *1 129.015,133.77
X$28450 432 612 433 644 645 cell_1rw
* cell instance $28451 r0 *1 129.015,133.77
X$28451 432 613 433 644 645 cell_1rw
* cell instance $28452 m0 *1 129.015,136.5
X$28452 432 615 433 644 645 cell_1rw
* cell instance $28453 r0 *1 129.015,136.5
X$28453 432 614 433 644 645 cell_1rw
* cell instance $28454 m0 *1 129.015,139.23
X$28454 432 617 433 644 645 cell_1rw
* cell instance $28455 r0 *1 129.015,139.23
X$28455 432 616 433 644 645 cell_1rw
* cell instance $28456 m0 *1 129.015,141.96
X$28456 432 618 433 644 645 cell_1rw
* cell instance $28457 r0 *1 129.015,141.96
X$28457 432 619 433 644 645 cell_1rw
* cell instance $28458 m0 *1 129.015,144.69
X$28458 432 620 433 644 645 cell_1rw
* cell instance $28459 r0 *1 129.015,144.69
X$28459 432 621 433 644 645 cell_1rw
* cell instance $28460 m0 *1 129.015,147.42
X$28460 432 622 433 644 645 cell_1rw
* cell instance $28461 r0 *1 129.015,147.42
X$28461 432 623 433 644 645 cell_1rw
* cell instance $28462 m0 *1 129.015,150.15
X$28462 432 624 433 644 645 cell_1rw
* cell instance $28463 r0 *1 129.015,150.15
X$28463 432 625 433 644 645 cell_1rw
* cell instance $28464 m0 *1 129.015,152.88
X$28464 432 626 433 644 645 cell_1rw
* cell instance $28465 r0 *1 129.015,152.88
X$28465 432 627 433 644 645 cell_1rw
* cell instance $28466 m0 *1 129.015,155.61
X$28466 432 628 433 644 645 cell_1rw
* cell instance $28467 r0 *1 129.015,155.61
X$28467 432 629 433 644 645 cell_1rw
* cell instance $28468 m0 *1 129.015,158.34
X$28468 432 630 433 644 645 cell_1rw
* cell instance $28469 r0 *1 129.015,158.34
X$28469 432 631 433 644 645 cell_1rw
* cell instance $28470 m0 *1 129.015,161.07
X$28470 432 632 433 644 645 cell_1rw
* cell instance $28471 m0 *1 129.015,163.8
X$28471 432 634 433 644 645 cell_1rw
* cell instance $28472 r0 *1 129.015,161.07
X$28472 432 633 433 644 645 cell_1rw
* cell instance $28473 r0 *1 129.015,163.8
X$28473 432 635 433 644 645 cell_1rw
* cell instance $28474 m0 *1 129.015,166.53
X$28474 432 637 433 644 645 cell_1rw
* cell instance $28475 r0 *1 129.015,166.53
X$28475 432 636 433 644 645 cell_1rw
* cell instance $28476 m0 *1 129.015,169.26
X$28476 432 639 433 644 645 cell_1rw
* cell instance $28477 r0 *1 129.015,169.26
X$28477 432 638 433 644 645 cell_1rw
* cell instance $28478 m0 *1 129.015,171.99
X$28478 432 640 433 644 645 cell_1rw
* cell instance $28479 r0 *1 129.015,171.99
X$28479 432 641 433 644 645 cell_1rw
* cell instance $28480 m0 *1 129.015,174.72
X$28480 432 642 433 644 645 cell_1rw
* cell instance $28481 r0 *1 129.015,174.72
X$28481 432 643 433 644 645 cell_1rw
* cell instance $28482 m0 *1 129.72,90.09
X$28482 434 581 435 644 645 cell_1rw
* cell instance $28483 r0 *1 129.72,90.09
X$28483 434 580 435 644 645 cell_1rw
* cell instance $28484 m0 *1 129.72,92.82
X$28484 434 583 435 644 645 cell_1rw
* cell instance $28485 r0 *1 129.72,92.82
X$28485 434 582 435 644 645 cell_1rw
* cell instance $28486 m0 *1 129.72,95.55
X$28486 434 584 435 644 645 cell_1rw
* cell instance $28487 r0 *1 129.72,95.55
X$28487 434 585 435 644 645 cell_1rw
* cell instance $28488 m0 *1 129.72,98.28
X$28488 434 586 435 644 645 cell_1rw
* cell instance $28489 r0 *1 129.72,98.28
X$28489 434 587 435 644 645 cell_1rw
* cell instance $28490 m0 *1 129.72,101.01
X$28490 434 588 435 644 645 cell_1rw
* cell instance $28491 r0 *1 129.72,101.01
X$28491 434 589 435 644 645 cell_1rw
* cell instance $28492 m0 *1 129.72,103.74
X$28492 434 590 435 644 645 cell_1rw
* cell instance $28493 r0 *1 129.72,103.74
X$28493 434 591 435 644 645 cell_1rw
* cell instance $28494 m0 *1 129.72,106.47
X$28494 434 593 435 644 645 cell_1rw
* cell instance $28495 r0 *1 129.72,106.47
X$28495 434 592 435 644 645 cell_1rw
* cell instance $28496 m0 *1 129.72,109.2
X$28496 434 594 435 644 645 cell_1rw
* cell instance $28497 m0 *1 129.72,111.93
X$28497 434 597 435 644 645 cell_1rw
* cell instance $28498 r0 *1 129.72,109.2
X$28498 434 595 435 644 645 cell_1rw
* cell instance $28499 r0 *1 129.72,111.93
X$28499 434 596 435 644 645 cell_1rw
* cell instance $28500 m0 *1 129.72,114.66
X$28500 434 598 435 644 645 cell_1rw
* cell instance $28501 r0 *1 129.72,114.66
X$28501 434 599 435 644 645 cell_1rw
* cell instance $28502 m0 *1 129.72,117.39
X$28502 434 600 435 644 645 cell_1rw
* cell instance $28503 r0 *1 129.72,117.39
X$28503 434 601 435 644 645 cell_1rw
* cell instance $28504 m0 *1 129.72,120.12
X$28504 434 602 435 644 645 cell_1rw
* cell instance $28505 r0 *1 129.72,120.12
X$28505 434 603 435 644 645 cell_1rw
* cell instance $28506 m0 *1 129.72,122.85
X$28506 434 604 435 644 645 cell_1rw
* cell instance $28507 r0 *1 129.72,122.85
X$28507 434 605 435 644 645 cell_1rw
* cell instance $28508 m0 *1 129.72,125.58
X$28508 434 606 435 644 645 cell_1rw
* cell instance $28509 r0 *1 129.72,125.58
X$28509 434 607 435 644 645 cell_1rw
* cell instance $28510 m0 *1 129.72,128.31
X$28510 434 609 435 644 645 cell_1rw
* cell instance $28511 m0 *1 129.72,131.04
X$28511 434 610 435 644 645 cell_1rw
* cell instance $28512 r0 *1 129.72,128.31
X$28512 434 608 435 644 645 cell_1rw
* cell instance $28513 r0 *1 129.72,131.04
X$28513 434 611 435 644 645 cell_1rw
* cell instance $28514 m0 *1 129.72,133.77
X$28514 434 612 435 644 645 cell_1rw
* cell instance $28515 r0 *1 129.72,133.77
X$28515 434 613 435 644 645 cell_1rw
* cell instance $28516 m0 *1 129.72,136.5
X$28516 434 615 435 644 645 cell_1rw
* cell instance $28517 r0 *1 129.72,136.5
X$28517 434 614 435 644 645 cell_1rw
* cell instance $28518 m0 *1 129.72,139.23
X$28518 434 617 435 644 645 cell_1rw
* cell instance $28519 r0 *1 129.72,139.23
X$28519 434 616 435 644 645 cell_1rw
* cell instance $28520 m0 *1 129.72,141.96
X$28520 434 618 435 644 645 cell_1rw
* cell instance $28521 r0 *1 129.72,141.96
X$28521 434 619 435 644 645 cell_1rw
* cell instance $28522 m0 *1 129.72,144.69
X$28522 434 620 435 644 645 cell_1rw
* cell instance $28523 r0 *1 129.72,144.69
X$28523 434 621 435 644 645 cell_1rw
* cell instance $28524 m0 *1 129.72,147.42
X$28524 434 622 435 644 645 cell_1rw
* cell instance $28525 m0 *1 129.72,150.15
X$28525 434 624 435 644 645 cell_1rw
* cell instance $28526 r0 *1 129.72,147.42
X$28526 434 623 435 644 645 cell_1rw
* cell instance $28527 r0 *1 129.72,150.15
X$28527 434 625 435 644 645 cell_1rw
* cell instance $28528 m0 *1 129.72,152.88
X$28528 434 626 435 644 645 cell_1rw
* cell instance $28529 m0 *1 129.72,155.61
X$28529 434 628 435 644 645 cell_1rw
* cell instance $28530 r0 *1 129.72,152.88
X$28530 434 627 435 644 645 cell_1rw
* cell instance $28531 r0 *1 129.72,155.61
X$28531 434 629 435 644 645 cell_1rw
* cell instance $28532 m0 *1 129.72,158.34
X$28532 434 630 435 644 645 cell_1rw
* cell instance $28533 m0 *1 129.72,161.07
X$28533 434 632 435 644 645 cell_1rw
* cell instance $28534 r0 *1 129.72,158.34
X$28534 434 631 435 644 645 cell_1rw
* cell instance $28535 r0 *1 129.72,161.07
X$28535 434 633 435 644 645 cell_1rw
* cell instance $28536 m0 *1 129.72,163.8
X$28536 434 634 435 644 645 cell_1rw
* cell instance $28537 r0 *1 129.72,163.8
X$28537 434 635 435 644 645 cell_1rw
* cell instance $28538 m0 *1 129.72,166.53
X$28538 434 637 435 644 645 cell_1rw
* cell instance $28539 r0 *1 129.72,166.53
X$28539 434 636 435 644 645 cell_1rw
* cell instance $28540 m0 *1 129.72,169.26
X$28540 434 639 435 644 645 cell_1rw
* cell instance $28541 m0 *1 129.72,171.99
X$28541 434 640 435 644 645 cell_1rw
* cell instance $28542 r0 *1 129.72,169.26
X$28542 434 638 435 644 645 cell_1rw
* cell instance $28543 m0 *1 129.72,174.72
X$28543 434 642 435 644 645 cell_1rw
* cell instance $28544 r0 *1 129.72,171.99
X$28544 434 641 435 644 645 cell_1rw
* cell instance $28545 r0 *1 129.72,174.72
X$28545 434 643 435 644 645 cell_1rw
* cell instance $28546 m0 *1 130.425,90.09
X$28546 436 581 437 644 645 cell_1rw
* cell instance $28547 r0 *1 130.425,90.09
X$28547 436 580 437 644 645 cell_1rw
* cell instance $28548 m0 *1 130.425,92.82
X$28548 436 583 437 644 645 cell_1rw
* cell instance $28549 m0 *1 130.425,95.55
X$28549 436 584 437 644 645 cell_1rw
* cell instance $28550 r0 *1 130.425,92.82
X$28550 436 582 437 644 645 cell_1rw
* cell instance $28551 m0 *1 130.425,98.28
X$28551 436 586 437 644 645 cell_1rw
* cell instance $28552 r0 *1 130.425,95.55
X$28552 436 585 437 644 645 cell_1rw
* cell instance $28553 r0 *1 130.425,98.28
X$28553 436 587 437 644 645 cell_1rw
* cell instance $28554 m0 *1 130.425,101.01
X$28554 436 588 437 644 645 cell_1rw
* cell instance $28555 r0 *1 130.425,101.01
X$28555 436 589 437 644 645 cell_1rw
* cell instance $28556 m0 *1 130.425,103.74
X$28556 436 590 437 644 645 cell_1rw
* cell instance $28557 r0 *1 130.425,103.74
X$28557 436 591 437 644 645 cell_1rw
* cell instance $28558 m0 *1 130.425,106.47
X$28558 436 593 437 644 645 cell_1rw
* cell instance $28559 r0 *1 130.425,106.47
X$28559 436 592 437 644 645 cell_1rw
* cell instance $28560 m0 *1 130.425,109.2
X$28560 436 594 437 644 645 cell_1rw
* cell instance $28561 r0 *1 130.425,109.2
X$28561 436 595 437 644 645 cell_1rw
* cell instance $28562 m0 *1 130.425,111.93
X$28562 436 597 437 644 645 cell_1rw
* cell instance $28563 r0 *1 130.425,111.93
X$28563 436 596 437 644 645 cell_1rw
* cell instance $28564 m0 *1 130.425,114.66
X$28564 436 598 437 644 645 cell_1rw
* cell instance $28565 m0 *1 130.425,117.39
X$28565 436 600 437 644 645 cell_1rw
* cell instance $28566 r0 *1 130.425,114.66
X$28566 436 599 437 644 645 cell_1rw
* cell instance $28567 r0 *1 130.425,117.39
X$28567 436 601 437 644 645 cell_1rw
* cell instance $28568 m0 *1 130.425,120.12
X$28568 436 602 437 644 645 cell_1rw
* cell instance $28569 r0 *1 130.425,120.12
X$28569 436 603 437 644 645 cell_1rw
* cell instance $28570 m0 *1 130.425,122.85
X$28570 436 604 437 644 645 cell_1rw
* cell instance $28571 r0 *1 130.425,122.85
X$28571 436 605 437 644 645 cell_1rw
* cell instance $28572 m0 *1 130.425,125.58
X$28572 436 606 437 644 645 cell_1rw
* cell instance $28573 r0 *1 130.425,125.58
X$28573 436 607 437 644 645 cell_1rw
* cell instance $28574 m0 *1 130.425,128.31
X$28574 436 609 437 644 645 cell_1rw
* cell instance $28575 r0 *1 130.425,128.31
X$28575 436 608 437 644 645 cell_1rw
* cell instance $28576 m0 *1 130.425,131.04
X$28576 436 610 437 644 645 cell_1rw
* cell instance $28577 r0 *1 130.425,131.04
X$28577 436 611 437 644 645 cell_1rw
* cell instance $28578 m0 *1 130.425,133.77
X$28578 436 612 437 644 645 cell_1rw
* cell instance $28579 r0 *1 130.425,133.77
X$28579 436 613 437 644 645 cell_1rw
* cell instance $28580 m0 *1 130.425,136.5
X$28580 436 615 437 644 645 cell_1rw
* cell instance $28581 m0 *1 130.425,139.23
X$28581 436 617 437 644 645 cell_1rw
* cell instance $28582 r0 *1 130.425,136.5
X$28582 436 614 437 644 645 cell_1rw
* cell instance $28583 r0 *1 130.425,139.23
X$28583 436 616 437 644 645 cell_1rw
* cell instance $28584 m0 *1 130.425,141.96
X$28584 436 618 437 644 645 cell_1rw
* cell instance $28585 r0 *1 130.425,141.96
X$28585 436 619 437 644 645 cell_1rw
* cell instance $28586 m0 *1 130.425,144.69
X$28586 436 620 437 644 645 cell_1rw
* cell instance $28587 r0 *1 130.425,144.69
X$28587 436 621 437 644 645 cell_1rw
* cell instance $28588 m0 *1 130.425,147.42
X$28588 436 622 437 644 645 cell_1rw
* cell instance $28589 r0 *1 130.425,147.42
X$28589 436 623 437 644 645 cell_1rw
* cell instance $28590 m0 *1 130.425,150.15
X$28590 436 624 437 644 645 cell_1rw
* cell instance $28591 m0 *1 130.425,152.88
X$28591 436 626 437 644 645 cell_1rw
* cell instance $28592 r0 *1 130.425,150.15
X$28592 436 625 437 644 645 cell_1rw
* cell instance $28593 r0 *1 130.425,152.88
X$28593 436 627 437 644 645 cell_1rw
* cell instance $28594 m0 *1 130.425,155.61
X$28594 436 628 437 644 645 cell_1rw
* cell instance $28595 r0 *1 130.425,155.61
X$28595 436 629 437 644 645 cell_1rw
* cell instance $28596 m0 *1 130.425,158.34
X$28596 436 630 437 644 645 cell_1rw
* cell instance $28597 r0 *1 130.425,158.34
X$28597 436 631 437 644 645 cell_1rw
* cell instance $28598 m0 *1 130.425,161.07
X$28598 436 632 437 644 645 cell_1rw
* cell instance $28599 r0 *1 130.425,161.07
X$28599 436 633 437 644 645 cell_1rw
* cell instance $28600 m0 *1 130.425,163.8
X$28600 436 634 437 644 645 cell_1rw
* cell instance $28601 r0 *1 130.425,163.8
X$28601 436 635 437 644 645 cell_1rw
* cell instance $28602 m0 *1 130.425,166.53
X$28602 436 637 437 644 645 cell_1rw
* cell instance $28603 r0 *1 130.425,166.53
X$28603 436 636 437 644 645 cell_1rw
* cell instance $28604 m0 *1 130.425,169.26
X$28604 436 639 437 644 645 cell_1rw
* cell instance $28605 r0 *1 130.425,169.26
X$28605 436 638 437 644 645 cell_1rw
* cell instance $28606 m0 *1 130.425,171.99
X$28606 436 640 437 644 645 cell_1rw
* cell instance $28607 r0 *1 130.425,171.99
X$28607 436 641 437 644 645 cell_1rw
* cell instance $28608 m0 *1 130.425,174.72
X$28608 436 642 437 644 645 cell_1rw
* cell instance $28609 r0 *1 130.425,174.72
X$28609 436 643 437 644 645 cell_1rw
* cell instance $28610 m0 *1 131.13,90.09
X$28610 438 581 439 644 645 cell_1rw
* cell instance $28611 m0 *1 131.13,92.82
X$28611 438 583 439 644 645 cell_1rw
* cell instance $28612 r0 *1 131.13,90.09
X$28612 438 580 439 644 645 cell_1rw
* cell instance $28613 r0 *1 131.13,92.82
X$28613 438 582 439 644 645 cell_1rw
* cell instance $28614 m0 *1 131.13,95.55
X$28614 438 584 439 644 645 cell_1rw
* cell instance $28615 m0 *1 131.13,98.28
X$28615 438 586 439 644 645 cell_1rw
* cell instance $28616 r0 *1 131.13,95.55
X$28616 438 585 439 644 645 cell_1rw
* cell instance $28617 r0 *1 131.13,98.28
X$28617 438 587 439 644 645 cell_1rw
* cell instance $28618 m0 *1 131.13,101.01
X$28618 438 588 439 644 645 cell_1rw
* cell instance $28619 r0 *1 131.13,101.01
X$28619 438 589 439 644 645 cell_1rw
* cell instance $28620 m0 *1 131.13,103.74
X$28620 438 590 439 644 645 cell_1rw
* cell instance $28621 m0 *1 131.13,106.47
X$28621 438 593 439 644 645 cell_1rw
* cell instance $28622 r0 *1 131.13,103.74
X$28622 438 591 439 644 645 cell_1rw
* cell instance $28623 r0 *1 131.13,106.47
X$28623 438 592 439 644 645 cell_1rw
* cell instance $28624 m0 *1 131.13,109.2
X$28624 438 594 439 644 645 cell_1rw
* cell instance $28625 r0 *1 131.13,109.2
X$28625 438 595 439 644 645 cell_1rw
* cell instance $28626 m0 *1 131.13,111.93
X$28626 438 597 439 644 645 cell_1rw
* cell instance $28627 r0 *1 131.13,111.93
X$28627 438 596 439 644 645 cell_1rw
* cell instance $28628 m0 *1 131.13,114.66
X$28628 438 598 439 644 645 cell_1rw
* cell instance $28629 m0 *1 131.13,117.39
X$28629 438 600 439 644 645 cell_1rw
* cell instance $28630 r0 *1 131.13,114.66
X$28630 438 599 439 644 645 cell_1rw
* cell instance $28631 r0 *1 131.13,117.39
X$28631 438 601 439 644 645 cell_1rw
* cell instance $28632 m0 *1 131.13,120.12
X$28632 438 602 439 644 645 cell_1rw
* cell instance $28633 r0 *1 131.13,120.12
X$28633 438 603 439 644 645 cell_1rw
* cell instance $28634 m0 *1 131.13,122.85
X$28634 438 604 439 644 645 cell_1rw
* cell instance $28635 r0 *1 131.13,122.85
X$28635 438 605 439 644 645 cell_1rw
* cell instance $28636 m0 *1 131.13,125.58
X$28636 438 606 439 644 645 cell_1rw
* cell instance $28637 r0 *1 131.13,125.58
X$28637 438 607 439 644 645 cell_1rw
* cell instance $28638 m0 *1 131.13,128.31
X$28638 438 609 439 644 645 cell_1rw
* cell instance $28639 m0 *1 131.13,131.04
X$28639 438 610 439 644 645 cell_1rw
* cell instance $28640 r0 *1 131.13,128.31
X$28640 438 608 439 644 645 cell_1rw
* cell instance $28641 r0 *1 131.13,131.04
X$28641 438 611 439 644 645 cell_1rw
* cell instance $28642 m0 *1 131.13,133.77
X$28642 438 612 439 644 645 cell_1rw
* cell instance $28643 r0 *1 131.13,133.77
X$28643 438 613 439 644 645 cell_1rw
* cell instance $28644 m0 *1 131.13,136.5
X$28644 438 615 439 644 645 cell_1rw
* cell instance $28645 m0 *1 131.13,139.23
X$28645 438 617 439 644 645 cell_1rw
* cell instance $28646 r0 *1 131.13,136.5
X$28646 438 614 439 644 645 cell_1rw
* cell instance $28647 m0 *1 131.13,141.96
X$28647 438 618 439 644 645 cell_1rw
* cell instance $28648 r0 *1 131.13,139.23
X$28648 438 616 439 644 645 cell_1rw
* cell instance $28649 r0 *1 131.13,141.96
X$28649 438 619 439 644 645 cell_1rw
* cell instance $28650 m0 *1 131.13,144.69
X$28650 438 620 439 644 645 cell_1rw
* cell instance $28651 r0 *1 131.13,144.69
X$28651 438 621 439 644 645 cell_1rw
* cell instance $28652 m0 *1 131.13,147.42
X$28652 438 622 439 644 645 cell_1rw
* cell instance $28653 r0 *1 131.13,147.42
X$28653 438 623 439 644 645 cell_1rw
* cell instance $28654 m0 *1 131.13,150.15
X$28654 438 624 439 644 645 cell_1rw
* cell instance $28655 r0 *1 131.13,150.15
X$28655 438 625 439 644 645 cell_1rw
* cell instance $28656 m0 *1 131.13,152.88
X$28656 438 626 439 644 645 cell_1rw
* cell instance $28657 r0 *1 131.13,152.88
X$28657 438 627 439 644 645 cell_1rw
* cell instance $28658 m0 *1 131.13,155.61
X$28658 438 628 439 644 645 cell_1rw
* cell instance $28659 r0 *1 131.13,155.61
X$28659 438 629 439 644 645 cell_1rw
* cell instance $28660 m0 *1 131.13,158.34
X$28660 438 630 439 644 645 cell_1rw
* cell instance $28661 r0 *1 131.13,158.34
X$28661 438 631 439 644 645 cell_1rw
* cell instance $28662 m0 *1 131.13,161.07
X$28662 438 632 439 644 645 cell_1rw
* cell instance $28663 r0 *1 131.13,161.07
X$28663 438 633 439 644 645 cell_1rw
* cell instance $28664 m0 *1 131.13,163.8
X$28664 438 634 439 644 645 cell_1rw
* cell instance $28665 r0 *1 131.13,163.8
X$28665 438 635 439 644 645 cell_1rw
* cell instance $28666 m0 *1 131.13,166.53
X$28666 438 637 439 644 645 cell_1rw
* cell instance $28667 r0 *1 131.13,166.53
X$28667 438 636 439 644 645 cell_1rw
* cell instance $28668 m0 *1 131.13,169.26
X$28668 438 639 439 644 645 cell_1rw
* cell instance $28669 r0 *1 131.13,169.26
X$28669 438 638 439 644 645 cell_1rw
* cell instance $28670 m0 *1 131.13,171.99
X$28670 438 640 439 644 645 cell_1rw
* cell instance $28671 r0 *1 131.13,171.99
X$28671 438 641 439 644 645 cell_1rw
* cell instance $28672 m0 *1 131.13,174.72
X$28672 438 642 439 644 645 cell_1rw
* cell instance $28673 r0 *1 131.13,174.72
X$28673 438 643 439 644 645 cell_1rw
* cell instance $28674 m0 *1 131.835,90.09
X$28674 440 581 441 644 645 cell_1rw
* cell instance $28675 r0 *1 131.835,90.09
X$28675 440 580 441 644 645 cell_1rw
* cell instance $28676 m0 *1 131.835,92.82
X$28676 440 583 441 644 645 cell_1rw
* cell instance $28677 m0 *1 131.835,95.55
X$28677 440 584 441 644 645 cell_1rw
* cell instance $28678 r0 *1 131.835,92.82
X$28678 440 582 441 644 645 cell_1rw
* cell instance $28679 r0 *1 131.835,95.55
X$28679 440 585 441 644 645 cell_1rw
* cell instance $28680 m0 *1 131.835,98.28
X$28680 440 586 441 644 645 cell_1rw
* cell instance $28681 m0 *1 131.835,101.01
X$28681 440 588 441 644 645 cell_1rw
* cell instance $28682 r0 *1 131.835,98.28
X$28682 440 587 441 644 645 cell_1rw
* cell instance $28683 r0 *1 131.835,101.01
X$28683 440 589 441 644 645 cell_1rw
* cell instance $28684 m0 *1 131.835,103.74
X$28684 440 590 441 644 645 cell_1rw
* cell instance $28685 r0 *1 131.835,103.74
X$28685 440 591 441 644 645 cell_1rw
* cell instance $28686 m0 *1 131.835,106.47
X$28686 440 593 441 644 645 cell_1rw
* cell instance $28687 m0 *1 131.835,109.2
X$28687 440 594 441 644 645 cell_1rw
* cell instance $28688 r0 *1 131.835,106.47
X$28688 440 592 441 644 645 cell_1rw
* cell instance $28689 r0 *1 131.835,109.2
X$28689 440 595 441 644 645 cell_1rw
* cell instance $28690 m0 *1 131.835,111.93
X$28690 440 597 441 644 645 cell_1rw
* cell instance $28691 r0 *1 131.835,111.93
X$28691 440 596 441 644 645 cell_1rw
* cell instance $28692 m0 *1 131.835,114.66
X$28692 440 598 441 644 645 cell_1rw
* cell instance $28693 r0 *1 131.835,114.66
X$28693 440 599 441 644 645 cell_1rw
* cell instance $28694 m0 *1 131.835,117.39
X$28694 440 600 441 644 645 cell_1rw
* cell instance $28695 r0 *1 131.835,117.39
X$28695 440 601 441 644 645 cell_1rw
* cell instance $28696 m0 *1 131.835,120.12
X$28696 440 602 441 644 645 cell_1rw
* cell instance $28697 m0 *1 131.835,122.85
X$28697 440 604 441 644 645 cell_1rw
* cell instance $28698 r0 *1 131.835,120.12
X$28698 440 603 441 644 645 cell_1rw
* cell instance $28699 r0 *1 131.835,122.85
X$28699 440 605 441 644 645 cell_1rw
* cell instance $28700 m0 *1 131.835,125.58
X$28700 440 606 441 644 645 cell_1rw
* cell instance $28701 r0 *1 131.835,125.58
X$28701 440 607 441 644 645 cell_1rw
* cell instance $28702 m0 *1 131.835,128.31
X$28702 440 609 441 644 645 cell_1rw
* cell instance $28703 r0 *1 131.835,128.31
X$28703 440 608 441 644 645 cell_1rw
* cell instance $28704 m0 *1 131.835,131.04
X$28704 440 610 441 644 645 cell_1rw
* cell instance $28705 r0 *1 131.835,131.04
X$28705 440 611 441 644 645 cell_1rw
* cell instance $28706 m0 *1 131.835,133.77
X$28706 440 612 441 644 645 cell_1rw
* cell instance $28707 m0 *1 131.835,136.5
X$28707 440 615 441 644 645 cell_1rw
* cell instance $28708 r0 *1 131.835,133.77
X$28708 440 613 441 644 645 cell_1rw
* cell instance $28709 m0 *1 131.835,139.23
X$28709 440 617 441 644 645 cell_1rw
* cell instance $28710 r0 *1 131.835,136.5
X$28710 440 614 441 644 645 cell_1rw
* cell instance $28711 r0 *1 131.835,139.23
X$28711 440 616 441 644 645 cell_1rw
* cell instance $28712 m0 *1 131.835,141.96
X$28712 440 618 441 644 645 cell_1rw
* cell instance $28713 m0 *1 131.835,144.69
X$28713 440 620 441 644 645 cell_1rw
* cell instance $28714 r0 *1 131.835,141.96
X$28714 440 619 441 644 645 cell_1rw
* cell instance $28715 r0 *1 131.835,144.69
X$28715 440 621 441 644 645 cell_1rw
* cell instance $28716 m0 *1 131.835,147.42
X$28716 440 622 441 644 645 cell_1rw
* cell instance $28717 m0 *1 131.835,150.15
X$28717 440 624 441 644 645 cell_1rw
* cell instance $28718 r0 *1 131.835,147.42
X$28718 440 623 441 644 645 cell_1rw
* cell instance $28719 r0 *1 131.835,150.15
X$28719 440 625 441 644 645 cell_1rw
* cell instance $28720 m0 *1 131.835,152.88
X$28720 440 626 441 644 645 cell_1rw
* cell instance $28721 r0 *1 131.835,152.88
X$28721 440 627 441 644 645 cell_1rw
* cell instance $28722 m0 *1 131.835,155.61
X$28722 440 628 441 644 645 cell_1rw
* cell instance $28723 r0 *1 131.835,155.61
X$28723 440 629 441 644 645 cell_1rw
* cell instance $28724 m0 *1 131.835,158.34
X$28724 440 630 441 644 645 cell_1rw
* cell instance $28725 r0 *1 131.835,158.34
X$28725 440 631 441 644 645 cell_1rw
* cell instance $28726 m0 *1 131.835,161.07
X$28726 440 632 441 644 645 cell_1rw
* cell instance $28727 r0 *1 131.835,161.07
X$28727 440 633 441 644 645 cell_1rw
* cell instance $28728 m0 *1 131.835,163.8
X$28728 440 634 441 644 645 cell_1rw
* cell instance $28729 r0 *1 131.835,163.8
X$28729 440 635 441 644 645 cell_1rw
* cell instance $28730 m0 *1 131.835,166.53
X$28730 440 637 441 644 645 cell_1rw
* cell instance $28731 m0 *1 131.835,169.26
X$28731 440 639 441 644 645 cell_1rw
* cell instance $28732 r0 *1 131.835,166.53
X$28732 440 636 441 644 645 cell_1rw
* cell instance $28733 r0 *1 131.835,169.26
X$28733 440 638 441 644 645 cell_1rw
* cell instance $28734 m0 *1 131.835,171.99
X$28734 440 640 441 644 645 cell_1rw
* cell instance $28735 m0 *1 131.835,174.72
X$28735 440 642 441 644 645 cell_1rw
* cell instance $28736 r0 *1 131.835,171.99
X$28736 440 641 441 644 645 cell_1rw
* cell instance $28737 r0 *1 131.835,174.72
X$28737 440 643 441 644 645 cell_1rw
* cell instance $28738 m0 *1 132.54,90.09
X$28738 442 581 443 644 645 cell_1rw
* cell instance $28739 r0 *1 132.54,90.09
X$28739 442 580 443 644 645 cell_1rw
* cell instance $28740 m0 *1 132.54,92.82
X$28740 442 583 443 644 645 cell_1rw
* cell instance $28741 r0 *1 132.54,92.82
X$28741 442 582 443 644 645 cell_1rw
* cell instance $28742 m0 *1 132.54,95.55
X$28742 442 584 443 644 645 cell_1rw
* cell instance $28743 r0 *1 132.54,95.55
X$28743 442 585 443 644 645 cell_1rw
* cell instance $28744 m0 *1 132.54,98.28
X$28744 442 586 443 644 645 cell_1rw
* cell instance $28745 r0 *1 132.54,98.28
X$28745 442 587 443 644 645 cell_1rw
* cell instance $28746 m0 *1 132.54,101.01
X$28746 442 588 443 644 645 cell_1rw
* cell instance $28747 r0 *1 132.54,101.01
X$28747 442 589 443 644 645 cell_1rw
* cell instance $28748 m0 *1 132.54,103.74
X$28748 442 590 443 644 645 cell_1rw
* cell instance $28749 r0 *1 132.54,103.74
X$28749 442 591 443 644 645 cell_1rw
* cell instance $28750 m0 *1 132.54,106.47
X$28750 442 593 443 644 645 cell_1rw
* cell instance $28751 m0 *1 132.54,109.2
X$28751 442 594 443 644 645 cell_1rw
* cell instance $28752 r0 *1 132.54,106.47
X$28752 442 592 443 644 645 cell_1rw
* cell instance $28753 r0 *1 132.54,109.2
X$28753 442 595 443 644 645 cell_1rw
* cell instance $28754 m0 *1 132.54,111.93
X$28754 442 597 443 644 645 cell_1rw
* cell instance $28755 m0 *1 132.54,114.66
X$28755 442 598 443 644 645 cell_1rw
* cell instance $28756 r0 *1 132.54,111.93
X$28756 442 596 443 644 645 cell_1rw
* cell instance $28757 r0 *1 132.54,114.66
X$28757 442 599 443 644 645 cell_1rw
* cell instance $28758 m0 *1 132.54,117.39
X$28758 442 600 443 644 645 cell_1rw
* cell instance $28759 r0 *1 132.54,117.39
X$28759 442 601 443 644 645 cell_1rw
* cell instance $28760 m0 *1 132.54,120.12
X$28760 442 602 443 644 645 cell_1rw
* cell instance $28761 r0 *1 132.54,120.12
X$28761 442 603 443 644 645 cell_1rw
* cell instance $28762 m0 *1 132.54,122.85
X$28762 442 604 443 644 645 cell_1rw
* cell instance $28763 r0 *1 132.54,122.85
X$28763 442 605 443 644 645 cell_1rw
* cell instance $28764 m0 *1 132.54,125.58
X$28764 442 606 443 644 645 cell_1rw
* cell instance $28765 r0 *1 132.54,125.58
X$28765 442 607 443 644 645 cell_1rw
* cell instance $28766 m0 *1 132.54,128.31
X$28766 442 609 443 644 645 cell_1rw
* cell instance $28767 r0 *1 132.54,128.31
X$28767 442 608 443 644 645 cell_1rw
* cell instance $28768 m0 *1 132.54,131.04
X$28768 442 610 443 644 645 cell_1rw
* cell instance $28769 r0 *1 132.54,131.04
X$28769 442 611 443 644 645 cell_1rw
* cell instance $28770 m0 *1 132.54,133.77
X$28770 442 612 443 644 645 cell_1rw
* cell instance $28771 r0 *1 132.54,133.77
X$28771 442 613 443 644 645 cell_1rw
* cell instance $28772 m0 *1 132.54,136.5
X$28772 442 615 443 644 645 cell_1rw
* cell instance $28773 m0 *1 132.54,139.23
X$28773 442 617 443 644 645 cell_1rw
* cell instance $28774 r0 *1 132.54,136.5
X$28774 442 614 443 644 645 cell_1rw
* cell instance $28775 m0 *1 132.54,141.96
X$28775 442 618 443 644 645 cell_1rw
* cell instance $28776 r0 *1 132.54,139.23
X$28776 442 616 443 644 645 cell_1rw
* cell instance $28777 r0 *1 132.54,141.96
X$28777 442 619 443 644 645 cell_1rw
* cell instance $28778 m0 *1 132.54,144.69
X$28778 442 620 443 644 645 cell_1rw
* cell instance $28779 r0 *1 132.54,144.69
X$28779 442 621 443 644 645 cell_1rw
* cell instance $28780 m0 *1 132.54,147.42
X$28780 442 622 443 644 645 cell_1rw
* cell instance $28781 r0 *1 132.54,147.42
X$28781 442 623 443 644 645 cell_1rw
* cell instance $28782 m0 *1 132.54,150.15
X$28782 442 624 443 644 645 cell_1rw
* cell instance $28783 m0 *1 132.54,152.88
X$28783 442 626 443 644 645 cell_1rw
* cell instance $28784 r0 *1 132.54,150.15
X$28784 442 625 443 644 645 cell_1rw
* cell instance $28785 m0 *1 132.54,155.61
X$28785 442 628 443 644 645 cell_1rw
* cell instance $28786 r0 *1 132.54,152.88
X$28786 442 627 443 644 645 cell_1rw
* cell instance $28787 r0 *1 132.54,155.61
X$28787 442 629 443 644 645 cell_1rw
* cell instance $28788 m0 *1 132.54,158.34
X$28788 442 630 443 644 645 cell_1rw
* cell instance $28789 r0 *1 132.54,158.34
X$28789 442 631 443 644 645 cell_1rw
* cell instance $28790 m0 *1 132.54,161.07
X$28790 442 632 443 644 645 cell_1rw
* cell instance $28791 r0 *1 132.54,161.07
X$28791 442 633 443 644 645 cell_1rw
* cell instance $28792 m0 *1 132.54,163.8
X$28792 442 634 443 644 645 cell_1rw
* cell instance $28793 r0 *1 132.54,163.8
X$28793 442 635 443 644 645 cell_1rw
* cell instance $28794 m0 *1 132.54,166.53
X$28794 442 637 443 644 645 cell_1rw
* cell instance $28795 r0 *1 132.54,166.53
X$28795 442 636 443 644 645 cell_1rw
* cell instance $28796 m0 *1 132.54,169.26
X$28796 442 639 443 644 645 cell_1rw
* cell instance $28797 r0 *1 132.54,169.26
X$28797 442 638 443 644 645 cell_1rw
* cell instance $28798 m0 *1 132.54,171.99
X$28798 442 640 443 644 645 cell_1rw
* cell instance $28799 r0 *1 132.54,171.99
X$28799 442 641 443 644 645 cell_1rw
* cell instance $28800 m0 *1 132.54,174.72
X$28800 442 642 443 644 645 cell_1rw
* cell instance $28801 r0 *1 132.54,174.72
X$28801 442 643 443 644 645 cell_1rw
* cell instance $28802 m0 *1 133.245,90.09
X$28802 444 581 445 644 645 cell_1rw
* cell instance $28803 r0 *1 133.245,90.09
X$28803 444 580 445 644 645 cell_1rw
* cell instance $28804 m0 *1 133.245,92.82
X$28804 444 583 445 644 645 cell_1rw
* cell instance $28805 m0 *1 133.245,95.55
X$28805 444 584 445 644 645 cell_1rw
* cell instance $28806 r0 *1 133.245,92.82
X$28806 444 582 445 644 645 cell_1rw
* cell instance $28807 r0 *1 133.245,95.55
X$28807 444 585 445 644 645 cell_1rw
* cell instance $28808 m0 *1 133.245,98.28
X$28808 444 586 445 644 645 cell_1rw
* cell instance $28809 r0 *1 133.245,98.28
X$28809 444 587 445 644 645 cell_1rw
* cell instance $28810 m0 *1 133.245,101.01
X$28810 444 588 445 644 645 cell_1rw
* cell instance $28811 r0 *1 133.245,101.01
X$28811 444 589 445 644 645 cell_1rw
* cell instance $28812 m0 *1 133.245,103.74
X$28812 444 590 445 644 645 cell_1rw
* cell instance $28813 r0 *1 133.245,103.74
X$28813 444 591 445 644 645 cell_1rw
* cell instance $28814 m0 *1 133.245,106.47
X$28814 444 593 445 644 645 cell_1rw
* cell instance $28815 m0 *1 133.245,109.2
X$28815 444 594 445 644 645 cell_1rw
* cell instance $28816 r0 *1 133.245,106.47
X$28816 444 592 445 644 645 cell_1rw
* cell instance $28817 r0 *1 133.245,109.2
X$28817 444 595 445 644 645 cell_1rw
* cell instance $28818 m0 *1 133.245,111.93
X$28818 444 597 445 644 645 cell_1rw
* cell instance $28819 m0 *1 133.245,114.66
X$28819 444 598 445 644 645 cell_1rw
* cell instance $28820 r0 *1 133.245,111.93
X$28820 444 596 445 644 645 cell_1rw
* cell instance $28821 r0 *1 133.245,114.66
X$28821 444 599 445 644 645 cell_1rw
* cell instance $28822 m0 *1 133.245,117.39
X$28822 444 600 445 644 645 cell_1rw
* cell instance $28823 m0 *1 133.245,120.12
X$28823 444 602 445 644 645 cell_1rw
* cell instance $28824 r0 *1 133.245,117.39
X$28824 444 601 445 644 645 cell_1rw
* cell instance $28825 r0 *1 133.245,120.12
X$28825 444 603 445 644 645 cell_1rw
* cell instance $28826 m0 *1 133.245,122.85
X$28826 444 604 445 644 645 cell_1rw
* cell instance $28827 r0 *1 133.245,122.85
X$28827 444 605 445 644 645 cell_1rw
* cell instance $28828 m0 *1 133.245,125.58
X$28828 444 606 445 644 645 cell_1rw
* cell instance $28829 r0 *1 133.245,125.58
X$28829 444 607 445 644 645 cell_1rw
* cell instance $28830 m0 *1 133.245,128.31
X$28830 444 609 445 644 645 cell_1rw
* cell instance $28831 r0 *1 133.245,128.31
X$28831 444 608 445 644 645 cell_1rw
* cell instance $28832 m0 *1 133.245,131.04
X$28832 444 610 445 644 645 cell_1rw
* cell instance $28833 r0 *1 133.245,131.04
X$28833 444 611 445 644 645 cell_1rw
* cell instance $28834 m0 *1 133.245,133.77
X$28834 444 612 445 644 645 cell_1rw
* cell instance $28835 r0 *1 133.245,133.77
X$28835 444 613 445 644 645 cell_1rw
* cell instance $28836 m0 *1 133.245,136.5
X$28836 444 615 445 644 645 cell_1rw
* cell instance $28837 r0 *1 133.245,136.5
X$28837 444 614 445 644 645 cell_1rw
* cell instance $28838 m0 *1 133.245,139.23
X$28838 444 617 445 644 645 cell_1rw
* cell instance $28839 r0 *1 133.245,139.23
X$28839 444 616 445 644 645 cell_1rw
* cell instance $28840 m0 *1 133.245,141.96
X$28840 444 618 445 644 645 cell_1rw
* cell instance $28841 r0 *1 133.245,141.96
X$28841 444 619 445 644 645 cell_1rw
* cell instance $28842 m0 *1 133.245,144.69
X$28842 444 620 445 644 645 cell_1rw
* cell instance $28843 r0 *1 133.245,144.69
X$28843 444 621 445 644 645 cell_1rw
* cell instance $28844 m0 *1 133.245,147.42
X$28844 444 622 445 644 645 cell_1rw
* cell instance $28845 r0 *1 133.245,147.42
X$28845 444 623 445 644 645 cell_1rw
* cell instance $28846 m0 *1 133.245,150.15
X$28846 444 624 445 644 645 cell_1rw
* cell instance $28847 r0 *1 133.245,150.15
X$28847 444 625 445 644 645 cell_1rw
* cell instance $28848 m0 *1 133.245,152.88
X$28848 444 626 445 644 645 cell_1rw
* cell instance $28849 r0 *1 133.245,152.88
X$28849 444 627 445 644 645 cell_1rw
* cell instance $28850 m0 *1 133.245,155.61
X$28850 444 628 445 644 645 cell_1rw
* cell instance $28851 r0 *1 133.245,155.61
X$28851 444 629 445 644 645 cell_1rw
* cell instance $28852 m0 *1 133.245,158.34
X$28852 444 630 445 644 645 cell_1rw
* cell instance $28853 m0 *1 133.245,161.07
X$28853 444 632 445 644 645 cell_1rw
* cell instance $28854 r0 *1 133.245,158.34
X$28854 444 631 445 644 645 cell_1rw
* cell instance $28855 m0 *1 133.245,163.8
X$28855 444 634 445 644 645 cell_1rw
* cell instance $28856 r0 *1 133.245,161.07
X$28856 444 633 445 644 645 cell_1rw
* cell instance $28857 r0 *1 133.245,163.8
X$28857 444 635 445 644 645 cell_1rw
* cell instance $28858 m0 *1 133.245,166.53
X$28858 444 637 445 644 645 cell_1rw
* cell instance $28859 m0 *1 133.245,169.26
X$28859 444 639 445 644 645 cell_1rw
* cell instance $28860 r0 *1 133.245,166.53
X$28860 444 636 445 644 645 cell_1rw
* cell instance $28861 r0 *1 133.245,169.26
X$28861 444 638 445 644 645 cell_1rw
* cell instance $28862 m0 *1 133.245,171.99
X$28862 444 640 445 644 645 cell_1rw
* cell instance $28863 r0 *1 133.245,171.99
X$28863 444 641 445 644 645 cell_1rw
* cell instance $28864 m0 *1 133.245,174.72
X$28864 444 642 445 644 645 cell_1rw
* cell instance $28865 r0 *1 133.245,174.72
X$28865 444 643 445 644 645 cell_1rw
* cell instance $28866 m0 *1 133.95,90.09
X$28866 446 581 447 644 645 cell_1rw
* cell instance $28867 r0 *1 133.95,90.09
X$28867 446 580 447 644 645 cell_1rw
* cell instance $28868 m0 *1 133.95,92.82
X$28868 446 583 447 644 645 cell_1rw
* cell instance $28869 r0 *1 133.95,92.82
X$28869 446 582 447 644 645 cell_1rw
* cell instance $28870 m0 *1 133.95,95.55
X$28870 446 584 447 644 645 cell_1rw
* cell instance $28871 r0 *1 133.95,95.55
X$28871 446 585 447 644 645 cell_1rw
* cell instance $28872 m0 *1 133.95,98.28
X$28872 446 586 447 644 645 cell_1rw
* cell instance $28873 r0 *1 133.95,98.28
X$28873 446 587 447 644 645 cell_1rw
* cell instance $28874 m0 *1 133.95,101.01
X$28874 446 588 447 644 645 cell_1rw
* cell instance $28875 r0 *1 133.95,101.01
X$28875 446 589 447 644 645 cell_1rw
* cell instance $28876 m0 *1 133.95,103.74
X$28876 446 590 447 644 645 cell_1rw
* cell instance $28877 m0 *1 133.95,106.47
X$28877 446 593 447 644 645 cell_1rw
* cell instance $28878 r0 *1 133.95,103.74
X$28878 446 591 447 644 645 cell_1rw
* cell instance $28879 r0 *1 133.95,106.47
X$28879 446 592 447 644 645 cell_1rw
* cell instance $28880 m0 *1 133.95,109.2
X$28880 446 594 447 644 645 cell_1rw
* cell instance $28881 r0 *1 133.95,109.2
X$28881 446 595 447 644 645 cell_1rw
* cell instance $28882 m0 *1 133.95,111.93
X$28882 446 597 447 644 645 cell_1rw
* cell instance $28883 m0 *1 133.95,114.66
X$28883 446 598 447 644 645 cell_1rw
* cell instance $28884 r0 *1 133.95,111.93
X$28884 446 596 447 644 645 cell_1rw
* cell instance $28885 r0 *1 133.95,114.66
X$28885 446 599 447 644 645 cell_1rw
* cell instance $28886 m0 *1 133.95,117.39
X$28886 446 600 447 644 645 cell_1rw
* cell instance $28887 r0 *1 133.95,117.39
X$28887 446 601 447 644 645 cell_1rw
* cell instance $28888 m0 *1 133.95,120.12
X$28888 446 602 447 644 645 cell_1rw
* cell instance $28889 r0 *1 133.95,120.12
X$28889 446 603 447 644 645 cell_1rw
* cell instance $28890 m0 *1 133.95,122.85
X$28890 446 604 447 644 645 cell_1rw
* cell instance $28891 r0 *1 133.95,122.85
X$28891 446 605 447 644 645 cell_1rw
* cell instance $28892 m0 *1 133.95,125.58
X$28892 446 606 447 644 645 cell_1rw
* cell instance $28893 r0 *1 133.95,125.58
X$28893 446 607 447 644 645 cell_1rw
* cell instance $28894 m0 *1 133.95,128.31
X$28894 446 609 447 644 645 cell_1rw
* cell instance $28895 r0 *1 133.95,128.31
X$28895 446 608 447 644 645 cell_1rw
* cell instance $28896 m0 *1 133.95,131.04
X$28896 446 610 447 644 645 cell_1rw
* cell instance $28897 r0 *1 133.95,131.04
X$28897 446 611 447 644 645 cell_1rw
* cell instance $28898 m0 *1 133.95,133.77
X$28898 446 612 447 644 645 cell_1rw
* cell instance $28899 r0 *1 133.95,133.77
X$28899 446 613 447 644 645 cell_1rw
* cell instance $28900 m0 *1 133.95,136.5
X$28900 446 615 447 644 645 cell_1rw
* cell instance $28901 r0 *1 133.95,136.5
X$28901 446 614 447 644 645 cell_1rw
* cell instance $28902 m0 *1 133.95,139.23
X$28902 446 617 447 644 645 cell_1rw
* cell instance $28903 m0 *1 133.95,141.96
X$28903 446 618 447 644 645 cell_1rw
* cell instance $28904 r0 *1 133.95,139.23
X$28904 446 616 447 644 645 cell_1rw
* cell instance $28905 r0 *1 133.95,141.96
X$28905 446 619 447 644 645 cell_1rw
* cell instance $28906 m0 *1 133.95,144.69
X$28906 446 620 447 644 645 cell_1rw
* cell instance $28907 m0 *1 133.95,147.42
X$28907 446 622 447 644 645 cell_1rw
* cell instance $28908 r0 *1 133.95,144.69
X$28908 446 621 447 644 645 cell_1rw
* cell instance $28909 m0 *1 133.95,150.15
X$28909 446 624 447 644 645 cell_1rw
* cell instance $28910 r0 *1 133.95,147.42
X$28910 446 623 447 644 645 cell_1rw
* cell instance $28911 r0 *1 133.95,150.15
X$28911 446 625 447 644 645 cell_1rw
* cell instance $28912 m0 *1 133.95,152.88
X$28912 446 626 447 644 645 cell_1rw
* cell instance $28913 r0 *1 133.95,152.88
X$28913 446 627 447 644 645 cell_1rw
* cell instance $28914 m0 *1 133.95,155.61
X$28914 446 628 447 644 645 cell_1rw
* cell instance $28915 r0 *1 133.95,155.61
X$28915 446 629 447 644 645 cell_1rw
* cell instance $28916 m0 *1 133.95,158.34
X$28916 446 630 447 644 645 cell_1rw
* cell instance $28917 r0 *1 133.95,158.34
X$28917 446 631 447 644 645 cell_1rw
* cell instance $28918 m0 *1 133.95,161.07
X$28918 446 632 447 644 645 cell_1rw
* cell instance $28919 r0 *1 133.95,161.07
X$28919 446 633 447 644 645 cell_1rw
* cell instance $28920 m0 *1 133.95,163.8
X$28920 446 634 447 644 645 cell_1rw
* cell instance $28921 r0 *1 133.95,163.8
X$28921 446 635 447 644 645 cell_1rw
* cell instance $28922 m0 *1 133.95,166.53
X$28922 446 637 447 644 645 cell_1rw
* cell instance $28923 r0 *1 133.95,166.53
X$28923 446 636 447 644 645 cell_1rw
* cell instance $28924 m0 *1 133.95,169.26
X$28924 446 639 447 644 645 cell_1rw
* cell instance $28925 r0 *1 133.95,169.26
X$28925 446 638 447 644 645 cell_1rw
* cell instance $28926 m0 *1 133.95,171.99
X$28926 446 640 447 644 645 cell_1rw
* cell instance $28927 m0 *1 133.95,174.72
X$28927 446 642 447 644 645 cell_1rw
* cell instance $28928 r0 *1 133.95,171.99
X$28928 446 641 447 644 645 cell_1rw
* cell instance $28929 r0 *1 133.95,174.72
X$28929 446 643 447 644 645 cell_1rw
* cell instance $28930 m0 *1 134.655,90.09
X$28930 448 581 449 644 645 cell_1rw
* cell instance $28931 r0 *1 134.655,90.09
X$28931 448 580 449 644 645 cell_1rw
* cell instance $28932 m0 *1 134.655,92.82
X$28932 448 583 449 644 645 cell_1rw
* cell instance $28933 r0 *1 134.655,92.82
X$28933 448 582 449 644 645 cell_1rw
* cell instance $28934 m0 *1 134.655,95.55
X$28934 448 584 449 644 645 cell_1rw
* cell instance $28935 r0 *1 134.655,95.55
X$28935 448 585 449 644 645 cell_1rw
* cell instance $28936 m0 *1 134.655,98.28
X$28936 448 586 449 644 645 cell_1rw
* cell instance $28937 r0 *1 134.655,98.28
X$28937 448 587 449 644 645 cell_1rw
* cell instance $28938 m0 *1 134.655,101.01
X$28938 448 588 449 644 645 cell_1rw
* cell instance $28939 r0 *1 134.655,101.01
X$28939 448 589 449 644 645 cell_1rw
* cell instance $28940 m0 *1 134.655,103.74
X$28940 448 590 449 644 645 cell_1rw
* cell instance $28941 m0 *1 134.655,106.47
X$28941 448 593 449 644 645 cell_1rw
* cell instance $28942 r0 *1 134.655,103.74
X$28942 448 591 449 644 645 cell_1rw
* cell instance $28943 r0 *1 134.655,106.47
X$28943 448 592 449 644 645 cell_1rw
* cell instance $28944 m0 *1 134.655,109.2
X$28944 448 594 449 644 645 cell_1rw
* cell instance $28945 r0 *1 134.655,109.2
X$28945 448 595 449 644 645 cell_1rw
* cell instance $28946 m0 *1 134.655,111.93
X$28946 448 597 449 644 645 cell_1rw
* cell instance $28947 r0 *1 134.655,111.93
X$28947 448 596 449 644 645 cell_1rw
* cell instance $28948 m0 *1 134.655,114.66
X$28948 448 598 449 644 645 cell_1rw
* cell instance $28949 r0 *1 134.655,114.66
X$28949 448 599 449 644 645 cell_1rw
* cell instance $28950 m0 *1 134.655,117.39
X$28950 448 600 449 644 645 cell_1rw
* cell instance $28951 r0 *1 134.655,117.39
X$28951 448 601 449 644 645 cell_1rw
* cell instance $28952 m0 *1 134.655,120.12
X$28952 448 602 449 644 645 cell_1rw
* cell instance $28953 r0 *1 134.655,120.12
X$28953 448 603 449 644 645 cell_1rw
* cell instance $28954 m0 *1 134.655,122.85
X$28954 448 604 449 644 645 cell_1rw
* cell instance $28955 m0 *1 134.655,125.58
X$28955 448 606 449 644 645 cell_1rw
* cell instance $28956 r0 *1 134.655,122.85
X$28956 448 605 449 644 645 cell_1rw
* cell instance $28957 r0 *1 134.655,125.58
X$28957 448 607 449 644 645 cell_1rw
* cell instance $28958 m0 *1 134.655,128.31
X$28958 448 609 449 644 645 cell_1rw
* cell instance $28959 r0 *1 134.655,128.31
X$28959 448 608 449 644 645 cell_1rw
* cell instance $28960 m0 *1 134.655,131.04
X$28960 448 610 449 644 645 cell_1rw
* cell instance $28961 r0 *1 134.655,131.04
X$28961 448 611 449 644 645 cell_1rw
* cell instance $28962 m0 *1 134.655,133.77
X$28962 448 612 449 644 645 cell_1rw
* cell instance $28963 r0 *1 134.655,133.77
X$28963 448 613 449 644 645 cell_1rw
* cell instance $28964 m0 *1 134.655,136.5
X$28964 448 615 449 644 645 cell_1rw
* cell instance $28965 r0 *1 134.655,136.5
X$28965 448 614 449 644 645 cell_1rw
* cell instance $28966 m0 *1 134.655,139.23
X$28966 448 617 449 644 645 cell_1rw
* cell instance $28967 r0 *1 134.655,139.23
X$28967 448 616 449 644 645 cell_1rw
* cell instance $28968 m0 *1 134.655,141.96
X$28968 448 618 449 644 645 cell_1rw
* cell instance $28969 r0 *1 134.655,141.96
X$28969 448 619 449 644 645 cell_1rw
* cell instance $28970 m0 *1 134.655,144.69
X$28970 448 620 449 644 645 cell_1rw
* cell instance $28971 r0 *1 134.655,144.69
X$28971 448 621 449 644 645 cell_1rw
* cell instance $28972 m0 *1 134.655,147.42
X$28972 448 622 449 644 645 cell_1rw
* cell instance $28973 r0 *1 134.655,147.42
X$28973 448 623 449 644 645 cell_1rw
* cell instance $28974 m0 *1 134.655,150.15
X$28974 448 624 449 644 645 cell_1rw
* cell instance $28975 r0 *1 134.655,150.15
X$28975 448 625 449 644 645 cell_1rw
* cell instance $28976 m0 *1 134.655,152.88
X$28976 448 626 449 644 645 cell_1rw
* cell instance $28977 r0 *1 134.655,152.88
X$28977 448 627 449 644 645 cell_1rw
* cell instance $28978 m0 *1 134.655,155.61
X$28978 448 628 449 644 645 cell_1rw
* cell instance $28979 r0 *1 134.655,155.61
X$28979 448 629 449 644 645 cell_1rw
* cell instance $28980 m0 *1 134.655,158.34
X$28980 448 630 449 644 645 cell_1rw
* cell instance $28981 r0 *1 134.655,158.34
X$28981 448 631 449 644 645 cell_1rw
* cell instance $28982 m0 *1 134.655,161.07
X$28982 448 632 449 644 645 cell_1rw
* cell instance $28983 r0 *1 134.655,161.07
X$28983 448 633 449 644 645 cell_1rw
* cell instance $28984 m0 *1 134.655,163.8
X$28984 448 634 449 644 645 cell_1rw
* cell instance $28985 r0 *1 134.655,163.8
X$28985 448 635 449 644 645 cell_1rw
* cell instance $28986 m0 *1 134.655,166.53
X$28986 448 637 449 644 645 cell_1rw
* cell instance $28987 m0 *1 134.655,169.26
X$28987 448 639 449 644 645 cell_1rw
* cell instance $28988 r0 *1 134.655,166.53
X$28988 448 636 449 644 645 cell_1rw
* cell instance $28989 r0 *1 134.655,169.26
X$28989 448 638 449 644 645 cell_1rw
* cell instance $28990 m0 *1 134.655,171.99
X$28990 448 640 449 644 645 cell_1rw
* cell instance $28991 r0 *1 134.655,171.99
X$28991 448 641 449 644 645 cell_1rw
* cell instance $28992 m0 *1 134.655,174.72
X$28992 448 642 449 644 645 cell_1rw
* cell instance $28993 r0 *1 134.655,174.72
X$28993 448 643 449 644 645 cell_1rw
* cell instance $28994 m0 *1 135.36,90.09
X$28994 450 581 451 644 645 cell_1rw
* cell instance $28995 m0 *1 135.36,92.82
X$28995 450 583 451 644 645 cell_1rw
* cell instance $28996 r0 *1 135.36,90.09
X$28996 450 580 451 644 645 cell_1rw
* cell instance $28997 r0 *1 135.36,92.82
X$28997 450 582 451 644 645 cell_1rw
* cell instance $28998 m0 *1 135.36,95.55
X$28998 450 584 451 644 645 cell_1rw
* cell instance $28999 r0 *1 135.36,95.55
X$28999 450 585 451 644 645 cell_1rw
* cell instance $29000 m0 *1 135.36,98.28
X$29000 450 586 451 644 645 cell_1rw
* cell instance $29001 r0 *1 135.36,98.28
X$29001 450 587 451 644 645 cell_1rw
* cell instance $29002 m0 *1 135.36,101.01
X$29002 450 588 451 644 645 cell_1rw
* cell instance $29003 r0 *1 135.36,101.01
X$29003 450 589 451 644 645 cell_1rw
* cell instance $29004 m0 *1 135.36,103.74
X$29004 450 590 451 644 645 cell_1rw
* cell instance $29005 r0 *1 135.36,103.74
X$29005 450 591 451 644 645 cell_1rw
* cell instance $29006 m0 *1 135.36,106.47
X$29006 450 593 451 644 645 cell_1rw
* cell instance $29007 m0 *1 135.36,109.2
X$29007 450 594 451 644 645 cell_1rw
* cell instance $29008 r0 *1 135.36,106.47
X$29008 450 592 451 644 645 cell_1rw
* cell instance $29009 r0 *1 135.36,109.2
X$29009 450 595 451 644 645 cell_1rw
* cell instance $29010 m0 *1 135.36,111.93
X$29010 450 597 451 644 645 cell_1rw
* cell instance $29011 r0 *1 135.36,111.93
X$29011 450 596 451 644 645 cell_1rw
* cell instance $29012 m0 *1 135.36,114.66
X$29012 450 598 451 644 645 cell_1rw
* cell instance $29013 r0 *1 135.36,114.66
X$29013 450 599 451 644 645 cell_1rw
* cell instance $29014 m0 *1 135.36,117.39
X$29014 450 600 451 644 645 cell_1rw
* cell instance $29015 r0 *1 135.36,117.39
X$29015 450 601 451 644 645 cell_1rw
* cell instance $29016 m0 *1 135.36,120.12
X$29016 450 602 451 644 645 cell_1rw
* cell instance $29017 r0 *1 135.36,120.12
X$29017 450 603 451 644 645 cell_1rw
* cell instance $29018 m0 *1 135.36,122.85
X$29018 450 604 451 644 645 cell_1rw
* cell instance $29019 m0 *1 135.36,125.58
X$29019 450 606 451 644 645 cell_1rw
* cell instance $29020 r0 *1 135.36,122.85
X$29020 450 605 451 644 645 cell_1rw
* cell instance $29021 r0 *1 135.36,125.58
X$29021 450 607 451 644 645 cell_1rw
* cell instance $29022 m0 *1 135.36,128.31
X$29022 450 609 451 644 645 cell_1rw
* cell instance $29023 r0 *1 135.36,128.31
X$29023 450 608 451 644 645 cell_1rw
* cell instance $29024 m0 *1 135.36,131.04
X$29024 450 610 451 644 645 cell_1rw
* cell instance $29025 r0 *1 135.36,131.04
X$29025 450 611 451 644 645 cell_1rw
* cell instance $29026 m0 *1 135.36,133.77
X$29026 450 612 451 644 645 cell_1rw
* cell instance $29027 r0 *1 135.36,133.77
X$29027 450 613 451 644 645 cell_1rw
* cell instance $29028 m0 *1 135.36,136.5
X$29028 450 615 451 644 645 cell_1rw
* cell instance $29029 r0 *1 135.36,136.5
X$29029 450 614 451 644 645 cell_1rw
* cell instance $29030 m0 *1 135.36,139.23
X$29030 450 617 451 644 645 cell_1rw
* cell instance $29031 r0 *1 135.36,139.23
X$29031 450 616 451 644 645 cell_1rw
* cell instance $29032 m0 *1 135.36,141.96
X$29032 450 618 451 644 645 cell_1rw
* cell instance $29033 m0 *1 135.36,144.69
X$29033 450 620 451 644 645 cell_1rw
* cell instance $29034 r0 *1 135.36,141.96
X$29034 450 619 451 644 645 cell_1rw
* cell instance $29035 r0 *1 135.36,144.69
X$29035 450 621 451 644 645 cell_1rw
* cell instance $29036 m0 *1 135.36,147.42
X$29036 450 622 451 644 645 cell_1rw
* cell instance $29037 r0 *1 135.36,147.42
X$29037 450 623 451 644 645 cell_1rw
* cell instance $29038 m0 *1 135.36,150.15
X$29038 450 624 451 644 645 cell_1rw
* cell instance $29039 r0 *1 135.36,150.15
X$29039 450 625 451 644 645 cell_1rw
* cell instance $29040 m0 *1 135.36,152.88
X$29040 450 626 451 644 645 cell_1rw
* cell instance $29041 r0 *1 135.36,152.88
X$29041 450 627 451 644 645 cell_1rw
* cell instance $29042 m0 *1 135.36,155.61
X$29042 450 628 451 644 645 cell_1rw
* cell instance $29043 r0 *1 135.36,155.61
X$29043 450 629 451 644 645 cell_1rw
* cell instance $29044 m0 *1 135.36,158.34
X$29044 450 630 451 644 645 cell_1rw
* cell instance $29045 r0 *1 135.36,158.34
X$29045 450 631 451 644 645 cell_1rw
* cell instance $29046 m0 *1 135.36,161.07
X$29046 450 632 451 644 645 cell_1rw
* cell instance $29047 r0 *1 135.36,161.07
X$29047 450 633 451 644 645 cell_1rw
* cell instance $29048 m0 *1 135.36,163.8
X$29048 450 634 451 644 645 cell_1rw
* cell instance $29049 r0 *1 135.36,163.8
X$29049 450 635 451 644 645 cell_1rw
* cell instance $29050 m0 *1 135.36,166.53
X$29050 450 637 451 644 645 cell_1rw
* cell instance $29051 r0 *1 135.36,166.53
X$29051 450 636 451 644 645 cell_1rw
* cell instance $29052 m0 *1 135.36,169.26
X$29052 450 639 451 644 645 cell_1rw
* cell instance $29053 r0 *1 135.36,169.26
X$29053 450 638 451 644 645 cell_1rw
* cell instance $29054 m0 *1 135.36,171.99
X$29054 450 640 451 644 645 cell_1rw
* cell instance $29055 m0 *1 135.36,174.72
X$29055 450 642 451 644 645 cell_1rw
* cell instance $29056 r0 *1 135.36,171.99
X$29056 450 641 451 644 645 cell_1rw
* cell instance $29057 r0 *1 135.36,174.72
X$29057 450 643 451 644 645 cell_1rw
* cell instance $29058 m0 *1 136.065,90.09
X$29058 452 581 453 644 645 cell_1rw
* cell instance $29059 r0 *1 136.065,90.09
X$29059 452 580 453 644 645 cell_1rw
* cell instance $29060 m0 *1 136.065,92.82
X$29060 452 583 453 644 645 cell_1rw
* cell instance $29061 m0 *1 136.065,95.55
X$29061 452 584 453 644 645 cell_1rw
* cell instance $29062 r0 *1 136.065,92.82
X$29062 452 582 453 644 645 cell_1rw
* cell instance $29063 m0 *1 136.065,98.28
X$29063 452 586 453 644 645 cell_1rw
* cell instance $29064 r0 *1 136.065,95.55
X$29064 452 585 453 644 645 cell_1rw
* cell instance $29065 r0 *1 136.065,98.28
X$29065 452 587 453 644 645 cell_1rw
* cell instance $29066 m0 *1 136.065,101.01
X$29066 452 588 453 644 645 cell_1rw
* cell instance $29067 r0 *1 136.065,101.01
X$29067 452 589 453 644 645 cell_1rw
* cell instance $29068 m0 *1 136.065,103.74
X$29068 452 590 453 644 645 cell_1rw
* cell instance $29069 r0 *1 136.065,103.74
X$29069 452 591 453 644 645 cell_1rw
* cell instance $29070 m0 *1 136.065,106.47
X$29070 452 593 453 644 645 cell_1rw
* cell instance $29071 r0 *1 136.065,106.47
X$29071 452 592 453 644 645 cell_1rw
* cell instance $29072 m0 *1 136.065,109.2
X$29072 452 594 453 644 645 cell_1rw
* cell instance $29073 r0 *1 136.065,109.2
X$29073 452 595 453 644 645 cell_1rw
* cell instance $29074 m0 *1 136.065,111.93
X$29074 452 597 453 644 645 cell_1rw
* cell instance $29075 r0 *1 136.065,111.93
X$29075 452 596 453 644 645 cell_1rw
* cell instance $29076 m0 *1 136.065,114.66
X$29076 452 598 453 644 645 cell_1rw
* cell instance $29077 m0 *1 136.065,117.39
X$29077 452 600 453 644 645 cell_1rw
* cell instance $29078 r0 *1 136.065,114.66
X$29078 452 599 453 644 645 cell_1rw
* cell instance $29079 m0 *1 136.065,120.12
X$29079 452 602 453 644 645 cell_1rw
* cell instance $29080 r0 *1 136.065,117.39
X$29080 452 601 453 644 645 cell_1rw
* cell instance $29081 r0 *1 136.065,120.12
X$29081 452 603 453 644 645 cell_1rw
* cell instance $29082 m0 *1 136.065,122.85
X$29082 452 604 453 644 645 cell_1rw
* cell instance $29083 r0 *1 136.065,122.85
X$29083 452 605 453 644 645 cell_1rw
* cell instance $29084 m0 *1 136.065,125.58
X$29084 452 606 453 644 645 cell_1rw
* cell instance $29085 m0 *1 136.065,128.31
X$29085 452 609 453 644 645 cell_1rw
* cell instance $29086 r0 *1 136.065,125.58
X$29086 452 607 453 644 645 cell_1rw
* cell instance $29087 r0 *1 136.065,128.31
X$29087 452 608 453 644 645 cell_1rw
* cell instance $29088 m0 *1 136.065,131.04
X$29088 452 610 453 644 645 cell_1rw
* cell instance $29089 r0 *1 136.065,131.04
X$29089 452 611 453 644 645 cell_1rw
* cell instance $29090 m0 *1 136.065,133.77
X$29090 452 612 453 644 645 cell_1rw
* cell instance $29091 r0 *1 136.065,133.77
X$29091 452 613 453 644 645 cell_1rw
* cell instance $29092 m0 *1 136.065,136.5
X$29092 452 615 453 644 645 cell_1rw
* cell instance $29093 r0 *1 136.065,136.5
X$29093 452 614 453 644 645 cell_1rw
* cell instance $29094 m0 *1 136.065,139.23
X$29094 452 617 453 644 645 cell_1rw
* cell instance $29095 m0 *1 136.065,141.96
X$29095 452 618 453 644 645 cell_1rw
* cell instance $29096 r0 *1 136.065,139.23
X$29096 452 616 453 644 645 cell_1rw
* cell instance $29097 r0 *1 136.065,141.96
X$29097 452 619 453 644 645 cell_1rw
* cell instance $29098 m0 *1 136.065,144.69
X$29098 452 620 453 644 645 cell_1rw
* cell instance $29099 r0 *1 136.065,144.69
X$29099 452 621 453 644 645 cell_1rw
* cell instance $29100 m0 *1 136.065,147.42
X$29100 452 622 453 644 645 cell_1rw
* cell instance $29101 r0 *1 136.065,147.42
X$29101 452 623 453 644 645 cell_1rw
* cell instance $29102 m0 *1 136.065,150.15
X$29102 452 624 453 644 645 cell_1rw
* cell instance $29103 r0 *1 136.065,150.15
X$29103 452 625 453 644 645 cell_1rw
* cell instance $29104 m0 *1 136.065,152.88
X$29104 452 626 453 644 645 cell_1rw
* cell instance $29105 r0 *1 136.065,152.88
X$29105 452 627 453 644 645 cell_1rw
* cell instance $29106 m0 *1 136.065,155.61
X$29106 452 628 453 644 645 cell_1rw
* cell instance $29107 r0 *1 136.065,155.61
X$29107 452 629 453 644 645 cell_1rw
* cell instance $29108 m0 *1 136.065,158.34
X$29108 452 630 453 644 645 cell_1rw
* cell instance $29109 r0 *1 136.065,158.34
X$29109 452 631 453 644 645 cell_1rw
* cell instance $29110 m0 *1 136.065,161.07
X$29110 452 632 453 644 645 cell_1rw
* cell instance $29111 r0 *1 136.065,161.07
X$29111 452 633 453 644 645 cell_1rw
* cell instance $29112 m0 *1 136.065,163.8
X$29112 452 634 453 644 645 cell_1rw
* cell instance $29113 r0 *1 136.065,163.8
X$29113 452 635 453 644 645 cell_1rw
* cell instance $29114 m0 *1 136.065,166.53
X$29114 452 637 453 644 645 cell_1rw
* cell instance $29115 r0 *1 136.065,166.53
X$29115 452 636 453 644 645 cell_1rw
* cell instance $29116 m0 *1 136.065,169.26
X$29116 452 639 453 644 645 cell_1rw
* cell instance $29117 r0 *1 136.065,169.26
X$29117 452 638 453 644 645 cell_1rw
* cell instance $29118 m0 *1 136.065,171.99
X$29118 452 640 453 644 645 cell_1rw
* cell instance $29119 r0 *1 136.065,171.99
X$29119 452 641 453 644 645 cell_1rw
* cell instance $29120 m0 *1 136.065,174.72
X$29120 452 642 453 644 645 cell_1rw
* cell instance $29121 r0 *1 136.065,174.72
X$29121 452 643 453 644 645 cell_1rw
* cell instance $29122 m0 *1 136.77,90.09
X$29122 454 581 455 644 645 cell_1rw
* cell instance $29123 m0 *1 136.77,92.82
X$29123 454 583 455 644 645 cell_1rw
* cell instance $29124 r0 *1 136.77,90.09
X$29124 454 580 455 644 645 cell_1rw
* cell instance $29125 r0 *1 136.77,92.82
X$29125 454 582 455 644 645 cell_1rw
* cell instance $29126 m0 *1 136.77,95.55
X$29126 454 584 455 644 645 cell_1rw
* cell instance $29127 r0 *1 136.77,95.55
X$29127 454 585 455 644 645 cell_1rw
* cell instance $29128 m0 *1 136.77,98.28
X$29128 454 586 455 644 645 cell_1rw
* cell instance $29129 r0 *1 136.77,98.28
X$29129 454 587 455 644 645 cell_1rw
* cell instance $29130 m0 *1 136.77,101.01
X$29130 454 588 455 644 645 cell_1rw
* cell instance $29131 r0 *1 136.77,101.01
X$29131 454 589 455 644 645 cell_1rw
* cell instance $29132 m0 *1 136.77,103.74
X$29132 454 590 455 644 645 cell_1rw
* cell instance $29133 r0 *1 136.77,103.74
X$29133 454 591 455 644 645 cell_1rw
* cell instance $29134 m0 *1 136.77,106.47
X$29134 454 593 455 644 645 cell_1rw
* cell instance $29135 m0 *1 136.77,109.2
X$29135 454 594 455 644 645 cell_1rw
* cell instance $29136 r0 *1 136.77,106.47
X$29136 454 592 455 644 645 cell_1rw
* cell instance $29137 m0 *1 136.77,111.93
X$29137 454 597 455 644 645 cell_1rw
* cell instance $29138 r0 *1 136.77,109.2
X$29138 454 595 455 644 645 cell_1rw
* cell instance $29139 r0 *1 136.77,111.93
X$29139 454 596 455 644 645 cell_1rw
* cell instance $29140 m0 *1 136.77,114.66
X$29140 454 598 455 644 645 cell_1rw
* cell instance $29141 r0 *1 136.77,114.66
X$29141 454 599 455 644 645 cell_1rw
* cell instance $29142 m0 *1 136.77,117.39
X$29142 454 600 455 644 645 cell_1rw
* cell instance $29143 r0 *1 136.77,117.39
X$29143 454 601 455 644 645 cell_1rw
* cell instance $29144 m0 *1 136.77,120.12
X$29144 454 602 455 644 645 cell_1rw
* cell instance $29145 r0 *1 136.77,120.12
X$29145 454 603 455 644 645 cell_1rw
* cell instance $29146 m0 *1 136.77,122.85
X$29146 454 604 455 644 645 cell_1rw
* cell instance $29147 r0 *1 136.77,122.85
X$29147 454 605 455 644 645 cell_1rw
* cell instance $29148 m0 *1 136.77,125.58
X$29148 454 606 455 644 645 cell_1rw
* cell instance $29149 m0 *1 136.77,128.31
X$29149 454 609 455 644 645 cell_1rw
* cell instance $29150 r0 *1 136.77,125.58
X$29150 454 607 455 644 645 cell_1rw
* cell instance $29151 m0 *1 136.77,131.04
X$29151 454 610 455 644 645 cell_1rw
* cell instance $29152 r0 *1 136.77,128.31
X$29152 454 608 455 644 645 cell_1rw
* cell instance $29153 r0 *1 136.77,131.04
X$29153 454 611 455 644 645 cell_1rw
* cell instance $29154 m0 *1 136.77,133.77
X$29154 454 612 455 644 645 cell_1rw
* cell instance $29155 r0 *1 136.77,133.77
X$29155 454 613 455 644 645 cell_1rw
* cell instance $29156 m0 *1 136.77,136.5
X$29156 454 615 455 644 645 cell_1rw
* cell instance $29157 r0 *1 136.77,136.5
X$29157 454 614 455 644 645 cell_1rw
* cell instance $29158 m0 *1 136.77,139.23
X$29158 454 617 455 644 645 cell_1rw
* cell instance $29159 r0 *1 136.77,139.23
X$29159 454 616 455 644 645 cell_1rw
* cell instance $29160 m0 *1 136.77,141.96
X$29160 454 618 455 644 645 cell_1rw
* cell instance $29161 r0 *1 136.77,141.96
X$29161 454 619 455 644 645 cell_1rw
* cell instance $29162 m0 *1 136.77,144.69
X$29162 454 620 455 644 645 cell_1rw
* cell instance $29163 m0 *1 136.77,147.42
X$29163 454 622 455 644 645 cell_1rw
* cell instance $29164 r0 *1 136.77,144.69
X$29164 454 621 455 644 645 cell_1rw
* cell instance $29165 r0 *1 136.77,147.42
X$29165 454 623 455 644 645 cell_1rw
* cell instance $29166 m0 *1 136.77,150.15
X$29166 454 624 455 644 645 cell_1rw
* cell instance $29167 r0 *1 136.77,150.15
X$29167 454 625 455 644 645 cell_1rw
* cell instance $29168 m0 *1 136.77,152.88
X$29168 454 626 455 644 645 cell_1rw
* cell instance $29169 m0 *1 136.77,155.61
X$29169 454 628 455 644 645 cell_1rw
* cell instance $29170 r0 *1 136.77,152.88
X$29170 454 627 455 644 645 cell_1rw
* cell instance $29171 r0 *1 136.77,155.61
X$29171 454 629 455 644 645 cell_1rw
* cell instance $29172 m0 *1 136.77,158.34
X$29172 454 630 455 644 645 cell_1rw
* cell instance $29173 r0 *1 136.77,158.34
X$29173 454 631 455 644 645 cell_1rw
* cell instance $29174 m0 *1 136.77,161.07
X$29174 454 632 455 644 645 cell_1rw
* cell instance $29175 r0 *1 136.77,161.07
X$29175 454 633 455 644 645 cell_1rw
* cell instance $29176 m0 *1 136.77,163.8
X$29176 454 634 455 644 645 cell_1rw
* cell instance $29177 r0 *1 136.77,163.8
X$29177 454 635 455 644 645 cell_1rw
* cell instance $29178 m0 *1 136.77,166.53
X$29178 454 637 455 644 645 cell_1rw
* cell instance $29179 r0 *1 136.77,166.53
X$29179 454 636 455 644 645 cell_1rw
* cell instance $29180 m0 *1 136.77,169.26
X$29180 454 639 455 644 645 cell_1rw
* cell instance $29181 r0 *1 136.77,169.26
X$29181 454 638 455 644 645 cell_1rw
* cell instance $29182 m0 *1 136.77,171.99
X$29182 454 640 455 644 645 cell_1rw
* cell instance $29183 m0 *1 136.77,174.72
X$29183 454 642 455 644 645 cell_1rw
* cell instance $29184 r0 *1 136.77,171.99
X$29184 454 641 455 644 645 cell_1rw
* cell instance $29185 r0 *1 136.77,174.72
X$29185 454 643 455 644 645 cell_1rw
* cell instance $29186 m0 *1 137.475,90.09
X$29186 456 581 457 644 645 cell_1rw
* cell instance $29187 r0 *1 137.475,90.09
X$29187 456 580 457 644 645 cell_1rw
* cell instance $29188 m0 *1 137.475,92.82
X$29188 456 583 457 644 645 cell_1rw
* cell instance $29189 m0 *1 137.475,95.55
X$29189 456 584 457 644 645 cell_1rw
* cell instance $29190 r0 *1 137.475,92.82
X$29190 456 582 457 644 645 cell_1rw
* cell instance $29191 r0 *1 137.475,95.55
X$29191 456 585 457 644 645 cell_1rw
* cell instance $29192 m0 *1 137.475,98.28
X$29192 456 586 457 644 645 cell_1rw
* cell instance $29193 r0 *1 137.475,98.28
X$29193 456 587 457 644 645 cell_1rw
* cell instance $29194 m0 *1 137.475,101.01
X$29194 456 588 457 644 645 cell_1rw
* cell instance $29195 r0 *1 137.475,101.01
X$29195 456 589 457 644 645 cell_1rw
* cell instance $29196 m0 *1 137.475,103.74
X$29196 456 590 457 644 645 cell_1rw
* cell instance $29197 r0 *1 137.475,103.74
X$29197 456 591 457 644 645 cell_1rw
* cell instance $29198 m0 *1 137.475,106.47
X$29198 456 593 457 644 645 cell_1rw
* cell instance $29199 r0 *1 137.475,106.47
X$29199 456 592 457 644 645 cell_1rw
* cell instance $29200 m0 *1 137.475,109.2
X$29200 456 594 457 644 645 cell_1rw
* cell instance $29201 r0 *1 137.475,109.2
X$29201 456 595 457 644 645 cell_1rw
* cell instance $29202 m0 *1 137.475,111.93
X$29202 456 597 457 644 645 cell_1rw
* cell instance $29203 r0 *1 137.475,111.93
X$29203 456 596 457 644 645 cell_1rw
* cell instance $29204 m0 *1 137.475,114.66
X$29204 456 598 457 644 645 cell_1rw
* cell instance $29205 r0 *1 137.475,114.66
X$29205 456 599 457 644 645 cell_1rw
* cell instance $29206 m0 *1 137.475,117.39
X$29206 456 600 457 644 645 cell_1rw
* cell instance $29207 r0 *1 137.475,117.39
X$29207 456 601 457 644 645 cell_1rw
* cell instance $29208 m0 *1 137.475,120.12
X$29208 456 602 457 644 645 cell_1rw
* cell instance $29209 r0 *1 137.475,120.12
X$29209 456 603 457 644 645 cell_1rw
* cell instance $29210 m0 *1 137.475,122.85
X$29210 456 604 457 644 645 cell_1rw
* cell instance $29211 r0 *1 137.475,122.85
X$29211 456 605 457 644 645 cell_1rw
* cell instance $29212 m0 *1 137.475,125.58
X$29212 456 606 457 644 645 cell_1rw
* cell instance $29213 r0 *1 137.475,125.58
X$29213 456 607 457 644 645 cell_1rw
* cell instance $29214 m0 *1 137.475,128.31
X$29214 456 609 457 644 645 cell_1rw
* cell instance $29215 r0 *1 137.475,128.31
X$29215 456 608 457 644 645 cell_1rw
* cell instance $29216 m0 *1 137.475,131.04
X$29216 456 610 457 644 645 cell_1rw
* cell instance $29217 r0 *1 137.475,131.04
X$29217 456 611 457 644 645 cell_1rw
* cell instance $29218 m0 *1 137.475,133.77
X$29218 456 612 457 644 645 cell_1rw
* cell instance $29219 m0 *1 137.475,136.5
X$29219 456 615 457 644 645 cell_1rw
* cell instance $29220 r0 *1 137.475,133.77
X$29220 456 613 457 644 645 cell_1rw
* cell instance $29221 r0 *1 137.475,136.5
X$29221 456 614 457 644 645 cell_1rw
* cell instance $29222 m0 *1 137.475,139.23
X$29222 456 617 457 644 645 cell_1rw
* cell instance $29223 r0 *1 137.475,139.23
X$29223 456 616 457 644 645 cell_1rw
* cell instance $29224 m0 *1 137.475,141.96
X$29224 456 618 457 644 645 cell_1rw
* cell instance $29225 r0 *1 137.475,141.96
X$29225 456 619 457 644 645 cell_1rw
* cell instance $29226 m0 *1 137.475,144.69
X$29226 456 620 457 644 645 cell_1rw
* cell instance $29227 r0 *1 137.475,144.69
X$29227 456 621 457 644 645 cell_1rw
* cell instance $29228 m0 *1 137.475,147.42
X$29228 456 622 457 644 645 cell_1rw
* cell instance $29229 r0 *1 137.475,147.42
X$29229 456 623 457 644 645 cell_1rw
* cell instance $29230 m0 *1 137.475,150.15
X$29230 456 624 457 644 645 cell_1rw
* cell instance $29231 r0 *1 137.475,150.15
X$29231 456 625 457 644 645 cell_1rw
* cell instance $29232 m0 *1 137.475,152.88
X$29232 456 626 457 644 645 cell_1rw
* cell instance $29233 r0 *1 137.475,152.88
X$29233 456 627 457 644 645 cell_1rw
* cell instance $29234 m0 *1 137.475,155.61
X$29234 456 628 457 644 645 cell_1rw
* cell instance $29235 r0 *1 137.475,155.61
X$29235 456 629 457 644 645 cell_1rw
* cell instance $29236 m0 *1 137.475,158.34
X$29236 456 630 457 644 645 cell_1rw
* cell instance $29237 r0 *1 137.475,158.34
X$29237 456 631 457 644 645 cell_1rw
* cell instance $29238 m0 *1 137.475,161.07
X$29238 456 632 457 644 645 cell_1rw
* cell instance $29239 r0 *1 137.475,161.07
X$29239 456 633 457 644 645 cell_1rw
* cell instance $29240 m0 *1 137.475,163.8
X$29240 456 634 457 644 645 cell_1rw
* cell instance $29241 m0 *1 137.475,166.53
X$29241 456 637 457 644 645 cell_1rw
* cell instance $29242 r0 *1 137.475,163.8
X$29242 456 635 457 644 645 cell_1rw
* cell instance $29243 r0 *1 137.475,166.53
X$29243 456 636 457 644 645 cell_1rw
* cell instance $29244 m0 *1 137.475,169.26
X$29244 456 639 457 644 645 cell_1rw
* cell instance $29245 r0 *1 137.475,169.26
X$29245 456 638 457 644 645 cell_1rw
* cell instance $29246 m0 *1 137.475,171.99
X$29246 456 640 457 644 645 cell_1rw
* cell instance $29247 r0 *1 137.475,171.99
X$29247 456 641 457 644 645 cell_1rw
* cell instance $29248 m0 *1 137.475,174.72
X$29248 456 642 457 644 645 cell_1rw
* cell instance $29249 r0 *1 137.475,174.72
X$29249 456 643 457 644 645 cell_1rw
* cell instance $29250 m0 *1 138.18,90.09
X$29250 458 581 459 644 645 cell_1rw
* cell instance $29251 r0 *1 138.18,90.09
X$29251 458 580 459 644 645 cell_1rw
* cell instance $29252 m0 *1 138.18,92.82
X$29252 458 583 459 644 645 cell_1rw
* cell instance $29253 r0 *1 138.18,92.82
X$29253 458 582 459 644 645 cell_1rw
* cell instance $29254 m0 *1 138.18,95.55
X$29254 458 584 459 644 645 cell_1rw
* cell instance $29255 r0 *1 138.18,95.55
X$29255 458 585 459 644 645 cell_1rw
* cell instance $29256 m0 *1 138.18,98.28
X$29256 458 586 459 644 645 cell_1rw
* cell instance $29257 r0 *1 138.18,98.28
X$29257 458 587 459 644 645 cell_1rw
* cell instance $29258 m0 *1 138.18,101.01
X$29258 458 588 459 644 645 cell_1rw
* cell instance $29259 r0 *1 138.18,101.01
X$29259 458 589 459 644 645 cell_1rw
* cell instance $29260 m0 *1 138.18,103.74
X$29260 458 590 459 644 645 cell_1rw
* cell instance $29261 r0 *1 138.18,103.74
X$29261 458 591 459 644 645 cell_1rw
* cell instance $29262 m0 *1 138.18,106.47
X$29262 458 593 459 644 645 cell_1rw
* cell instance $29263 r0 *1 138.18,106.47
X$29263 458 592 459 644 645 cell_1rw
* cell instance $29264 m0 *1 138.18,109.2
X$29264 458 594 459 644 645 cell_1rw
* cell instance $29265 r0 *1 138.18,109.2
X$29265 458 595 459 644 645 cell_1rw
* cell instance $29266 m0 *1 138.18,111.93
X$29266 458 597 459 644 645 cell_1rw
* cell instance $29267 r0 *1 138.18,111.93
X$29267 458 596 459 644 645 cell_1rw
* cell instance $29268 m0 *1 138.18,114.66
X$29268 458 598 459 644 645 cell_1rw
* cell instance $29269 r0 *1 138.18,114.66
X$29269 458 599 459 644 645 cell_1rw
* cell instance $29270 m0 *1 138.18,117.39
X$29270 458 600 459 644 645 cell_1rw
* cell instance $29271 r0 *1 138.18,117.39
X$29271 458 601 459 644 645 cell_1rw
* cell instance $29272 m0 *1 138.18,120.12
X$29272 458 602 459 644 645 cell_1rw
* cell instance $29273 r0 *1 138.18,120.12
X$29273 458 603 459 644 645 cell_1rw
* cell instance $29274 m0 *1 138.18,122.85
X$29274 458 604 459 644 645 cell_1rw
* cell instance $29275 r0 *1 138.18,122.85
X$29275 458 605 459 644 645 cell_1rw
* cell instance $29276 m0 *1 138.18,125.58
X$29276 458 606 459 644 645 cell_1rw
* cell instance $29277 r0 *1 138.18,125.58
X$29277 458 607 459 644 645 cell_1rw
* cell instance $29278 m0 *1 138.18,128.31
X$29278 458 609 459 644 645 cell_1rw
* cell instance $29279 r0 *1 138.18,128.31
X$29279 458 608 459 644 645 cell_1rw
* cell instance $29280 m0 *1 138.18,131.04
X$29280 458 610 459 644 645 cell_1rw
* cell instance $29281 r0 *1 138.18,131.04
X$29281 458 611 459 644 645 cell_1rw
* cell instance $29282 m0 *1 138.18,133.77
X$29282 458 612 459 644 645 cell_1rw
* cell instance $29283 r0 *1 138.18,133.77
X$29283 458 613 459 644 645 cell_1rw
* cell instance $29284 m0 *1 138.18,136.5
X$29284 458 615 459 644 645 cell_1rw
* cell instance $29285 m0 *1 138.18,139.23
X$29285 458 617 459 644 645 cell_1rw
* cell instance $29286 r0 *1 138.18,136.5
X$29286 458 614 459 644 645 cell_1rw
* cell instance $29287 r0 *1 138.18,139.23
X$29287 458 616 459 644 645 cell_1rw
* cell instance $29288 m0 *1 138.18,141.96
X$29288 458 618 459 644 645 cell_1rw
* cell instance $29289 r0 *1 138.18,141.96
X$29289 458 619 459 644 645 cell_1rw
* cell instance $29290 m0 *1 138.18,144.69
X$29290 458 620 459 644 645 cell_1rw
* cell instance $29291 m0 *1 138.18,147.42
X$29291 458 622 459 644 645 cell_1rw
* cell instance $29292 r0 *1 138.18,144.69
X$29292 458 621 459 644 645 cell_1rw
* cell instance $29293 m0 *1 138.18,150.15
X$29293 458 624 459 644 645 cell_1rw
* cell instance $29294 r0 *1 138.18,147.42
X$29294 458 623 459 644 645 cell_1rw
* cell instance $29295 r0 *1 138.18,150.15
X$29295 458 625 459 644 645 cell_1rw
* cell instance $29296 m0 *1 138.18,152.88
X$29296 458 626 459 644 645 cell_1rw
* cell instance $29297 r0 *1 138.18,152.88
X$29297 458 627 459 644 645 cell_1rw
* cell instance $29298 m0 *1 138.18,155.61
X$29298 458 628 459 644 645 cell_1rw
* cell instance $29299 m0 *1 138.18,158.34
X$29299 458 630 459 644 645 cell_1rw
* cell instance $29300 r0 *1 138.18,155.61
X$29300 458 629 459 644 645 cell_1rw
* cell instance $29301 r0 *1 138.18,158.34
X$29301 458 631 459 644 645 cell_1rw
* cell instance $29302 m0 *1 138.18,161.07
X$29302 458 632 459 644 645 cell_1rw
* cell instance $29303 r0 *1 138.18,161.07
X$29303 458 633 459 644 645 cell_1rw
* cell instance $29304 m0 *1 138.18,163.8
X$29304 458 634 459 644 645 cell_1rw
* cell instance $29305 r0 *1 138.18,163.8
X$29305 458 635 459 644 645 cell_1rw
* cell instance $29306 m0 *1 138.18,166.53
X$29306 458 637 459 644 645 cell_1rw
* cell instance $29307 m0 *1 138.18,169.26
X$29307 458 639 459 644 645 cell_1rw
* cell instance $29308 r0 *1 138.18,166.53
X$29308 458 636 459 644 645 cell_1rw
* cell instance $29309 r0 *1 138.18,169.26
X$29309 458 638 459 644 645 cell_1rw
* cell instance $29310 m0 *1 138.18,171.99
X$29310 458 640 459 644 645 cell_1rw
* cell instance $29311 r0 *1 138.18,171.99
X$29311 458 641 459 644 645 cell_1rw
* cell instance $29312 m0 *1 138.18,174.72
X$29312 458 642 459 644 645 cell_1rw
* cell instance $29313 r0 *1 138.18,174.72
X$29313 458 643 459 644 645 cell_1rw
* cell instance $29314 m0 *1 138.885,90.09
X$29314 460 581 461 644 645 cell_1rw
* cell instance $29315 r0 *1 138.885,90.09
X$29315 460 580 461 644 645 cell_1rw
* cell instance $29316 m0 *1 138.885,92.82
X$29316 460 583 461 644 645 cell_1rw
* cell instance $29317 r0 *1 138.885,92.82
X$29317 460 582 461 644 645 cell_1rw
* cell instance $29318 m0 *1 138.885,95.55
X$29318 460 584 461 644 645 cell_1rw
* cell instance $29319 r0 *1 138.885,95.55
X$29319 460 585 461 644 645 cell_1rw
* cell instance $29320 m0 *1 138.885,98.28
X$29320 460 586 461 644 645 cell_1rw
* cell instance $29321 r0 *1 138.885,98.28
X$29321 460 587 461 644 645 cell_1rw
* cell instance $29322 m0 *1 138.885,101.01
X$29322 460 588 461 644 645 cell_1rw
* cell instance $29323 r0 *1 138.885,101.01
X$29323 460 589 461 644 645 cell_1rw
* cell instance $29324 m0 *1 138.885,103.74
X$29324 460 590 461 644 645 cell_1rw
* cell instance $29325 m0 *1 138.885,106.47
X$29325 460 593 461 644 645 cell_1rw
* cell instance $29326 r0 *1 138.885,103.74
X$29326 460 591 461 644 645 cell_1rw
* cell instance $29327 r0 *1 138.885,106.47
X$29327 460 592 461 644 645 cell_1rw
* cell instance $29328 m0 *1 138.885,109.2
X$29328 460 594 461 644 645 cell_1rw
* cell instance $29329 m0 *1 138.885,111.93
X$29329 460 597 461 644 645 cell_1rw
* cell instance $29330 r0 *1 138.885,109.2
X$29330 460 595 461 644 645 cell_1rw
* cell instance $29331 r0 *1 138.885,111.93
X$29331 460 596 461 644 645 cell_1rw
* cell instance $29332 m0 *1 138.885,114.66
X$29332 460 598 461 644 645 cell_1rw
* cell instance $29333 m0 *1 138.885,117.39
X$29333 460 600 461 644 645 cell_1rw
* cell instance $29334 r0 *1 138.885,114.66
X$29334 460 599 461 644 645 cell_1rw
* cell instance $29335 r0 *1 138.885,117.39
X$29335 460 601 461 644 645 cell_1rw
* cell instance $29336 m0 *1 138.885,120.12
X$29336 460 602 461 644 645 cell_1rw
* cell instance $29337 m0 *1 138.885,122.85
X$29337 460 604 461 644 645 cell_1rw
* cell instance $29338 r0 *1 138.885,120.12
X$29338 460 603 461 644 645 cell_1rw
* cell instance $29339 r0 *1 138.885,122.85
X$29339 460 605 461 644 645 cell_1rw
* cell instance $29340 m0 *1 138.885,125.58
X$29340 460 606 461 644 645 cell_1rw
* cell instance $29341 r0 *1 138.885,125.58
X$29341 460 607 461 644 645 cell_1rw
* cell instance $29342 m0 *1 138.885,128.31
X$29342 460 609 461 644 645 cell_1rw
* cell instance $29343 r0 *1 138.885,128.31
X$29343 460 608 461 644 645 cell_1rw
* cell instance $29344 m0 *1 138.885,131.04
X$29344 460 610 461 644 645 cell_1rw
* cell instance $29345 r0 *1 138.885,131.04
X$29345 460 611 461 644 645 cell_1rw
* cell instance $29346 m0 *1 138.885,133.77
X$29346 460 612 461 644 645 cell_1rw
* cell instance $29347 r0 *1 138.885,133.77
X$29347 460 613 461 644 645 cell_1rw
* cell instance $29348 m0 *1 138.885,136.5
X$29348 460 615 461 644 645 cell_1rw
* cell instance $29349 r0 *1 138.885,136.5
X$29349 460 614 461 644 645 cell_1rw
* cell instance $29350 m0 *1 138.885,139.23
X$29350 460 617 461 644 645 cell_1rw
* cell instance $29351 r0 *1 138.885,139.23
X$29351 460 616 461 644 645 cell_1rw
* cell instance $29352 m0 *1 138.885,141.96
X$29352 460 618 461 644 645 cell_1rw
* cell instance $29353 r0 *1 138.885,141.96
X$29353 460 619 461 644 645 cell_1rw
* cell instance $29354 m0 *1 138.885,144.69
X$29354 460 620 461 644 645 cell_1rw
* cell instance $29355 r0 *1 138.885,144.69
X$29355 460 621 461 644 645 cell_1rw
* cell instance $29356 m0 *1 138.885,147.42
X$29356 460 622 461 644 645 cell_1rw
* cell instance $29357 r0 *1 138.885,147.42
X$29357 460 623 461 644 645 cell_1rw
* cell instance $29358 m0 *1 138.885,150.15
X$29358 460 624 461 644 645 cell_1rw
* cell instance $29359 r0 *1 138.885,150.15
X$29359 460 625 461 644 645 cell_1rw
* cell instance $29360 m0 *1 138.885,152.88
X$29360 460 626 461 644 645 cell_1rw
* cell instance $29361 r0 *1 138.885,152.88
X$29361 460 627 461 644 645 cell_1rw
* cell instance $29362 m0 *1 138.885,155.61
X$29362 460 628 461 644 645 cell_1rw
* cell instance $29363 r0 *1 138.885,155.61
X$29363 460 629 461 644 645 cell_1rw
* cell instance $29364 m0 *1 138.885,158.34
X$29364 460 630 461 644 645 cell_1rw
* cell instance $29365 r0 *1 138.885,158.34
X$29365 460 631 461 644 645 cell_1rw
* cell instance $29366 m0 *1 138.885,161.07
X$29366 460 632 461 644 645 cell_1rw
* cell instance $29367 r0 *1 138.885,161.07
X$29367 460 633 461 644 645 cell_1rw
* cell instance $29368 m0 *1 138.885,163.8
X$29368 460 634 461 644 645 cell_1rw
* cell instance $29369 r0 *1 138.885,163.8
X$29369 460 635 461 644 645 cell_1rw
* cell instance $29370 m0 *1 138.885,166.53
X$29370 460 637 461 644 645 cell_1rw
* cell instance $29371 m0 *1 138.885,169.26
X$29371 460 639 461 644 645 cell_1rw
* cell instance $29372 r0 *1 138.885,166.53
X$29372 460 636 461 644 645 cell_1rw
* cell instance $29373 r0 *1 138.885,169.26
X$29373 460 638 461 644 645 cell_1rw
* cell instance $29374 m0 *1 138.885,171.99
X$29374 460 640 461 644 645 cell_1rw
* cell instance $29375 r0 *1 138.885,171.99
X$29375 460 641 461 644 645 cell_1rw
* cell instance $29376 m0 *1 138.885,174.72
X$29376 460 642 461 644 645 cell_1rw
* cell instance $29377 r0 *1 138.885,174.72
X$29377 460 643 461 644 645 cell_1rw
* cell instance $29378 m0 *1 139.59,90.09
X$29378 462 581 463 644 645 cell_1rw
* cell instance $29379 r0 *1 139.59,90.09
X$29379 462 580 463 644 645 cell_1rw
* cell instance $29380 m0 *1 139.59,92.82
X$29380 462 583 463 644 645 cell_1rw
* cell instance $29381 r0 *1 139.59,92.82
X$29381 462 582 463 644 645 cell_1rw
* cell instance $29382 m0 *1 139.59,95.55
X$29382 462 584 463 644 645 cell_1rw
* cell instance $29383 r0 *1 139.59,95.55
X$29383 462 585 463 644 645 cell_1rw
* cell instance $29384 m0 *1 139.59,98.28
X$29384 462 586 463 644 645 cell_1rw
* cell instance $29385 r0 *1 139.59,98.28
X$29385 462 587 463 644 645 cell_1rw
* cell instance $29386 m0 *1 139.59,101.01
X$29386 462 588 463 644 645 cell_1rw
* cell instance $29387 r0 *1 139.59,101.01
X$29387 462 589 463 644 645 cell_1rw
* cell instance $29388 m0 *1 139.59,103.74
X$29388 462 590 463 644 645 cell_1rw
* cell instance $29389 r0 *1 139.59,103.74
X$29389 462 591 463 644 645 cell_1rw
* cell instance $29390 m0 *1 139.59,106.47
X$29390 462 593 463 644 645 cell_1rw
* cell instance $29391 r0 *1 139.59,106.47
X$29391 462 592 463 644 645 cell_1rw
* cell instance $29392 m0 *1 139.59,109.2
X$29392 462 594 463 644 645 cell_1rw
* cell instance $29393 m0 *1 139.59,111.93
X$29393 462 597 463 644 645 cell_1rw
* cell instance $29394 r0 *1 139.59,109.2
X$29394 462 595 463 644 645 cell_1rw
* cell instance $29395 r0 *1 139.59,111.93
X$29395 462 596 463 644 645 cell_1rw
* cell instance $29396 m0 *1 139.59,114.66
X$29396 462 598 463 644 645 cell_1rw
* cell instance $29397 r0 *1 139.59,114.66
X$29397 462 599 463 644 645 cell_1rw
* cell instance $29398 m0 *1 139.59,117.39
X$29398 462 600 463 644 645 cell_1rw
* cell instance $29399 r0 *1 139.59,117.39
X$29399 462 601 463 644 645 cell_1rw
* cell instance $29400 m0 *1 139.59,120.12
X$29400 462 602 463 644 645 cell_1rw
* cell instance $29401 r0 *1 139.59,120.12
X$29401 462 603 463 644 645 cell_1rw
* cell instance $29402 m0 *1 139.59,122.85
X$29402 462 604 463 644 645 cell_1rw
* cell instance $29403 m0 *1 139.59,125.58
X$29403 462 606 463 644 645 cell_1rw
* cell instance $29404 r0 *1 139.59,122.85
X$29404 462 605 463 644 645 cell_1rw
* cell instance $29405 r0 *1 139.59,125.58
X$29405 462 607 463 644 645 cell_1rw
* cell instance $29406 m0 *1 139.59,128.31
X$29406 462 609 463 644 645 cell_1rw
* cell instance $29407 r0 *1 139.59,128.31
X$29407 462 608 463 644 645 cell_1rw
* cell instance $29408 m0 *1 139.59,131.04
X$29408 462 610 463 644 645 cell_1rw
* cell instance $29409 m0 *1 139.59,133.77
X$29409 462 612 463 644 645 cell_1rw
* cell instance $29410 r0 *1 139.59,131.04
X$29410 462 611 463 644 645 cell_1rw
* cell instance $29411 r0 *1 139.59,133.77
X$29411 462 613 463 644 645 cell_1rw
* cell instance $29412 m0 *1 139.59,136.5
X$29412 462 615 463 644 645 cell_1rw
* cell instance $29413 r0 *1 139.59,136.5
X$29413 462 614 463 644 645 cell_1rw
* cell instance $29414 m0 *1 139.59,139.23
X$29414 462 617 463 644 645 cell_1rw
* cell instance $29415 m0 *1 139.59,141.96
X$29415 462 618 463 644 645 cell_1rw
* cell instance $29416 r0 *1 139.59,139.23
X$29416 462 616 463 644 645 cell_1rw
* cell instance $29417 r0 *1 139.59,141.96
X$29417 462 619 463 644 645 cell_1rw
* cell instance $29418 m0 *1 139.59,144.69
X$29418 462 620 463 644 645 cell_1rw
* cell instance $29419 m0 *1 139.59,147.42
X$29419 462 622 463 644 645 cell_1rw
* cell instance $29420 r0 *1 139.59,144.69
X$29420 462 621 463 644 645 cell_1rw
* cell instance $29421 r0 *1 139.59,147.42
X$29421 462 623 463 644 645 cell_1rw
* cell instance $29422 m0 *1 139.59,150.15
X$29422 462 624 463 644 645 cell_1rw
* cell instance $29423 m0 *1 139.59,152.88
X$29423 462 626 463 644 645 cell_1rw
* cell instance $29424 r0 *1 139.59,150.15
X$29424 462 625 463 644 645 cell_1rw
* cell instance $29425 r0 *1 139.59,152.88
X$29425 462 627 463 644 645 cell_1rw
* cell instance $29426 m0 *1 139.59,155.61
X$29426 462 628 463 644 645 cell_1rw
* cell instance $29427 r0 *1 139.59,155.61
X$29427 462 629 463 644 645 cell_1rw
* cell instance $29428 m0 *1 139.59,158.34
X$29428 462 630 463 644 645 cell_1rw
* cell instance $29429 r0 *1 139.59,158.34
X$29429 462 631 463 644 645 cell_1rw
* cell instance $29430 m0 *1 139.59,161.07
X$29430 462 632 463 644 645 cell_1rw
* cell instance $29431 m0 *1 139.59,163.8
X$29431 462 634 463 644 645 cell_1rw
* cell instance $29432 r0 *1 139.59,161.07
X$29432 462 633 463 644 645 cell_1rw
* cell instance $29433 m0 *1 139.59,166.53
X$29433 462 637 463 644 645 cell_1rw
* cell instance $29434 r0 *1 139.59,163.8
X$29434 462 635 463 644 645 cell_1rw
* cell instance $29435 r0 *1 139.59,166.53
X$29435 462 636 463 644 645 cell_1rw
* cell instance $29436 m0 *1 139.59,169.26
X$29436 462 639 463 644 645 cell_1rw
* cell instance $29437 r0 *1 139.59,169.26
X$29437 462 638 463 644 645 cell_1rw
* cell instance $29438 m0 *1 139.59,171.99
X$29438 462 640 463 644 645 cell_1rw
* cell instance $29439 r0 *1 139.59,171.99
X$29439 462 641 463 644 645 cell_1rw
* cell instance $29440 m0 *1 139.59,174.72
X$29440 462 642 463 644 645 cell_1rw
* cell instance $29441 r0 *1 139.59,174.72
X$29441 462 643 463 644 645 cell_1rw
* cell instance $29442 m0 *1 140.295,90.09
X$29442 464 581 465 644 645 cell_1rw
* cell instance $29443 r0 *1 140.295,90.09
X$29443 464 580 465 644 645 cell_1rw
* cell instance $29444 m0 *1 140.295,92.82
X$29444 464 583 465 644 645 cell_1rw
* cell instance $29445 r0 *1 140.295,92.82
X$29445 464 582 465 644 645 cell_1rw
* cell instance $29446 m0 *1 140.295,95.55
X$29446 464 584 465 644 645 cell_1rw
* cell instance $29447 r0 *1 140.295,95.55
X$29447 464 585 465 644 645 cell_1rw
* cell instance $29448 m0 *1 140.295,98.28
X$29448 464 586 465 644 645 cell_1rw
* cell instance $29449 r0 *1 140.295,98.28
X$29449 464 587 465 644 645 cell_1rw
* cell instance $29450 m0 *1 140.295,101.01
X$29450 464 588 465 644 645 cell_1rw
* cell instance $29451 m0 *1 140.295,103.74
X$29451 464 590 465 644 645 cell_1rw
* cell instance $29452 r0 *1 140.295,101.01
X$29452 464 589 465 644 645 cell_1rw
* cell instance $29453 r0 *1 140.295,103.74
X$29453 464 591 465 644 645 cell_1rw
* cell instance $29454 m0 *1 140.295,106.47
X$29454 464 593 465 644 645 cell_1rw
* cell instance $29455 r0 *1 140.295,106.47
X$29455 464 592 465 644 645 cell_1rw
* cell instance $29456 m0 *1 140.295,109.2
X$29456 464 594 465 644 645 cell_1rw
* cell instance $29457 r0 *1 140.295,109.2
X$29457 464 595 465 644 645 cell_1rw
* cell instance $29458 m0 *1 140.295,111.93
X$29458 464 597 465 644 645 cell_1rw
* cell instance $29459 r0 *1 140.295,111.93
X$29459 464 596 465 644 645 cell_1rw
* cell instance $29460 m0 *1 140.295,114.66
X$29460 464 598 465 644 645 cell_1rw
* cell instance $29461 r0 *1 140.295,114.66
X$29461 464 599 465 644 645 cell_1rw
* cell instance $29462 m0 *1 140.295,117.39
X$29462 464 600 465 644 645 cell_1rw
* cell instance $29463 m0 *1 140.295,120.12
X$29463 464 602 465 644 645 cell_1rw
* cell instance $29464 r0 *1 140.295,117.39
X$29464 464 601 465 644 645 cell_1rw
* cell instance $29465 r0 *1 140.295,120.12
X$29465 464 603 465 644 645 cell_1rw
* cell instance $29466 m0 *1 140.295,122.85
X$29466 464 604 465 644 645 cell_1rw
* cell instance $29467 r0 *1 140.295,122.85
X$29467 464 605 465 644 645 cell_1rw
* cell instance $29468 m0 *1 140.295,125.58
X$29468 464 606 465 644 645 cell_1rw
* cell instance $29469 r0 *1 140.295,125.58
X$29469 464 607 465 644 645 cell_1rw
* cell instance $29470 m0 *1 140.295,128.31
X$29470 464 609 465 644 645 cell_1rw
* cell instance $29471 r0 *1 140.295,128.31
X$29471 464 608 465 644 645 cell_1rw
* cell instance $29472 m0 *1 140.295,131.04
X$29472 464 610 465 644 645 cell_1rw
* cell instance $29473 r0 *1 140.295,131.04
X$29473 464 611 465 644 645 cell_1rw
* cell instance $29474 m0 *1 140.295,133.77
X$29474 464 612 465 644 645 cell_1rw
* cell instance $29475 r0 *1 140.295,133.77
X$29475 464 613 465 644 645 cell_1rw
* cell instance $29476 m0 *1 140.295,136.5
X$29476 464 615 465 644 645 cell_1rw
* cell instance $29477 r0 *1 140.295,136.5
X$29477 464 614 465 644 645 cell_1rw
* cell instance $29478 m0 *1 140.295,139.23
X$29478 464 617 465 644 645 cell_1rw
* cell instance $29479 r0 *1 140.295,139.23
X$29479 464 616 465 644 645 cell_1rw
* cell instance $29480 m0 *1 140.295,141.96
X$29480 464 618 465 644 645 cell_1rw
* cell instance $29481 r0 *1 140.295,141.96
X$29481 464 619 465 644 645 cell_1rw
* cell instance $29482 m0 *1 140.295,144.69
X$29482 464 620 465 644 645 cell_1rw
* cell instance $29483 r0 *1 140.295,144.69
X$29483 464 621 465 644 645 cell_1rw
* cell instance $29484 m0 *1 140.295,147.42
X$29484 464 622 465 644 645 cell_1rw
* cell instance $29485 r0 *1 140.295,147.42
X$29485 464 623 465 644 645 cell_1rw
* cell instance $29486 m0 *1 140.295,150.15
X$29486 464 624 465 644 645 cell_1rw
* cell instance $29487 r0 *1 140.295,150.15
X$29487 464 625 465 644 645 cell_1rw
* cell instance $29488 m0 *1 140.295,152.88
X$29488 464 626 465 644 645 cell_1rw
* cell instance $29489 m0 *1 140.295,155.61
X$29489 464 628 465 644 645 cell_1rw
* cell instance $29490 r0 *1 140.295,152.88
X$29490 464 627 465 644 645 cell_1rw
* cell instance $29491 r0 *1 140.295,155.61
X$29491 464 629 465 644 645 cell_1rw
* cell instance $29492 m0 *1 140.295,158.34
X$29492 464 630 465 644 645 cell_1rw
* cell instance $29493 r0 *1 140.295,158.34
X$29493 464 631 465 644 645 cell_1rw
* cell instance $29494 m0 *1 140.295,161.07
X$29494 464 632 465 644 645 cell_1rw
* cell instance $29495 r0 *1 140.295,161.07
X$29495 464 633 465 644 645 cell_1rw
* cell instance $29496 m0 *1 140.295,163.8
X$29496 464 634 465 644 645 cell_1rw
* cell instance $29497 m0 *1 140.295,166.53
X$29497 464 637 465 644 645 cell_1rw
* cell instance $29498 r0 *1 140.295,163.8
X$29498 464 635 465 644 645 cell_1rw
* cell instance $29499 r0 *1 140.295,166.53
X$29499 464 636 465 644 645 cell_1rw
* cell instance $29500 m0 *1 140.295,169.26
X$29500 464 639 465 644 645 cell_1rw
* cell instance $29501 m0 *1 140.295,171.99
X$29501 464 640 465 644 645 cell_1rw
* cell instance $29502 r0 *1 140.295,169.26
X$29502 464 638 465 644 645 cell_1rw
* cell instance $29503 r0 *1 140.295,171.99
X$29503 464 641 465 644 645 cell_1rw
* cell instance $29504 m0 *1 140.295,174.72
X$29504 464 642 465 644 645 cell_1rw
* cell instance $29505 r0 *1 140.295,174.72
X$29505 464 643 465 644 645 cell_1rw
* cell instance $29506 m0 *1 141,90.09
X$29506 466 581 467 644 645 cell_1rw
* cell instance $29507 r0 *1 141,90.09
X$29507 466 580 467 644 645 cell_1rw
* cell instance $29508 m0 *1 141,92.82
X$29508 466 583 467 644 645 cell_1rw
* cell instance $29509 r0 *1 141,92.82
X$29509 466 582 467 644 645 cell_1rw
* cell instance $29510 m0 *1 141,95.55
X$29510 466 584 467 644 645 cell_1rw
* cell instance $29511 m0 *1 141,98.28
X$29511 466 586 467 644 645 cell_1rw
* cell instance $29512 r0 *1 141,95.55
X$29512 466 585 467 644 645 cell_1rw
* cell instance $29513 r0 *1 141,98.28
X$29513 466 587 467 644 645 cell_1rw
* cell instance $29514 m0 *1 141,101.01
X$29514 466 588 467 644 645 cell_1rw
* cell instance $29515 r0 *1 141,101.01
X$29515 466 589 467 644 645 cell_1rw
* cell instance $29516 m0 *1 141,103.74
X$29516 466 590 467 644 645 cell_1rw
* cell instance $29517 r0 *1 141,103.74
X$29517 466 591 467 644 645 cell_1rw
* cell instance $29518 m0 *1 141,106.47
X$29518 466 593 467 644 645 cell_1rw
* cell instance $29519 r0 *1 141,106.47
X$29519 466 592 467 644 645 cell_1rw
* cell instance $29520 m0 *1 141,109.2
X$29520 466 594 467 644 645 cell_1rw
* cell instance $29521 r0 *1 141,109.2
X$29521 466 595 467 644 645 cell_1rw
* cell instance $29522 m0 *1 141,111.93
X$29522 466 597 467 644 645 cell_1rw
* cell instance $29523 r0 *1 141,111.93
X$29523 466 596 467 644 645 cell_1rw
* cell instance $29524 m0 *1 141,114.66
X$29524 466 598 467 644 645 cell_1rw
* cell instance $29525 r0 *1 141,114.66
X$29525 466 599 467 644 645 cell_1rw
* cell instance $29526 m0 *1 141,117.39
X$29526 466 600 467 644 645 cell_1rw
* cell instance $29527 m0 *1 141,120.12
X$29527 466 602 467 644 645 cell_1rw
* cell instance $29528 r0 *1 141,117.39
X$29528 466 601 467 644 645 cell_1rw
* cell instance $29529 m0 *1 141,122.85
X$29529 466 604 467 644 645 cell_1rw
* cell instance $29530 r0 *1 141,120.12
X$29530 466 603 467 644 645 cell_1rw
* cell instance $29531 m0 *1 141,125.58
X$29531 466 606 467 644 645 cell_1rw
* cell instance $29532 r0 *1 141,122.85
X$29532 466 605 467 644 645 cell_1rw
* cell instance $29533 m0 *1 141,128.31
X$29533 466 609 467 644 645 cell_1rw
* cell instance $29534 r0 *1 141,125.58
X$29534 466 607 467 644 645 cell_1rw
* cell instance $29535 r0 *1 141,128.31
X$29535 466 608 467 644 645 cell_1rw
* cell instance $29536 m0 *1 141,131.04
X$29536 466 610 467 644 645 cell_1rw
* cell instance $29537 m0 *1 141,133.77
X$29537 466 612 467 644 645 cell_1rw
* cell instance $29538 r0 *1 141,131.04
X$29538 466 611 467 644 645 cell_1rw
* cell instance $29539 r0 *1 141,133.77
X$29539 466 613 467 644 645 cell_1rw
* cell instance $29540 m0 *1 141,136.5
X$29540 466 615 467 644 645 cell_1rw
* cell instance $29541 r0 *1 141,136.5
X$29541 466 614 467 644 645 cell_1rw
* cell instance $29542 m0 *1 141,139.23
X$29542 466 617 467 644 645 cell_1rw
* cell instance $29543 r0 *1 141,139.23
X$29543 466 616 467 644 645 cell_1rw
* cell instance $29544 m0 *1 141,141.96
X$29544 466 618 467 644 645 cell_1rw
* cell instance $29545 r0 *1 141,141.96
X$29545 466 619 467 644 645 cell_1rw
* cell instance $29546 m0 *1 141,144.69
X$29546 466 620 467 644 645 cell_1rw
* cell instance $29547 r0 *1 141,144.69
X$29547 466 621 467 644 645 cell_1rw
* cell instance $29548 m0 *1 141,147.42
X$29548 466 622 467 644 645 cell_1rw
* cell instance $29549 r0 *1 141,147.42
X$29549 466 623 467 644 645 cell_1rw
* cell instance $29550 m0 *1 141,150.15
X$29550 466 624 467 644 645 cell_1rw
* cell instance $29551 r0 *1 141,150.15
X$29551 466 625 467 644 645 cell_1rw
* cell instance $29552 m0 *1 141,152.88
X$29552 466 626 467 644 645 cell_1rw
* cell instance $29553 r0 *1 141,152.88
X$29553 466 627 467 644 645 cell_1rw
* cell instance $29554 m0 *1 141,155.61
X$29554 466 628 467 644 645 cell_1rw
* cell instance $29555 m0 *1 141,158.34
X$29555 466 630 467 644 645 cell_1rw
* cell instance $29556 r0 *1 141,155.61
X$29556 466 629 467 644 645 cell_1rw
* cell instance $29557 r0 *1 141,158.34
X$29557 466 631 467 644 645 cell_1rw
* cell instance $29558 m0 *1 141,161.07
X$29558 466 632 467 644 645 cell_1rw
* cell instance $29559 r0 *1 141,161.07
X$29559 466 633 467 644 645 cell_1rw
* cell instance $29560 m0 *1 141,163.8
X$29560 466 634 467 644 645 cell_1rw
* cell instance $29561 r0 *1 141,163.8
X$29561 466 635 467 644 645 cell_1rw
* cell instance $29562 m0 *1 141,166.53
X$29562 466 637 467 644 645 cell_1rw
* cell instance $29563 m0 *1 141,169.26
X$29563 466 639 467 644 645 cell_1rw
* cell instance $29564 r0 *1 141,166.53
X$29564 466 636 467 644 645 cell_1rw
* cell instance $29565 r0 *1 141,169.26
X$29565 466 638 467 644 645 cell_1rw
* cell instance $29566 m0 *1 141,171.99
X$29566 466 640 467 644 645 cell_1rw
* cell instance $29567 m0 *1 141,174.72
X$29567 466 642 467 644 645 cell_1rw
* cell instance $29568 r0 *1 141,171.99
X$29568 466 641 467 644 645 cell_1rw
* cell instance $29569 r0 *1 141,174.72
X$29569 466 643 467 644 645 cell_1rw
* cell instance $29570 m0 *1 141.705,90.09
X$29570 468 581 469 644 645 cell_1rw
* cell instance $29571 r0 *1 141.705,90.09
X$29571 468 580 469 644 645 cell_1rw
* cell instance $29572 m0 *1 141.705,92.82
X$29572 468 583 469 644 645 cell_1rw
* cell instance $29573 m0 *1 141.705,95.55
X$29573 468 584 469 644 645 cell_1rw
* cell instance $29574 r0 *1 141.705,92.82
X$29574 468 582 469 644 645 cell_1rw
* cell instance $29575 r0 *1 141.705,95.55
X$29575 468 585 469 644 645 cell_1rw
* cell instance $29576 m0 *1 141.705,98.28
X$29576 468 586 469 644 645 cell_1rw
* cell instance $29577 r0 *1 141.705,98.28
X$29577 468 587 469 644 645 cell_1rw
* cell instance $29578 m0 *1 141.705,101.01
X$29578 468 588 469 644 645 cell_1rw
* cell instance $29579 m0 *1 141.705,103.74
X$29579 468 590 469 644 645 cell_1rw
* cell instance $29580 r0 *1 141.705,101.01
X$29580 468 589 469 644 645 cell_1rw
* cell instance $29581 r0 *1 141.705,103.74
X$29581 468 591 469 644 645 cell_1rw
* cell instance $29582 m0 *1 141.705,106.47
X$29582 468 593 469 644 645 cell_1rw
* cell instance $29583 r0 *1 141.705,106.47
X$29583 468 592 469 644 645 cell_1rw
* cell instance $29584 m0 *1 141.705,109.2
X$29584 468 594 469 644 645 cell_1rw
* cell instance $29585 m0 *1 141.705,111.93
X$29585 468 597 469 644 645 cell_1rw
* cell instance $29586 r0 *1 141.705,109.2
X$29586 468 595 469 644 645 cell_1rw
* cell instance $29587 r0 *1 141.705,111.93
X$29587 468 596 469 644 645 cell_1rw
* cell instance $29588 m0 *1 141.705,114.66
X$29588 468 598 469 644 645 cell_1rw
* cell instance $29589 r0 *1 141.705,114.66
X$29589 468 599 469 644 645 cell_1rw
* cell instance $29590 m0 *1 141.705,117.39
X$29590 468 600 469 644 645 cell_1rw
* cell instance $29591 r0 *1 141.705,117.39
X$29591 468 601 469 644 645 cell_1rw
* cell instance $29592 m0 *1 141.705,120.12
X$29592 468 602 469 644 645 cell_1rw
* cell instance $29593 m0 *1 141.705,122.85
X$29593 468 604 469 644 645 cell_1rw
* cell instance $29594 r0 *1 141.705,120.12
X$29594 468 603 469 644 645 cell_1rw
* cell instance $29595 m0 *1 141.705,125.58
X$29595 468 606 469 644 645 cell_1rw
* cell instance $29596 r0 *1 141.705,122.85
X$29596 468 605 469 644 645 cell_1rw
* cell instance $29597 r0 *1 141.705,125.58
X$29597 468 607 469 644 645 cell_1rw
* cell instance $29598 m0 *1 141.705,128.31
X$29598 468 609 469 644 645 cell_1rw
* cell instance $29599 m0 *1 141.705,131.04
X$29599 468 610 469 644 645 cell_1rw
* cell instance $29600 r0 *1 141.705,128.31
X$29600 468 608 469 644 645 cell_1rw
* cell instance $29601 r0 *1 141.705,131.04
X$29601 468 611 469 644 645 cell_1rw
* cell instance $29602 m0 *1 141.705,133.77
X$29602 468 612 469 644 645 cell_1rw
* cell instance $29603 r0 *1 141.705,133.77
X$29603 468 613 469 644 645 cell_1rw
* cell instance $29604 m0 *1 141.705,136.5
X$29604 468 615 469 644 645 cell_1rw
* cell instance $29605 r0 *1 141.705,136.5
X$29605 468 614 469 644 645 cell_1rw
* cell instance $29606 m0 *1 141.705,139.23
X$29606 468 617 469 644 645 cell_1rw
* cell instance $29607 r0 *1 141.705,139.23
X$29607 468 616 469 644 645 cell_1rw
* cell instance $29608 m0 *1 141.705,141.96
X$29608 468 618 469 644 645 cell_1rw
* cell instance $29609 r0 *1 141.705,141.96
X$29609 468 619 469 644 645 cell_1rw
* cell instance $29610 m0 *1 141.705,144.69
X$29610 468 620 469 644 645 cell_1rw
* cell instance $29611 r0 *1 141.705,144.69
X$29611 468 621 469 644 645 cell_1rw
* cell instance $29612 m0 *1 141.705,147.42
X$29612 468 622 469 644 645 cell_1rw
* cell instance $29613 r0 *1 141.705,147.42
X$29613 468 623 469 644 645 cell_1rw
* cell instance $29614 m0 *1 141.705,150.15
X$29614 468 624 469 644 645 cell_1rw
* cell instance $29615 r0 *1 141.705,150.15
X$29615 468 625 469 644 645 cell_1rw
* cell instance $29616 m0 *1 141.705,152.88
X$29616 468 626 469 644 645 cell_1rw
* cell instance $29617 r0 *1 141.705,152.88
X$29617 468 627 469 644 645 cell_1rw
* cell instance $29618 m0 *1 141.705,155.61
X$29618 468 628 469 644 645 cell_1rw
* cell instance $29619 r0 *1 141.705,155.61
X$29619 468 629 469 644 645 cell_1rw
* cell instance $29620 m0 *1 141.705,158.34
X$29620 468 630 469 644 645 cell_1rw
* cell instance $29621 r0 *1 141.705,158.34
X$29621 468 631 469 644 645 cell_1rw
* cell instance $29622 m0 *1 141.705,161.07
X$29622 468 632 469 644 645 cell_1rw
* cell instance $29623 r0 *1 141.705,161.07
X$29623 468 633 469 644 645 cell_1rw
* cell instance $29624 m0 *1 141.705,163.8
X$29624 468 634 469 644 645 cell_1rw
* cell instance $29625 r0 *1 141.705,163.8
X$29625 468 635 469 644 645 cell_1rw
* cell instance $29626 m0 *1 141.705,166.53
X$29626 468 637 469 644 645 cell_1rw
* cell instance $29627 r0 *1 141.705,166.53
X$29627 468 636 469 644 645 cell_1rw
* cell instance $29628 m0 *1 141.705,169.26
X$29628 468 639 469 644 645 cell_1rw
* cell instance $29629 r0 *1 141.705,169.26
X$29629 468 638 469 644 645 cell_1rw
* cell instance $29630 m0 *1 141.705,171.99
X$29630 468 640 469 644 645 cell_1rw
* cell instance $29631 r0 *1 141.705,171.99
X$29631 468 641 469 644 645 cell_1rw
* cell instance $29632 m0 *1 141.705,174.72
X$29632 468 642 469 644 645 cell_1rw
* cell instance $29633 r0 *1 141.705,174.72
X$29633 468 643 469 644 645 cell_1rw
* cell instance $29634 m0 *1 142.41,90.09
X$29634 470 581 471 644 645 cell_1rw
* cell instance $29635 r0 *1 142.41,90.09
X$29635 470 580 471 644 645 cell_1rw
* cell instance $29636 m0 *1 142.41,92.82
X$29636 470 583 471 644 645 cell_1rw
* cell instance $29637 m0 *1 142.41,95.55
X$29637 470 584 471 644 645 cell_1rw
* cell instance $29638 r0 *1 142.41,92.82
X$29638 470 582 471 644 645 cell_1rw
* cell instance $29639 r0 *1 142.41,95.55
X$29639 470 585 471 644 645 cell_1rw
* cell instance $29640 m0 *1 142.41,98.28
X$29640 470 586 471 644 645 cell_1rw
* cell instance $29641 r0 *1 142.41,98.28
X$29641 470 587 471 644 645 cell_1rw
* cell instance $29642 m0 *1 142.41,101.01
X$29642 470 588 471 644 645 cell_1rw
* cell instance $29643 m0 *1 142.41,103.74
X$29643 470 590 471 644 645 cell_1rw
* cell instance $29644 r0 *1 142.41,101.01
X$29644 470 589 471 644 645 cell_1rw
* cell instance $29645 m0 *1 142.41,106.47
X$29645 470 593 471 644 645 cell_1rw
* cell instance $29646 r0 *1 142.41,103.74
X$29646 470 591 471 644 645 cell_1rw
* cell instance $29647 m0 *1 142.41,109.2
X$29647 470 594 471 644 645 cell_1rw
* cell instance $29648 r0 *1 142.41,106.47
X$29648 470 592 471 644 645 cell_1rw
* cell instance $29649 m0 *1 142.41,111.93
X$29649 470 597 471 644 645 cell_1rw
* cell instance $29650 r0 *1 142.41,109.2
X$29650 470 595 471 644 645 cell_1rw
* cell instance $29651 r0 *1 142.41,111.93
X$29651 470 596 471 644 645 cell_1rw
* cell instance $29652 m0 *1 142.41,114.66
X$29652 470 598 471 644 645 cell_1rw
* cell instance $29653 r0 *1 142.41,114.66
X$29653 470 599 471 644 645 cell_1rw
* cell instance $29654 m0 *1 142.41,117.39
X$29654 470 600 471 644 645 cell_1rw
* cell instance $29655 r0 *1 142.41,117.39
X$29655 470 601 471 644 645 cell_1rw
* cell instance $29656 m0 *1 142.41,120.12
X$29656 470 602 471 644 645 cell_1rw
* cell instance $29657 r0 *1 142.41,120.12
X$29657 470 603 471 644 645 cell_1rw
* cell instance $29658 m0 *1 142.41,122.85
X$29658 470 604 471 644 645 cell_1rw
* cell instance $29659 r0 *1 142.41,122.85
X$29659 470 605 471 644 645 cell_1rw
* cell instance $29660 m0 *1 142.41,125.58
X$29660 470 606 471 644 645 cell_1rw
* cell instance $29661 m0 *1 142.41,128.31
X$29661 470 609 471 644 645 cell_1rw
* cell instance $29662 r0 *1 142.41,125.58
X$29662 470 607 471 644 645 cell_1rw
* cell instance $29663 r0 *1 142.41,128.31
X$29663 470 608 471 644 645 cell_1rw
* cell instance $29664 m0 *1 142.41,131.04
X$29664 470 610 471 644 645 cell_1rw
* cell instance $29665 r0 *1 142.41,131.04
X$29665 470 611 471 644 645 cell_1rw
* cell instance $29666 m0 *1 142.41,133.77
X$29666 470 612 471 644 645 cell_1rw
* cell instance $29667 r0 *1 142.41,133.77
X$29667 470 613 471 644 645 cell_1rw
* cell instance $29668 m0 *1 142.41,136.5
X$29668 470 615 471 644 645 cell_1rw
* cell instance $29669 r0 *1 142.41,136.5
X$29669 470 614 471 644 645 cell_1rw
* cell instance $29670 m0 *1 142.41,139.23
X$29670 470 617 471 644 645 cell_1rw
* cell instance $29671 r0 *1 142.41,139.23
X$29671 470 616 471 644 645 cell_1rw
* cell instance $29672 m0 *1 142.41,141.96
X$29672 470 618 471 644 645 cell_1rw
* cell instance $29673 r0 *1 142.41,141.96
X$29673 470 619 471 644 645 cell_1rw
* cell instance $29674 m0 *1 142.41,144.69
X$29674 470 620 471 644 645 cell_1rw
* cell instance $29675 r0 *1 142.41,144.69
X$29675 470 621 471 644 645 cell_1rw
* cell instance $29676 m0 *1 142.41,147.42
X$29676 470 622 471 644 645 cell_1rw
* cell instance $29677 r0 *1 142.41,147.42
X$29677 470 623 471 644 645 cell_1rw
* cell instance $29678 m0 *1 142.41,150.15
X$29678 470 624 471 644 645 cell_1rw
* cell instance $29679 r0 *1 142.41,150.15
X$29679 470 625 471 644 645 cell_1rw
* cell instance $29680 m0 *1 142.41,152.88
X$29680 470 626 471 644 645 cell_1rw
* cell instance $29681 r0 *1 142.41,152.88
X$29681 470 627 471 644 645 cell_1rw
* cell instance $29682 m0 *1 142.41,155.61
X$29682 470 628 471 644 645 cell_1rw
* cell instance $29683 r0 *1 142.41,155.61
X$29683 470 629 471 644 645 cell_1rw
* cell instance $29684 m0 *1 142.41,158.34
X$29684 470 630 471 644 645 cell_1rw
* cell instance $29685 r0 *1 142.41,158.34
X$29685 470 631 471 644 645 cell_1rw
* cell instance $29686 m0 *1 142.41,161.07
X$29686 470 632 471 644 645 cell_1rw
* cell instance $29687 r0 *1 142.41,161.07
X$29687 470 633 471 644 645 cell_1rw
* cell instance $29688 m0 *1 142.41,163.8
X$29688 470 634 471 644 645 cell_1rw
* cell instance $29689 r0 *1 142.41,163.8
X$29689 470 635 471 644 645 cell_1rw
* cell instance $29690 m0 *1 142.41,166.53
X$29690 470 637 471 644 645 cell_1rw
* cell instance $29691 r0 *1 142.41,166.53
X$29691 470 636 471 644 645 cell_1rw
* cell instance $29692 m0 *1 142.41,169.26
X$29692 470 639 471 644 645 cell_1rw
* cell instance $29693 r0 *1 142.41,169.26
X$29693 470 638 471 644 645 cell_1rw
* cell instance $29694 m0 *1 142.41,171.99
X$29694 470 640 471 644 645 cell_1rw
* cell instance $29695 m0 *1 142.41,174.72
X$29695 470 642 471 644 645 cell_1rw
* cell instance $29696 r0 *1 142.41,171.99
X$29696 470 641 471 644 645 cell_1rw
* cell instance $29697 r0 *1 142.41,174.72
X$29697 470 643 471 644 645 cell_1rw
* cell instance $29698 m0 *1 143.115,90.09
X$29698 472 581 473 644 645 cell_1rw
* cell instance $29699 r0 *1 143.115,90.09
X$29699 472 580 473 644 645 cell_1rw
* cell instance $29700 m0 *1 143.115,92.82
X$29700 472 583 473 644 645 cell_1rw
* cell instance $29701 r0 *1 143.115,92.82
X$29701 472 582 473 644 645 cell_1rw
* cell instance $29702 m0 *1 143.115,95.55
X$29702 472 584 473 644 645 cell_1rw
* cell instance $29703 r0 *1 143.115,95.55
X$29703 472 585 473 644 645 cell_1rw
* cell instance $29704 m0 *1 143.115,98.28
X$29704 472 586 473 644 645 cell_1rw
* cell instance $29705 r0 *1 143.115,98.28
X$29705 472 587 473 644 645 cell_1rw
* cell instance $29706 m0 *1 143.115,101.01
X$29706 472 588 473 644 645 cell_1rw
* cell instance $29707 r0 *1 143.115,101.01
X$29707 472 589 473 644 645 cell_1rw
* cell instance $29708 m0 *1 143.115,103.74
X$29708 472 590 473 644 645 cell_1rw
* cell instance $29709 r0 *1 143.115,103.74
X$29709 472 591 473 644 645 cell_1rw
* cell instance $29710 m0 *1 143.115,106.47
X$29710 472 593 473 644 645 cell_1rw
* cell instance $29711 r0 *1 143.115,106.47
X$29711 472 592 473 644 645 cell_1rw
* cell instance $29712 m0 *1 143.115,109.2
X$29712 472 594 473 644 645 cell_1rw
* cell instance $29713 r0 *1 143.115,109.2
X$29713 472 595 473 644 645 cell_1rw
* cell instance $29714 m0 *1 143.115,111.93
X$29714 472 597 473 644 645 cell_1rw
* cell instance $29715 r0 *1 143.115,111.93
X$29715 472 596 473 644 645 cell_1rw
* cell instance $29716 m0 *1 143.115,114.66
X$29716 472 598 473 644 645 cell_1rw
* cell instance $29717 r0 *1 143.115,114.66
X$29717 472 599 473 644 645 cell_1rw
* cell instance $29718 m0 *1 143.115,117.39
X$29718 472 600 473 644 645 cell_1rw
* cell instance $29719 r0 *1 143.115,117.39
X$29719 472 601 473 644 645 cell_1rw
* cell instance $29720 m0 *1 143.115,120.12
X$29720 472 602 473 644 645 cell_1rw
* cell instance $29721 m0 *1 143.115,122.85
X$29721 472 604 473 644 645 cell_1rw
* cell instance $29722 r0 *1 143.115,120.12
X$29722 472 603 473 644 645 cell_1rw
* cell instance $29723 r0 *1 143.115,122.85
X$29723 472 605 473 644 645 cell_1rw
* cell instance $29724 m0 *1 143.115,125.58
X$29724 472 606 473 644 645 cell_1rw
* cell instance $29725 r0 *1 143.115,125.58
X$29725 472 607 473 644 645 cell_1rw
* cell instance $29726 m0 *1 143.115,128.31
X$29726 472 609 473 644 645 cell_1rw
* cell instance $29727 r0 *1 143.115,128.31
X$29727 472 608 473 644 645 cell_1rw
* cell instance $29728 m0 *1 143.115,131.04
X$29728 472 610 473 644 645 cell_1rw
* cell instance $29729 m0 *1 143.115,133.77
X$29729 472 612 473 644 645 cell_1rw
* cell instance $29730 r0 *1 143.115,131.04
X$29730 472 611 473 644 645 cell_1rw
* cell instance $29731 r0 *1 143.115,133.77
X$29731 472 613 473 644 645 cell_1rw
* cell instance $29732 m0 *1 143.115,136.5
X$29732 472 615 473 644 645 cell_1rw
* cell instance $29733 m0 *1 143.115,139.23
X$29733 472 617 473 644 645 cell_1rw
* cell instance $29734 r0 *1 143.115,136.5
X$29734 472 614 473 644 645 cell_1rw
* cell instance $29735 r0 *1 143.115,139.23
X$29735 472 616 473 644 645 cell_1rw
* cell instance $29736 m0 *1 143.115,141.96
X$29736 472 618 473 644 645 cell_1rw
* cell instance $29737 r0 *1 143.115,141.96
X$29737 472 619 473 644 645 cell_1rw
* cell instance $29738 m0 *1 143.115,144.69
X$29738 472 620 473 644 645 cell_1rw
* cell instance $29739 r0 *1 143.115,144.69
X$29739 472 621 473 644 645 cell_1rw
* cell instance $29740 m0 *1 143.115,147.42
X$29740 472 622 473 644 645 cell_1rw
* cell instance $29741 r0 *1 143.115,147.42
X$29741 472 623 473 644 645 cell_1rw
* cell instance $29742 m0 *1 143.115,150.15
X$29742 472 624 473 644 645 cell_1rw
* cell instance $29743 r0 *1 143.115,150.15
X$29743 472 625 473 644 645 cell_1rw
* cell instance $29744 m0 *1 143.115,152.88
X$29744 472 626 473 644 645 cell_1rw
* cell instance $29745 r0 *1 143.115,152.88
X$29745 472 627 473 644 645 cell_1rw
* cell instance $29746 m0 *1 143.115,155.61
X$29746 472 628 473 644 645 cell_1rw
* cell instance $29747 r0 *1 143.115,155.61
X$29747 472 629 473 644 645 cell_1rw
* cell instance $29748 m0 *1 143.115,158.34
X$29748 472 630 473 644 645 cell_1rw
* cell instance $29749 r0 *1 143.115,158.34
X$29749 472 631 473 644 645 cell_1rw
* cell instance $29750 m0 *1 143.115,161.07
X$29750 472 632 473 644 645 cell_1rw
* cell instance $29751 r0 *1 143.115,161.07
X$29751 472 633 473 644 645 cell_1rw
* cell instance $29752 m0 *1 143.115,163.8
X$29752 472 634 473 644 645 cell_1rw
* cell instance $29753 m0 *1 143.115,166.53
X$29753 472 637 473 644 645 cell_1rw
* cell instance $29754 r0 *1 143.115,163.8
X$29754 472 635 473 644 645 cell_1rw
* cell instance $29755 r0 *1 143.115,166.53
X$29755 472 636 473 644 645 cell_1rw
* cell instance $29756 m0 *1 143.115,169.26
X$29756 472 639 473 644 645 cell_1rw
* cell instance $29757 r0 *1 143.115,169.26
X$29757 472 638 473 644 645 cell_1rw
* cell instance $29758 m0 *1 143.115,171.99
X$29758 472 640 473 644 645 cell_1rw
* cell instance $29759 r0 *1 143.115,171.99
X$29759 472 641 473 644 645 cell_1rw
* cell instance $29760 m0 *1 143.115,174.72
X$29760 472 642 473 644 645 cell_1rw
* cell instance $29761 r0 *1 143.115,174.72
X$29761 472 643 473 644 645 cell_1rw
* cell instance $29762 m0 *1 143.82,90.09
X$29762 474 581 475 644 645 cell_1rw
* cell instance $29763 r0 *1 143.82,90.09
X$29763 474 580 475 644 645 cell_1rw
* cell instance $29764 m0 *1 143.82,92.82
X$29764 474 583 475 644 645 cell_1rw
* cell instance $29765 r0 *1 143.82,92.82
X$29765 474 582 475 644 645 cell_1rw
* cell instance $29766 m0 *1 143.82,95.55
X$29766 474 584 475 644 645 cell_1rw
* cell instance $29767 r0 *1 143.82,95.55
X$29767 474 585 475 644 645 cell_1rw
* cell instance $29768 m0 *1 143.82,98.28
X$29768 474 586 475 644 645 cell_1rw
* cell instance $29769 r0 *1 143.82,98.28
X$29769 474 587 475 644 645 cell_1rw
* cell instance $29770 m0 *1 143.82,101.01
X$29770 474 588 475 644 645 cell_1rw
* cell instance $29771 r0 *1 143.82,101.01
X$29771 474 589 475 644 645 cell_1rw
* cell instance $29772 m0 *1 143.82,103.74
X$29772 474 590 475 644 645 cell_1rw
* cell instance $29773 r0 *1 143.82,103.74
X$29773 474 591 475 644 645 cell_1rw
* cell instance $29774 m0 *1 143.82,106.47
X$29774 474 593 475 644 645 cell_1rw
* cell instance $29775 r0 *1 143.82,106.47
X$29775 474 592 475 644 645 cell_1rw
* cell instance $29776 m0 *1 143.82,109.2
X$29776 474 594 475 644 645 cell_1rw
* cell instance $29777 r0 *1 143.82,109.2
X$29777 474 595 475 644 645 cell_1rw
* cell instance $29778 m0 *1 143.82,111.93
X$29778 474 597 475 644 645 cell_1rw
* cell instance $29779 r0 *1 143.82,111.93
X$29779 474 596 475 644 645 cell_1rw
* cell instance $29780 m0 *1 143.82,114.66
X$29780 474 598 475 644 645 cell_1rw
* cell instance $29781 m0 *1 143.82,117.39
X$29781 474 600 475 644 645 cell_1rw
* cell instance $29782 r0 *1 143.82,114.66
X$29782 474 599 475 644 645 cell_1rw
* cell instance $29783 r0 *1 143.82,117.39
X$29783 474 601 475 644 645 cell_1rw
* cell instance $29784 m0 *1 143.82,120.12
X$29784 474 602 475 644 645 cell_1rw
* cell instance $29785 r0 *1 143.82,120.12
X$29785 474 603 475 644 645 cell_1rw
* cell instance $29786 m0 *1 143.82,122.85
X$29786 474 604 475 644 645 cell_1rw
* cell instance $29787 r0 *1 143.82,122.85
X$29787 474 605 475 644 645 cell_1rw
* cell instance $29788 m0 *1 143.82,125.58
X$29788 474 606 475 644 645 cell_1rw
* cell instance $29789 r0 *1 143.82,125.58
X$29789 474 607 475 644 645 cell_1rw
* cell instance $29790 m0 *1 143.82,128.31
X$29790 474 609 475 644 645 cell_1rw
* cell instance $29791 r0 *1 143.82,128.31
X$29791 474 608 475 644 645 cell_1rw
* cell instance $29792 m0 *1 143.82,131.04
X$29792 474 610 475 644 645 cell_1rw
* cell instance $29793 r0 *1 143.82,131.04
X$29793 474 611 475 644 645 cell_1rw
* cell instance $29794 m0 *1 143.82,133.77
X$29794 474 612 475 644 645 cell_1rw
* cell instance $29795 r0 *1 143.82,133.77
X$29795 474 613 475 644 645 cell_1rw
* cell instance $29796 m0 *1 143.82,136.5
X$29796 474 615 475 644 645 cell_1rw
* cell instance $29797 m0 *1 143.82,139.23
X$29797 474 617 475 644 645 cell_1rw
* cell instance $29798 r0 *1 143.82,136.5
X$29798 474 614 475 644 645 cell_1rw
* cell instance $29799 r0 *1 143.82,139.23
X$29799 474 616 475 644 645 cell_1rw
* cell instance $29800 m0 *1 143.82,141.96
X$29800 474 618 475 644 645 cell_1rw
* cell instance $29801 m0 *1 143.82,144.69
X$29801 474 620 475 644 645 cell_1rw
* cell instance $29802 r0 *1 143.82,141.96
X$29802 474 619 475 644 645 cell_1rw
* cell instance $29803 m0 *1 143.82,147.42
X$29803 474 622 475 644 645 cell_1rw
* cell instance $29804 r0 *1 143.82,144.69
X$29804 474 621 475 644 645 cell_1rw
* cell instance $29805 r0 *1 143.82,147.42
X$29805 474 623 475 644 645 cell_1rw
* cell instance $29806 m0 *1 143.82,150.15
X$29806 474 624 475 644 645 cell_1rw
* cell instance $29807 r0 *1 143.82,150.15
X$29807 474 625 475 644 645 cell_1rw
* cell instance $29808 m0 *1 143.82,152.88
X$29808 474 626 475 644 645 cell_1rw
* cell instance $29809 r0 *1 143.82,152.88
X$29809 474 627 475 644 645 cell_1rw
* cell instance $29810 m0 *1 143.82,155.61
X$29810 474 628 475 644 645 cell_1rw
* cell instance $29811 m0 *1 143.82,158.34
X$29811 474 630 475 644 645 cell_1rw
* cell instance $29812 r0 *1 143.82,155.61
X$29812 474 629 475 644 645 cell_1rw
* cell instance $29813 r0 *1 143.82,158.34
X$29813 474 631 475 644 645 cell_1rw
* cell instance $29814 m0 *1 143.82,161.07
X$29814 474 632 475 644 645 cell_1rw
* cell instance $29815 r0 *1 143.82,161.07
X$29815 474 633 475 644 645 cell_1rw
* cell instance $29816 m0 *1 143.82,163.8
X$29816 474 634 475 644 645 cell_1rw
* cell instance $29817 m0 *1 143.82,166.53
X$29817 474 637 475 644 645 cell_1rw
* cell instance $29818 r0 *1 143.82,163.8
X$29818 474 635 475 644 645 cell_1rw
* cell instance $29819 r0 *1 143.82,166.53
X$29819 474 636 475 644 645 cell_1rw
* cell instance $29820 m0 *1 143.82,169.26
X$29820 474 639 475 644 645 cell_1rw
* cell instance $29821 r0 *1 143.82,169.26
X$29821 474 638 475 644 645 cell_1rw
* cell instance $29822 m0 *1 143.82,171.99
X$29822 474 640 475 644 645 cell_1rw
* cell instance $29823 r0 *1 143.82,171.99
X$29823 474 641 475 644 645 cell_1rw
* cell instance $29824 m0 *1 143.82,174.72
X$29824 474 642 475 644 645 cell_1rw
* cell instance $29825 r0 *1 143.82,174.72
X$29825 474 643 475 644 645 cell_1rw
* cell instance $29826 m0 *1 144.525,90.09
X$29826 476 581 477 644 645 cell_1rw
* cell instance $29827 m0 *1 144.525,92.82
X$29827 476 583 477 644 645 cell_1rw
* cell instance $29828 r0 *1 144.525,90.09
X$29828 476 580 477 644 645 cell_1rw
* cell instance $29829 r0 *1 144.525,92.82
X$29829 476 582 477 644 645 cell_1rw
* cell instance $29830 m0 *1 144.525,95.55
X$29830 476 584 477 644 645 cell_1rw
* cell instance $29831 r0 *1 144.525,95.55
X$29831 476 585 477 644 645 cell_1rw
* cell instance $29832 m0 *1 144.525,98.28
X$29832 476 586 477 644 645 cell_1rw
* cell instance $29833 r0 *1 144.525,98.28
X$29833 476 587 477 644 645 cell_1rw
* cell instance $29834 m0 *1 144.525,101.01
X$29834 476 588 477 644 645 cell_1rw
* cell instance $29835 r0 *1 144.525,101.01
X$29835 476 589 477 644 645 cell_1rw
* cell instance $29836 m0 *1 144.525,103.74
X$29836 476 590 477 644 645 cell_1rw
* cell instance $29837 r0 *1 144.525,103.74
X$29837 476 591 477 644 645 cell_1rw
* cell instance $29838 m0 *1 144.525,106.47
X$29838 476 593 477 644 645 cell_1rw
* cell instance $29839 r0 *1 144.525,106.47
X$29839 476 592 477 644 645 cell_1rw
* cell instance $29840 m0 *1 144.525,109.2
X$29840 476 594 477 644 645 cell_1rw
* cell instance $29841 m0 *1 144.525,111.93
X$29841 476 597 477 644 645 cell_1rw
* cell instance $29842 r0 *1 144.525,109.2
X$29842 476 595 477 644 645 cell_1rw
* cell instance $29843 r0 *1 144.525,111.93
X$29843 476 596 477 644 645 cell_1rw
* cell instance $29844 m0 *1 144.525,114.66
X$29844 476 598 477 644 645 cell_1rw
* cell instance $29845 m0 *1 144.525,117.39
X$29845 476 600 477 644 645 cell_1rw
* cell instance $29846 r0 *1 144.525,114.66
X$29846 476 599 477 644 645 cell_1rw
* cell instance $29847 r0 *1 144.525,117.39
X$29847 476 601 477 644 645 cell_1rw
* cell instance $29848 m0 *1 144.525,120.12
X$29848 476 602 477 644 645 cell_1rw
* cell instance $29849 r0 *1 144.525,120.12
X$29849 476 603 477 644 645 cell_1rw
* cell instance $29850 m0 *1 144.525,122.85
X$29850 476 604 477 644 645 cell_1rw
* cell instance $29851 r0 *1 144.525,122.85
X$29851 476 605 477 644 645 cell_1rw
* cell instance $29852 m0 *1 144.525,125.58
X$29852 476 606 477 644 645 cell_1rw
* cell instance $29853 r0 *1 144.525,125.58
X$29853 476 607 477 644 645 cell_1rw
* cell instance $29854 m0 *1 144.525,128.31
X$29854 476 609 477 644 645 cell_1rw
* cell instance $29855 r0 *1 144.525,128.31
X$29855 476 608 477 644 645 cell_1rw
* cell instance $29856 m0 *1 144.525,131.04
X$29856 476 610 477 644 645 cell_1rw
* cell instance $29857 r0 *1 144.525,131.04
X$29857 476 611 477 644 645 cell_1rw
* cell instance $29858 m0 *1 144.525,133.77
X$29858 476 612 477 644 645 cell_1rw
* cell instance $29859 m0 *1 144.525,136.5
X$29859 476 615 477 644 645 cell_1rw
* cell instance $29860 r0 *1 144.525,133.77
X$29860 476 613 477 644 645 cell_1rw
* cell instance $29861 r0 *1 144.525,136.5
X$29861 476 614 477 644 645 cell_1rw
* cell instance $29862 m0 *1 144.525,139.23
X$29862 476 617 477 644 645 cell_1rw
* cell instance $29863 r0 *1 144.525,139.23
X$29863 476 616 477 644 645 cell_1rw
* cell instance $29864 m0 *1 144.525,141.96
X$29864 476 618 477 644 645 cell_1rw
* cell instance $29865 m0 *1 144.525,144.69
X$29865 476 620 477 644 645 cell_1rw
* cell instance $29866 r0 *1 144.525,141.96
X$29866 476 619 477 644 645 cell_1rw
* cell instance $29867 r0 *1 144.525,144.69
X$29867 476 621 477 644 645 cell_1rw
* cell instance $29868 m0 *1 144.525,147.42
X$29868 476 622 477 644 645 cell_1rw
* cell instance $29869 r0 *1 144.525,147.42
X$29869 476 623 477 644 645 cell_1rw
* cell instance $29870 m0 *1 144.525,150.15
X$29870 476 624 477 644 645 cell_1rw
* cell instance $29871 m0 *1 144.525,152.88
X$29871 476 626 477 644 645 cell_1rw
* cell instance $29872 r0 *1 144.525,150.15
X$29872 476 625 477 644 645 cell_1rw
* cell instance $29873 r0 *1 144.525,152.88
X$29873 476 627 477 644 645 cell_1rw
* cell instance $29874 m0 *1 144.525,155.61
X$29874 476 628 477 644 645 cell_1rw
* cell instance $29875 r0 *1 144.525,155.61
X$29875 476 629 477 644 645 cell_1rw
* cell instance $29876 m0 *1 144.525,158.34
X$29876 476 630 477 644 645 cell_1rw
* cell instance $29877 r0 *1 144.525,158.34
X$29877 476 631 477 644 645 cell_1rw
* cell instance $29878 m0 *1 144.525,161.07
X$29878 476 632 477 644 645 cell_1rw
* cell instance $29879 r0 *1 144.525,161.07
X$29879 476 633 477 644 645 cell_1rw
* cell instance $29880 m0 *1 144.525,163.8
X$29880 476 634 477 644 645 cell_1rw
* cell instance $29881 r0 *1 144.525,163.8
X$29881 476 635 477 644 645 cell_1rw
* cell instance $29882 m0 *1 144.525,166.53
X$29882 476 637 477 644 645 cell_1rw
* cell instance $29883 r0 *1 144.525,166.53
X$29883 476 636 477 644 645 cell_1rw
* cell instance $29884 m0 *1 144.525,169.26
X$29884 476 639 477 644 645 cell_1rw
* cell instance $29885 r0 *1 144.525,169.26
X$29885 476 638 477 644 645 cell_1rw
* cell instance $29886 m0 *1 144.525,171.99
X$29886 476 640 477 644 645 cell_1rw
* cell instance $29887 r0 *1 144.525,171.99
X$29887 476 641 477 644 645 cell_1rw
* cell instance $29888 m0 *1 144.525,174.72
X$29888 476 642 477 644 645 cell_1rw
* cell instance $29889 r0 *1 144.525,174.72
X$29889 476 643 477 644 645 cell_1rw
* cell instance $29890 m0 *1 145.23,90.09
X$29890 478 581 479 644 645 cell_1rw
* cell instance $29891 m0 *1 145.23,92.82
X$29891 478 583 479 644 645 cell_1rw
* cell instance $29892 r0 *1 145.23,90.09
X$29892 478 580 479 644 645 cell_1rw
* cell instance $29893 r0 *1 145.23,92.82
X$29893 478 582 479 644 645 cell_1rw
* cell instance $29894 m0 *1 145.23,95.55
X$29894 478 584 479 644 645 cell_1rw
* cell instance $29895 r0 *1 145.23,95.55
X$29895 478 585 479 644 645 cell_1rw
* cell instance $29896 m0 *1 145.23,98.28
X$29896 478 586 479 644 645 cell_1rw
* cell instance $29897 r0 *1 145.23,98.28
X$29897 478 587 479 644 645 cell_1rw
* cell instance $29898 m0 *1 145.23,101.01
X$29898 478 588 479 644 645 cell_1rw
* cell instance $29899 r0 *1 145.23,101.01
X$29899 478 589 479 644 645 cell_1rw
* cell instance $29900 m0 *1 145.23,103.74
X$29900 478 590 479 644 645 cell_1rw
* cell instance $29901 m0 *1 145.23,106.47
X$29901 478 593 479 644 645 cell_1rw
* cell instance $29902 r0 *1 145.23,103.74
X$29902 478 591 479 644 645 cell_1rw
* cell instance $29903 r0 *1 145.23,106.47
X$29903 478 592 479 644 645 cell_1rw
* cell instance $29904 m0 *1 145.23,109.2
X$29904 478 594 479 644 645 cell_1rw
* cell instance $29905 m0 *1 145.23,111.93
X$29905 478 597 479 644 645 cell_1rw
* cell instance $29906 r0 *1 145.23,109.2
X$29906 478 595 479 644 645 cell_1rw
* cell instance $29907 m0 *1 145.23,114.66
X$29907 478 598 479 644 645 cell_1rw
* cell instance $29908 r0 *1 145.23,111.93
X$29908 478 596 479 644 645 cell_1rw
* cell instance $29909 r0 *1 145.23,114.66
X$29909 478 599 479 644 645 cell_1rw
* cell instance $29910 m0 *1 145.23,117.39
X$29910 478 600 479 644 645 cell_1rw
* cell instance $29911 r0 *1 145.23,117.39
X$29911 478 601 479 644 645 cell_1rw
* cell instance $29912 m0 *1 145.23,120.12
X$29912 478 602 479 644 645 cell_1rw
* cell instance $29913 r0 *1 145.23,120.12
X$29913 478 603 479 644 645 cell_1rw
* cell instance $29914 m0 *1 145.23,122.85
X$29914 478 604 479 644 645 cell_1rw
* cell instance $29915 r0 *1 145.23,122.85
X$29915 478 605 479 644 645 cell_1rw
* cell instance $29916 m0 *1 145.23,125.58
X$29916 478 606 479 644 645 cell_1rw
* cell instance $29917 r0 *1 145.23,125.58
X$29917 478 607 479 644 645 cell_1rw
* cell instance $29918 m0 *1 145.23,128.31
X$29918 478 609 479 644 645 cell_1rw
* cell instance $29919 r0 *1 145.23,128.31
X$29919 478 608 479 644 645 cell_1rw
* cell instance $29920 m0 *1 145.23,131.04
X$29920 478 610 479 644 645 cell_1rw
* cell instance $29921 r0 *1 145.23,131.04
X$29921 478 611 479 644 645 cell_1rw
* cell instance $29922 m0 *1 145.23,133.77
X$29922 478 612 479 644 645 cell_1rw
* cell instance $29923 r0 *1 145.23,133.77
X$29923 478 613 479 644 645 cell_1rw
* cell instance $29924 m0 *1 145.23,136.5
X$29924 478 615 479 644 645 cell_1rw
* cell instance $29925 r0 *1 145.23,136.5
X$29925 478 614 479 644 645 cell_1rw
* cell instance $29926 m0 *1 145.23,139.23
X$29926 478 617 479 644 645 cell_1rw
* cell instance $29927 r0 *1 145.23,139.23
X$29927 478 616 479 644 645 cell_1rw
* cell instance $29928 m0 *1 145.23,141.96
X$29928 478 618 479 644 645 cell_1rw
* cell instance $29929 r0 *1 145.23,141.96
X$29929 478 619 479 644 645 cell_1rw
* cell instance $29930 m0 *1 145.23,144.69
X$29930 478 620 479 644 645 cell_1rw
* cell instance $29931 r0 *1 145.23,144.69
X$29931 478 621 479 644 645 cell_1rw
* cell instance $29932 m0 *1 145.23,147.42
X$29932 478 622 479 644 645 cell_1rw
* cell instance $29933 m0 *1 145.23,150.15
X$29933 478 624 479 644 645 cell_1rw
* cell instance $29934 r0 *1 145.23,147.42
X$29934 478 623 479 644 645 cell_1rw
* cell instance $29935 r0 *1 145.23,150.15
X$29935 478 625 479 644 645 cell_1rw
* cell instance $29936 m0 *1 145.23,152.88
X$29936 478 626 479 644 645 cell_1rw
* cell instance $29937 r0 *1 145.23,152.88
X$29937 478 627 479 644 645 cell_1rw
* cell instance $29938 m0 *1 145.23,155.61
X$29938 478 628 479 644 645 cell_1rw
* cell instance $29939 r0 *1 145.23,155.61
X$29939 478 629 479 644 645 cell_1rw
* cell instance $29940 m0 *1 145.23,158.34
X$29940 478 630 479 644 645 cell_1rw
* cell instance $29941 r0 *1 145.23,158.34
X$29941 478 631 479 644 645 cell_1rw
* cell instance $29942 m0 *1 145.23,161.07
X$29942 478 632 479 644 645 cell_1rw
* cell instance $29943 r0 *1 145.23,161.07
X$29943 478 633 479 644 645 cell_1rw
* cell instance $29944 m0 *1 145.23,163.8
X$29944 478 634 479 644 645 cell_1rw
* cell instance $29945 r0 *1 145.23,163.8
X$29945 478 635 479 644 645 cell_1rw
* cell instance $29946 m0 *1 145.23,166.53
X$29946 478 637 479 644 645 cell_1rw
* cell instance $29947 r0 *1 145.23,166.53
X$29947 478 636 479 644 645 cell_1rw
* cell instance $29948 m0 *1 145.23,169.26
X$29948 478 639 479 644 645 cell_1rw
* cell instance $29949 r0 *1 145.23,169.26
X$29949 478 638 479 644 645 cell_1rw
* cell instance $29950 m0 *1 145.23,171.99
X$29950 478 640 479 644 645 cell_1rw
* cell instance $29951 r0 *1 145.23,171.99
X$29951 478 641 479 644 645 cell_1rw
* cell instance $29952 m0 *1 145.23,174.72
X$29952 478 642 479 644 645 cell_1rw
* cell instance $29953 r0 *1 145.23,174.72
X$29953 478 643 479 644 645 cell_1rw
* cell instance $29954 m0 *1 145.935,90.09
X$29954 480 581 481 644 645 cell_1rw
* cell instance $29955 m0 *1 145.935,92.82
X$29955 480 583 481 644 645 cell_1rw
* cell instance $29956 r0 *1 145.935,90.09
X$29956 480 580 481 644 645 cell_1rw
* cell instance $29957 r0 *1 145.935,92.82
X$29957 480 582 481 644 645 cell_1rw
* cell instance $29958 m0 *1 145.935,95.55
X$29958 480 584 481 644 645 cell_1rw
* cell instance $29959 r0 *1 145.935,95.55
X$29959 480 585 481 644 645 cell_1rw
* cell instance $29960 m0 *1 145.935,98.28
X$29960 480 586 481 644 645 cell_1rw
* cell instance $29961 r0 *1 145.935,98.28
X$29961 480 587 481 644 645 cell_1rw
* cell instance $29962 m0 *1 145.935,101.01
X$29962 480 588 481 644 645 cell_1rw
* cell instance $29963 m0 *1 145.935,103.74
X$29963 480 590 481 644 645 cell_1rw
* cell instance $29964 r0 *1 145.935,101.01
X$29964 480 589 481 644 645 cell_1rw
* cell instance $29965 r0 *1 145.935,103.74
X$29965 480 591 481 644 645 cell_1rw
* cell instance $29966 m0 *1 145.935,106.47
X$29966 480 593 481 644 645 cell_1rw
* cell instance $29967 r0 *1 145.935,106.47
X$29967 480 592 481 644 645 cell_1rw
* cell instance $29968 m0 *1 145.935,109.2
X$29968 480 594 481 644 645 cell_1rw
* cell instance $29969 r0 *1 145.935,109.2
X$29969 480 595 481 644 645 cell_1rw
* cell instance $29970 m0 *1 145.935,111.93
X$29970 480 597 481 644 645 cell_1rw
* cell instance $29971 r0 *1 145.935,111.93
X$29971 480 596 481 644 645 cell_1rw
* cell instance $29972 m0 *1 145.935,114.66
X$29972 480 598 481 644 645 cell_1rw
* cell instance $29973 r0 *1 145.935,114.66
X$29973 480 599 481 644 645 cell_1rw
* cell instance $29974 m0 *1 145.935,117.39
X$29974 480 600 481 644 645 cell_1rw
* cell instance $29975 r0 *1 145.935,117.39
X$29975 480 601 481 644 645 cell_1rw
* cell instance $29976 m0 *1 145.935,120.12
X$29976 480 602 481 644 645 cell_1rw
* cell instance $29977 r0 *1 145.935,120.12
X$29977 480 603 481 644 645 cell_1rw
* cell instance $29978 m0 *1 145.935,122.85
X$29978 480 604 481 644 645 cell_1rw
* cell instance $29979 r0 *1 145.935,122.85
X$29979 480 605 481 644 645 cell_1rw
* cell instance $29980 m0 *1 145.935,125.58
X$29980 480 606 481 644 645 cell_1rw
* cell instance $29981 r0 *1 145.935,125.58
X$29981 480 607 481 644 645 cell_1rw
* cell instance $29982 m0 *1 145.935,128.31
X$29982 480 609 481 644 645 cell_1rw
* cell instance $29983 r0 *1 145.935,128.31
X$29983 480 608 481 644 645 cell_1rw
* cell instance $29984 m0 *1 145.935,131.04
X$29984 480 610 481 644 645 cell_1rw
* cell instance $29985 r0 *1 145.935,131.04
X$29985 480 611 481 644 645 cell_1rw
* cell instance $29986 m0 *1 145.935,133.77
X$29986 480 612 481 644 645 cell_1rw
* cell instance $29987 r0 *1 145.935,133.77
X$29987 480 613 481 644 645 cell_1rw
* cell instance $29988 m0 *1 145.935,136.5
X$29988 480 615 481 644 645 cell_1rw
* cell instance $29989 r0 *1 145.935,136.5
X$29989 480 614 481 644 645 cell_1rw
* cell instance $29990 m0 *1 145.935,139.23
X$29990 480 617 481 644 645 cell_1rw
* cell instance $29991 r0 *1 145.935,139.23
X$29991 480 616 481 644 645 cell_1rw
* cell instance $29992 m0 *1 145.935,141.96
X$29992 480 618 481 644 645 cell_1rw
* cell instance $29993 r0 *1 145.935,141.96
X$29993 480 619 481 644 645 cell_1rw
* cell instance $29994 m0 *1 145.935,144.69
X$29994 480 620 481 644 645 cell_1rw
* cell instance $29995 r0 *1 145.935,144.69
X$29995 480 621 481 644 645 cell_1rw
* cell instance $29996 m0 *1 145.935,147.42
X$29996 480 622 481 644 645 cell_1rw
* cell instance $29997 r0 *1 145.935,147.42
X$29997 480 623 481 644 645 cell_1rw
* cell instance $29998 m0 *1 145.935,150.15
X$29998 480 624 481 644 645 cell_1rw
* cell instance $29999 r0 *1 145.935,150.15
X$29999 480 625 481 644 645 cell_1rw
* cell instance $30000 m0 *1 145.935,152.88
X$30000 480 626 481 644 645 cell_1rw
* cell instance $30001 r0 *1 145.935,152.88
X$30001 480 627 481 644 645 cell_1rw
* cell instance $30002 m0 *1 145.935,155.61
X$30002 480 628 481 644 645 cell_1rw
* cell instance $30003 r0 *1 145.935,155.61
X$30003 480 629 481 644 645 cell_1rw
* cell instance $30004 m0 *1 145.935,158.34
X$30004 480 630 481 644 645 cell_1rw
* cell instance $30005 r0 *1 145.935,158.34
X$30005 480 631 481 644 645 cell_1rw
* cell instance $30006 m0 *1 145.935,161.07
X$30006 480 632 481 644 645 cell_1rw
* cell instance $30007 m0 *1 145.935,163.8
X$30007 480 634 481 644 645 cell_1rw
* cell instance $30008 r0 *1 145.935,161.07
X$30008 480 633 481 644 645 cell_1rw
* cell instance $30009 m0 *1 145.935,166.53
X$30009 480 637 481 644 645 cell_1rw
* cell instance $30010 r0 *1 145.935,163.8
X$30010 480 635 481 644 645 cell_1rw
* cell instance $30011 m0 *1 145.935,169.26
X$30011 480 639 481 644 645 cell_1rw
* cell instance $30012 r0 *1 145.935,166.53
X$30012 480 636 481 644 645 cell_1rw
* cell instance $30013 r0 *1 145.935,169.26
X$30013 480 638 481 644 645 cell_1rw
* cell instance $30014 m0 *1 145.935,171.99
X$30014 480 640 481 644 645 cell_1rw
* cell instance $30015 r0 *1 145.935,171.99
X$30015 480 641 481 644 645 cell_1rw
* cell instance $30016 m0 *1 145.935,174.72
X$30016 480 642 481 644 645 cell_1rw
* cell instance $30017 r0 *1 145.935,174.72
X$30017 480 643 481 644 645 cell_1rw
* cell instance $30018 m0 *1 146.64,90.09
X$30018 482 581 483 644 645 cell_1rw
* cell instance $30019 r0 *1 146.64,90.09
X$30019 482 580 483 644 645 cell_1rw
* cell instance $30020 m0 *1 146.64,92.82
X$30020 482 583 483 644 645 cell_1rw
* cell instance $30021 r0 *1 146.64,92.82
X$30021 482 582 483 644 645 cell_1rw
* cell instance $30022 m0 *1 146.64,95.55
X$30022 482 584 483 644 645 cell_1rw
* cell instance $30023 r0 *1 146.64,95.55
X$30023 482 585 483 644 645 cell_1rw
* cell instance $30024 m0 *1 146.64,98.28
X$30024 482 586 483 644 645 cell_1rw
* cell instance $30025 r0 *1 146.64,98.28
X$30025 482 587 483 644 645 cell_1rw
* cell instance $30026 m0 *1 146.64,101.01
X$30026 482 588 483 644 645 cell_1rw
* cell instance $30027 r0 *1 146.64,101.01
X$30027 482 589 483 644 645 cell_1rw
* cell instance $30028 m0 *1 146.64,103.74
X$30028 482 590 483 644 645 cell_1rw
* cell instance $30029 r0 *1 146.64,103.74
X$30029 482 591 483 644 645 cell_1rw
* cell instance $30030 m0 *1 146.64,106.47
X$30030 482 593 483 644 645 cell_1rw
* cell instance $30031 r0 *1 146.64,106.47
X$30031 482 592 483 644 645 cell_1rw
* cell instance $30032 m0 *1 146.64,109.2
X$30032 482 594 483 644 645 cell_1rw
* cell instance $30033 m0 *1 146.64,111.93
X$30033 482 597 483 644 645 cell_1rw
* cell instance $30034 r0 *1 146.64,109.2
X$30034 482 595 483 644 645 cell_1rw
* cell instance $30035 r0 *1 146.64,111.93
X$30035 482 596 483 644 645 cell_1rw
* cell instance $30036 m0 *1 146.64,114.66
X$30036 482 598 483 644 645 cell_1rw
* cell instance $30037 r0 *1 146.64,114.66
X$30037 482 599 483 644 645 cell_1rw
* cell instance $30038 m0 *1 146.64,117.39
X$30038 482 600 483 644 645 cell_1rw
* cell instance $30039 r0 *1 146.64,117.39
X$30039 482 601 483 644 645 cell_1rw
* cell instance $30040 m0 *1 146.64,120.12
X$30040 482 602 483 644 645 cell_1rw
* cell instance $30041 r0 *1 146.64,120.12
X$30041 482 603 483 644 645 cell_1rw
* cell instance $30042 m0 *1 146.64,122.85
X$30042 482 604 483 644 645 cell_1rw
* cell instance $30043 m0 *1 146.64,125.58
X$30043 482 606 483 644 645 cell_1rw
* cell instance $30044 r0 *1 146.64,122.85
X$30044 482 605 483 644 645 cell_1rw
* cell instance $30045 r0 *1 146.64,125.58
X$30045 482 607 483 644 645 cell_1rw
* cell instance $30046 m0 *1 146.64,128.31
X$30046 482 609 483 644 645 cell_1rw
* cell instance $30047 m0 *1 146.64,131.04
X$30047 482 610 483 644 645 cell_1rw
* cell instance $30048 r0 *1 146.64,128.31
X$30048 482 608 483 644 645 cell_1rw
* cell instance $30049 m0 *1 146.64,133.77
X$30049 482 612 483 644 645 cell_1rw
* cell instance $30050 r0 *1 146.64,131.04
X$30050 482 611 483 644 645 cell_1rw
* cell instance $30051 m0 *1 146.64,136.5
X$30051 482 615 483 644 645 cell_1rw
* cell instance $30052 r0 *1 146.64,133.77
X$30052 482 613 483 644 645 cell_1rw
* cell instance $30053 r0 *1 146.64,136.5
X$30053 482 614 483 644 645 cell_1rw
* cell instance $30054 m0 *1 146.64,139.23
X$30054 482 617 483 644 645 cell_1rw
* cell instance $30055 r0 *1 146.64,139.23
X$30055 482 616 483 644 645 cell_1rw
* cell instance $30056 m0 *1 146.64,141.96
X$30056 482 618 483 644 645 cell_1rw
* cell instance $30057 r0 *1 146.64,141.96
X$30057 482 619 483 644 645 cell_1rw
* cell instance $30058 m0 *1 146.64,144.69
X$30058 482 620 483 644 645 cell_1rw
* cell instance $30059 m0 *1 146.64,147.42
X$30059 482 622 483 644 645 cell_1rw
* cell instance $30060 r0 *1 146.64,144.69
X$30060 482 621 483 644 645 cell_1rw
* cell instance $30061 m0 *1 146.64,150.15
X$30061 482 624 483 644 645 cell_1rw
* cell instance $30062 r0 *1 146.64,147.42
X$30062 482 623 483 644 645 cell_1rw
* cell instance $30063 m0 *1 146.64,152.88
X$30063 482 626 483 644 645 cell_1rw
* cell instance $30064 r0 *1 146.64,150.15
X$30064 482 625 483 644 645 cell_1rw
* cell instance $30065 r0 *1 146.64,152.88
X$30065 482 627 483 644 645 cell_1rw
* cell instance $30066 m0 *1 146.64,155.61
X$30066 482 628 483 644 645 cell_1rw
* cell instance $30067 r0 *1 146.64,155.61
X$30067 482 629 483 644 645 cell_1rw
* cell instance $30068 m0 *1 146.64,158.34
X$30068 482 630 483 644 645 cell_1rw
* cell instance $30069 r0 *1 146.64,158.34
X$30069 482 631 483 644 645 cell_1rw
* cell instance $30070 m0 *1 146.64,161.07
X$30070 482 632 483 644 645 cell_1rw
* cell instance $30071 r0 *1 146.64,161.07
X$30071 482 633 483 644 645 cell_1rw
* cell instance $30072 m0 *1 146.64,163.8
X$30072 482 634 483 644 645 cell_1rw
* cell instance $30073 r0 *1 146.64,163.8
X$30073 482 635 483 644 645 cell_1rw
* cell instance $30074 m0 *1 146.64,166.53
X$30074 482 637 483 644 645 cell_1rw
* cell instance $30075 r0 *1 146.64,166.53
X$30075 482 636 483 644 645 cell_1rw
* cell instance $30076 m0 *1 146.64,169.26
X$30076 482 639 483 644 645 cell_1rw
* cell instance $30077 r0 *1 146.64,169.26
X$30077 482 638 483 644 645 cell_1rw
* cell instance $30078 m0 *1 146.64,171.99
X$30078 482 640 483 644 645 cell_1rw
* cell instance $30079 m0 *1 146.64,174.72
X$30079 482 642 483 644 645 cell_1rw
* cell instance $30080 r0 *1 146.64,171.99
X$30080 482 641 483 644 645 cell_1rw
* cell instance $30081 r0 *1 146.64,174.72
X$30081 482 643 483 644 645 cell_1rw
* cell instance $30082 m0 *1 147.345,90.09
X$30082 484 581 485 644 645 cell_1rw
* cell instance $30083 r0 *1 147.345,90.09
X$30083 484 580 485 644 645 cell_1rw
* cell instance $30084 m0 *1 147.345,92.82
X$30084 484 583 485 644 645 cell_1rw
* cell instance $30085 r0 *1 147.345,92.82
X$30085 484 582 485 644 645 cell_1rw
* cell instance $30086 m0 *1 147.345,95.55
X$30086 484 584 485 644 645 cell_1rw
* cell instance $30087 r0 *1 147.345,95.55
X$30087 484 585 485 644 645 cell_1rw
* cell instance $30088 m0 *1 147.345,98.28
X$30088 484 586 485 644 645 cell_1rw
* cell instance $30089 r0 *1 147.345,98.28
X$30089 484 587 485 644 645 cell_1rw
* cell instance $30090 m0 *1 147.345,101.01
X$30090 484 588 485 644 645 cell_1rw
* cell instance $30091 r0 *1 147.345,101.01
X$30091 484 589 485 644 645 cell_1rw
* cell instance $30092 m0 *1 147.345,103.74
X$30092 484 590 485 644 645 cell_1rw
* cell instance $30093 r0 *1 147.345,103.74
X$30093 484 591 485 644 645 cell_1rw
* cell instance $30094 m0 *1 147.345,106.47
X$30094 484 593 485 644 645 cell_1rw
* cell instance $30095 r0 *1 147.345,106.47
X$30095 484 592 485 644 645 cell_1rw
* cell instance $30096 m0 *1 147.345,109.2
X$30096 484 594 485 644 645 cell_1rw
* cell instance $30097 m0 *1 147.345,111.93
X$30097 484 597 485 644 645 cell_1rw
* cell instance $30098 r0 *1 147.345,109.2
X$30098 484 595 485 644 645 cell_1rw
* cell instance $30099 r0 *1 147.345,111.93
X$30099 484 596 485 644 645 cell_1rw
* cell instance $30100 m0 *1 147.345,114.66
X$30100 484 598 485 644 645 cell_1rw
* cell instance $30101 r0 *1 147.345,114.66
X$30101 484 599 485 644 645 cell_1rw
* cell instance $30102 m0 *1 147.345,117.39
X$30102 484 600 485 644 645 cell_1rw
* cell instance $30103 r0 *1 147.345,117.39
X$30103 484 601 485 644 645 cell_1rw
* cell instance $30104 m0 *1 147.345,120.12
X$30104 484 602 485 644 645 cell_1rw
* cell instance $30105 m0 *1 147.345,122.85
X$30105 484 604 485 644 645 cell_1rw
* cell instance $30106 r0 *1 147.345,120.12
X$30106 484 603 485 644 645 cell_1rw
* cell instance $30107 r0 *1 147.345,122.85
X$30107 484 605 485 644 645 cell_1rw
* cell instance $30108 m0 *1 147.345,125.58
X$30108 484 606 485 644 645 cell_1rw
* cell instance $30109 m0 *1 147.345,128.31
X$30109 484 609 485 644 645 cell_1rw
* cell instance $30110 r0 *1 147.345,125.58
X$30110 484 607 485 644 645 cell_1rw
* cell instance $30111 m0 *1 147.345,131.04
X$30111 484 610 485 644 645 cell_1rw
* cell instance $30112 r0 *1 147.345,128.31
X$30112 484 608 485 644 645 cell_1rw
* cell instance $30113 m0 *1 147.345,133.77
X$30113 484 612 485 644 645 cell_1rw
* cell instance $30114 r0 *1 147.345,131.04
X$30114 484 611 485 644 645 cell_1rw
* cell instance $30115 r0 *1 147.345,133.77
X$30115 484 613 485 644 645 cell_1rw
* cell instance $30116 m0 *1 147.345,136.5
X$30116 484 615 485 644 645 cell_1rw
* cell instance $30117 r0 *1 147.345,136.5
X$30117 484 614 485 644 645 cell_1rw
* cell instance $30118 m0 *1 147.345,139.23
X$30118 484 617 485 644 645 cell_1rw
* cell instance $30119 r0 *1 147.345,139.23
X$30119 484 616 485 644 645 cell_1rw
* cell instance $30120 m0 *1 147.345,141.96
X$30120 484 618 485 644 645 cell_1rw
* cell instance $30121 m0 *1 147.345,144.69
X$30121 484 620 485 644 645 cell_1rw
* cell instance $30122 r0 *1 147.345,141.96
X$30122 484 619 485 644 645 cell_1rw
* cell instance $30123 r0 *1 147.345,144.69
X$30123 484 621 485 644 645 cell_1rw
* cell instance $30124 m0 *1 147.345,147.42
X$30124 484 622 485 644 645 cell_1rw
* cell instance $30125 m0 *1 147.345,150.15
X$30125 484 624 485 644 645 cell_1rw
* cell instance $30126 r0 *1 147.345,147.42
X$30126 484 623 485 644 645 cell_1rw
* cell instance $30127 r0 *1 147.345,150.15
X$30127 484 625 485 644 645 cell_1rw
* cell instance $30128 m0 *1 147.345,152.88
X$30128 484 626 485 644 645 cell_1rw
* cell instance $30129 r0 *1 147.345,152.88
X$30129 484 627 485 644 645 cell_1rw
* cell instance $30130 m0 *1 147.345,155.61
X$30130 484 628 485 644 645 cell_1rw
* cell instance $30131 r0 *1 147.345,155.61
X$30131 484 629 485 644 645 cell_1rw
* cell instance $30132 m0 *1 147.345,158.34
X$30132 484 630 485 644 645 cell_1rw
* cell instance $30133 m0 *1 147.345,161.07
X$30133 484 632 485 644 645 cell_1rw
* cell instance $30134 r0 *1 147.345,158.34
X$30134 484 631 485 644 645 cell_1rw
* cell instance $30135 r0 *1 147.345,161.07
X$30135 484 633 485 644 645 cell_1rw
* cell instance $30136 m0 *1 147.345,163.8
X$30136 484 634 485 644 645 cell_1rw
* cell instance $30137 r0 *1 147.345,163.8
X$30137 484 635 485 644 645 cell_1rw
* cell instance $30138 m0 *1 147.345,166.53
X$30138 484 637 485 644 645 cell_1rw
* cell instance $30139 r0 *1 147.345,166.53
X$30139 484 636 485 644 645 cell_1rw
* cell instance $30140 m0 *1 147.345,169.26
X$30140 484 639 485 644 645 cell_1rw
* cell instance $30141 r0 *1 147.345,169.26
X$30141 484 638 485 644 645 cell_1rw
* cell instance $30142 m0 *1 147.345,171.99
X$30142 484 640 485 644 645 cell_1rw
* cell instance $30143 r0 *1 147.345,171.99
X$30143 484 641 485 644 645 cell_1rw
* cell instance $30144 m0 *1 147.345,174.72
X$30144 484 642 485 644 645 cell_1rw
* cell instance $30145 r0 *1 147.345,174.72
X$30145 484 643 485 644 645 cell_1rw
* cell instance $30146 m0 *1 148.05,90.09
X$30146 486 581 487 644 645 cell_1rw
* cell instance $30147 r0 *1 148.05,90.09
X$30147 486 580 487 644 645 cell_1rw
* cell instance $30148 m0 *1 148.05,92.82
X$30148 486 583 487 644 645 cell_1rw
* cell instance $30149 r0 *1 148.05,92.82
X$30149 486 582 487 644 645 cell_1rw
* cell instance $30150 m0 *1 148.05,95.55
X$30150 486 584 487 644 645 cell_1rw
* cell instance $30151 r0 *1 148.05,95.55
X$30151 486 585 487 644 645 cell_1rw
* cell instance $30152 m0 *1 148.05,98.28
X$30152 486 586 487 644 645 cell_1rw
* cell instance $30153 r0 *1 148.05,98.28
X$30153 486 587 487 644 645 cell_1rw
* cell instance $30154 m0 *1 148.05,101.01
X$30154 486 588 487 644 645 cell_1rw
* cell instance $30155 r0 *1 148.05,101.01
X$30155 486 589 487 644 645 cell_1rw
* cell instance $30156 m0 *1 148.05,103.74
X$30156 486 590 487 644 645 cell_1rw
* cell instance $30157 r0 *1 148.05,103.74
X$30157 486 591 487 644 645 cell_1rw
* cell instance $30158 m0 *1 148.05,106.47
X$30158 486 593 487 644 645 cell_1rw
* cell instance $30159 r0 *1 148.05,106.47
X$30159 486 592 487 644 645 cell_1rw
* cell instance $30160 m0 *1 148.05,109.2
X$30160 486 594 487 644 645 cell_1rw
* cell instance $30161 r0 *1 148.05,109.2
X$30161 486 595 487 644 645 cell_1rw
* cell instance $30162 m0 *1 148.05,111.93
X$30162 486 597 487 644 645 cell_1rw
* cell instance $30163 m0 *1 148.05,114.66
X$30163 486 598 487 644 645 cell_1rw
* cell instance $30164 r0 *1 148.05,111.93
X$30164 486 596 487 644 645 cell_1rw
* cell instance $30165 r0 *1 148.05,114.66
X$30165 486 599 487 644 645 cell_1rw
* cell instance $30166 m0 *1 148.05,117.39
X$30166 486 600 487 644 645 cell_1rw
* cell instance $30167 r0 *1 148.05,117.39
X$30167 486 601 487 644 645 cell_1rw
* cell instance $30168 m0 *1 148.05,120.12
X$30168 486 602 487 644 645 cell_1rw
* cell instance $30169 r0 *1 148.05,120.12
X$30169 486 603 487 644 645 cell_1rw
* cell instance $30170 m0 *1 148.05,122.85
X$30170 486 604 487 644 645 cell_1rw
* cell instance $30171 r0 *1 148.05,122.85
X$30171 486 605 487 644 645 cell_1rw
* cell instance $30172 m0 *1 148.05,125.58
X$30172 486 606 487 644 645 cell_1rw
* cell instance $30173 m0 *1 148.05,128.31
X$30173 486 609 487 644 645 cell_1rw
* cell instance $30174 r0 *1 148.05,125.58
X$30174 486 607 487 644 645 cell_1rw
* cell instance $30175 r0 *1 148.05,128.31
X$30175 486 608 487 644 645 cell_1rw
* cell instance $30176 m0 *1 148.05,131.04
X$30176 486 610 487 644 645 cell_1rw
* cell instance $30177 m0 *1 148.05,133.77
X$30177 486 612 487 644 645 cell_1rw
* cell instance $30178 r0 *1 148.05,131.04
X$30178 486 611 487 644 645 cell_1rw
* cell instance $30179 r0 *1 148.05,133.77
X$30179 486 613 487 644 645 cell_1rw
* cell instance $30180 m0 *1 148.05,136.5
X$30180 486 615 487 644 645 cell_1rw
* cell instance $30181 r0 *1 148.05,136.5
X$30181 486 614 487 644 645 cell_1rw
* cell instance $30182 m0 *1 148.05,139.23
X$30182 486 617 487 644 645 cell_1rw
* cell instance $30183 m0 *1 148.05,141.96
X$30183 486 618 487 644 645 cell_1rw
* cell instance $30184 r0 *1 148.05,139.23
X$30184 486 616 487 644 645 cell_1rw
* cell instance $30185 r0 *1 148.05,141.96
X$30185 486 619 487 644 645 cell_1rw
* cell instance $30186 m0 *1 148.05,144.69
X$30186 486 620 487 644 645 cell_1rw
* cell instance $30187 r0 *1 148.05,144.69
X$30187 486 621 487 644 645 cell_1rw
* cell instance $30188 m0 *1 148.05,147.42
X$30188 486 622 487 644 645 cell_1rw
* cell instance $30189 r0 *1 148.05,147.42
X$30189 486 623 487 644 645 cell_1rw
* cell instance $30190 m0 *1 148.05,150.15
X$30190 486 624 487 644 645 cell_1rw
* cell instance $30191 r0 *1 148.05,150.15
X$30191 486 625 487 644 645 cell_1rw
* cell instance $30192 m0 *1 148.05,152.88
X$30192 486 626 487 644 645 cell_1rw
* cell instance $30193 r0 *1 148.05,152.88
X$30193 486 627 487 644 645 cell_1rw
* cell instance $30194 m0 *1 148.05,155.61
X$30194 486 628 487 644 645 cell_1rw
* cell instance $30195 m0 *1 148.05,158.34
X$30195 486 630 487 644 645 cell_1rw
* cell instance $30196 r0 *1 148.05,155.61
X$30196 486 629 487 644 645 cell_1rw
* cell instance $30197 r0 *1 148.05,158.34
X$30197 486 631 487 644 645 cell_1rw
* cell instance $30198 m0 *1 148.05,161.07
X$30198 486 632 487 644 645 cell_1rw
* cell instance $30199 m0 *1 148.05,163.8
X$30199 486 634 487 644 645 cell_1rw
* cell instance $30200 r0 *1 148.05,161.07
X$30200 486 633 487 644 645 cell_1rw
* cell instance $30201 r0 *1 148.05,163.8
X$30201 486 635 487 644 645 cell_1rw
* cell instance $30202 m0 *1 148.05,166.53
X$30202 486 637 487 644 645 cell_1rw
* cell instance $30203 r0 *1 148.05,166.53
X$30203 486 636 487 644 645 cell_1rw
* cell instance $30204 m0 *1 148.05,169.26
X$30204 486 639 487 644 645 cell_1rw
* cell instance $30205 r0 *1 148.05,169.26
X$30205 486 638 487 644 645 cell_1rw
* cell instance $30206 m0 *1 148.05,171.99
X$30206 486 640 487 644 645 cell_1rw
* cell instance $30207 r0 *1 148.05,171.99
X$30207 486 641 487 644 645 cell_1rw
* cell instance $30208 m0 *1 148.05,174.72
X$30208 486 642 487 644 645 cell_1rw
* cell instance $30209 r0 *1 148.05,174.72
X$30209 486 643 487 644 645 cell_1rw
* cell instance $30210 m0 *1 148.755,90.09
X$30210 488 581 489 644 645 cell_1rw
* cell instance $30211 r0 *1 148.755,90.09
X$30211 488 580 489 644 645 cell_1rw
* cell instance $30212 m0 *1 148.755,92.82
X$30212 488 583 489 644 645 cell_1rw
* cell instance $30213 r0 *1 148.755,92.82
X$30213 488 582 489 644 645 cell_1rw
* cell instance $30214 m0 *1 148.755,95.55
X$30214 488 584 489 644 645 cell_1rw
* cell instance $30215 m0 *1 148.755,98.28
X$30215 488 586 489 644 645 cell_1rw
* cell instance $30216 r0 *1 148.755,95.55
X$30216 488 585 489 644 645 cell_1rw
* cell instance $30217 r0 *1 148.755,98.28
X$30217 488 587 489 644 645 cell_1rw
* cell instance $30218 m0 *1 148.755,101.01
X$30218 488 588 489 644 645 cell_1rw
* cell instance $30219 m0 *1 148.755,103.74
X$30219 488 590 489 644 645 cell_1rw
* cell instance $30220 r0 *1 148.755,101.01
X$30220 488 589 489 644 645 cell_1rw
* cell instance $30221 r0 *1 148.755,103.74
X$30221 488 591 489 644 645 cell_1rw
* cell instance $30222 m0 *1 148.755,106.47
X$30222 488 593 489 644 645 cell_1rw
* cell instance $30223 r0 *1 148.755,106.47
X$30223 488 592 489 644 645 cell_1rw
* cell instance $30224 m0 *1 148.755,109.2
X$30224 488 594 489 644 645 cell_1rw
* cell instance $30225 r0 *1 148.755,109.2
X$30225 488 595 489 644 645 cell_1rw
* cell instance $30226 m0 *1 148.755,111.93
X$30226 488 597 489 644 645 cell_1rw
* cell instance $30227 m0 *1 148.755,114.66
X$30227 488 598 489 644 645 cell_1rw
* cell instance $30228 r0 *1 148.755,111.93
X$30228 488 596 489 644 645 cell_1rw
* cell instance $30229 r0 *1 148.755,114.66
X$30229 488 599 489 644 645 cell_1rw
* cell instance $30230 m0 *1 148.755,117.39
X$30230 488 600 489 644 645 cell_1rw
* cell instance $30231 m0 *1 148.755,120.12
X$30231 488 602 489 644 645 cell_1rw
* cell instance $30232 r0 *1 148.755,117.39
X$30232 488 601 489 644 645 cell_1rw
* cell instance $30233 m0 *1 148.755,122.85
X$30233 488 604 489 644 645 cell_1rw
* cell instance $30234 r0 *1 148.755,120.12
X$30234 488 603 489 644 645 cell_1rw
* cell instance $30235 r0 *1 148.755,122.85
X$30235 488 605 489 644 645 cell_1rw
* cell instance $30236 m0 *1 148.755,125.58
X$30236 488 606 489 644 645 cell_1rw
* cell instance $30237 r0 *1 148.755,125.58
X$30237 488 607 489 644 645 cell_1rw
* cell instance $30238 m0 *1 148.755,128.31
X$30238 488 609 489 644 645 cell_1rw
* cell instance $30239 r0 *1 148.755,128.31
X$30239 488 608 489 644 645 cell_1rw
* cell instance $30240 m0 *1 148.755,131.04
X$30240 488 610 489 644 645 cell_1rw
* cell instance $30241 r0 *1 148.755,131.04
X$30241 488 611 489 644 645 cell_1rw
* cell instance $30242 m0 *1 148.755,133.77
X$30242 488 612 489 644 645 cell_1rw
* cell instance $30243 r0 *1 148.755,133.77
X$30243 488 613 489 644 645 cell_1rw
* cell instance $30244 m0 *1 148.755,136.5
X$30244 488 615 489 644 645 cell_1rw
* cell instance $30245 r0 *1 148.755,136.5
X$30245 488 614 489 644 645 cell_1rw
* cell instance $30246 m0 *1 148.755,139.23
X$30246 488 617 489 644 645 cell_1rw
* cell instance $30247 r0 *1 148.755,139.23
X$30247 488 616 489 644 645 cell_1rw
* cell instance $30248 m0 *1 148.755,141.96
X$30248 488 618 489 644 645 cell_1rw
* cell instance $30249 m0 *1 148.755,144.69
X$30249 488 620 489 644 645 cell_1rw
* cell instance $30250 r0 *1 148.755,141.96
X$30250 488 619 489 644 645 cell_1rw
* cell instance $30251 r0 *1 148.755,144.69
X$30251 488 621 489 644 645 cell_1rw
* cell instance $30252 m0 *1 148.755,147.42
X$30252 488 622 489 644 645 cell_1rw
* cell instance $30253 m0 *1 148.755,150.15
X$30253 488 624 489 644 645 cell_1rw
* cell instance $30254 r0 *1 148.755,147.42
X$30254 488 623 489 644 645 cell_1rw
* cell instance $30255 m0 *1 148.755,152.88
X$30255 488 626 489 644 645 cell_1rw
* cell instance $30256 r0 *1 148.755,150.15
X$30256 488 625 489 644 645 cell_1rw
* cell instance $30257 m0 *1 148.755,155.61
X$30257 488 628 489 644 645 cell_1rw
* cell instance $30258 r0 *1 148.755,152.88
X$30258 488 627 489 644 645 cell_1rw
* cell instance $30259 r0 *1 148.755,155.61
X$30259 488 629 489 644 645 cell_1rw
* cell instance $30260 m0 *1 148.755,158.34
X$30260 488 630 489 644 645 cell_1rw
* cell instance $30261 r0 *1 148.755,158.34
X$30261 488 631 489 644 645 cell_1rw
* cell instance $30262 m0 *1 148.755,161.07
X$30262 488 632 489 644 645 cell_1rw
* cell instance $30263 r0 *1 148.755,161.07
X$30263 488 633 489 644 645 cell_1rw
* cell instance $30264 m0 *1 148.755,163.8
X$30264 488 634 489 644 645 cell_1rw
* cell instance $30265 r0 *1 148.755,163.8
X$30265 488 635 489 644 645 cell_1rw
* cell instance $30266 m0 *1 148.755,166.53
X$30266 488 637 489 644 645 cell_1rw
* cell instance $30267 m0 *1 148.755,169.26
X$30267 488 639 489 644 645 cell_1rw
* cell instance $30268 r0 *1 148.755,166.53
X$30268 488 636 489 644 645 cell_1rw
* cell instance $30269 r0 *1 148.755,169.26
X$30269 488 638 489 644 645 cell_1rw
* cell instance $30270 m0 *1 148.755,171.99
X$30270 488 640 489 644 645 cell_1rw
* cell instance $30271 r0 *1 148.755,171.99
X$30271 488 641 489 644 645 cell_1rw
* cell instance $30272 m0 *1 148.755,174.72
X$30272 488 642 489 644 645 cell_1rw
* cell instance $30273 r0 *1 148.755,174.72
X$30273 488 643 489 644 645 cell_1rw
* cell instance $30274 m0 *1 149.46,90.09
X$30274 490 581 491 644 645 cell_1rw
* cell instance $30275 m0 *1 149.46,92.82
X$30275 490 583 491 644 645 cell_1rw
* cell instance $30276 r0 *1 149.46,90.09
X$30276 490 580 491 644 645 cell_1rw
* cell instance $30277 m0 *1 149.46,95.55
X$30277 490 584 491 644 645 cell_1rw
* cell instance $30278 r0 *1 149.46,92.82
X$30278 490 582 491 644 645 cell_1rw
* cell instance $30279 r0 *1 149.46,95.55
X$30279 490 585 491 644 645 cell_1rw
* cell instance $30280 m0 *1 149.46,98.28
X$30280 490 586 491 644 645 cell_1rw
* cell instance $30281 r0 *1 149.46,98.28
X$30281 490 587 491 644 645 cell_1rw
* cell instance $30282 m0 *1 149.46,101.01
X$30282 490 588 491 644 645 cell_1rw
* cell instance $30283 r0 *1 149.46,101.01
X$30283 490 589 491 644 645 cell_1rw
* cell instance $30284 m0 *1 149.46,103.74
X$30284 490 590 491 644 645 cell_1rw
* cell instance $30285 r0 *1 149.46,103.74
X$30285 490 591 491 644 645 cell_1rw
* cell instance $30286 m0 *1 149.46,106.47
X$30286 490 593 491 644 645 cell_1rw
* cell instance $30287 r0 *1 149.46,106.47
X$30287 490 592 491 644 645 cell_1rw
* cell instance $30288 m0 *1 149.46,109.2
X$30288 490 594 491 644 645 cell_1rw
* cell instance $30289 r0 *1 149.46,109.2
X$30289 490 595 491 644 645 cell_1rw
* cell instance $30290 m0 *1 149.46,111.93
X$30290 490 597 491 644 645 cell_1rw
* cell instance $30291 m0 *1 149.46,114.66
X$30291 490 598 491 644 645 cell_1rw
* cell instance $30292 r0 *1 149.46,111.93
X$30292 490 596 491 644 645 cell_1rw
* cell instance $30293 r0 *1 149.46,114.66
X$30293 490 599 491 644 645 cell_1rw
* cell instance $30294 m0 *1 149.46,117.39
X$30294 490 600 491 644 645 cell_1rw
* cell instance $30295 m0 *1 149.46,120.12
X$30295 490 602 491 644 645 cell_1rw
* cell instance $30296 r0 *1 149.46,117.39
X$30296 490 601 491 644 645 cell_1rw
* cell instance $30297 r0 *1 149.46,120.12
X$30297 490 603 491 644 645 cell_1rw
* cell instance $30298 m0 *1 149.46,122.85
X$30298 490 604 491 644 645 cell_1rw
* cell instance $30299 r0 *1 149.46,122.85
X$30299 490 605 491 644 645 cell_1rw
* cell instance $30300 m0 *1 149.46,125.58
X$30300 490 606 491 644 645 cell_1rw
* cell instance $30301 r0 *1 149.46,125.58
X$30301 490 607 491 644 645 cell_1rw
* cell instance $30302 m0 *1 149.46,128.31
X$30302 490 609 491 644 645 cell_1rw
* cell instance $30303 r0 *1 149.46,128.31
X$30303 490 608 491 644 645 cell_1rw
* cell instance $30304 m0 *1 149.46,131.04
X$30304 490 610 491 644 645 cell_1rw
* cell instance $30305 r0 *1 149.46,131.04
X$30305 490 611 491 644 645 cell_1rw
* cell instance $30306 m0 *1 149.46,133.77
X$30306 490 612 491 644 645 cell_1rw
* cell instance $30307 r0 *1 149.46,133.77
X$30307 490 613 491 644 645 cell_1rw
* cell instance $30308 m0 *1 149.46,136.5
X$30308 490 615 491 644 645 cell_1rw
* cell instance $30309 r0 *1 149.46,136.5
X$30309 490 614 491 644 645 cell_1rw
* cell instance $30310 m0 *1 149.46,139.23
X$30310 490 617 491 644 645 cell_1rw
* cell instance $30311 m0 *1 149.46,141.96
X$30311 490 618 491 644 645 cell_1rw
* cell instance $30312 r0 *1 149.46,139.23
X$30312 490 616 491 644 645 cell_1rw
* cell instance $30313 m0 *1 149.46,144.69
X$30313 490 620 491 644 645 cell_1rw
* cell instance $30314 r0 *1 149.46,141.96
X$30314 490 619 491 644 645 cell_1rw
* cell instance $30315 r0 *1 149.46,144.69
X$30315 490 621 491 644 645 cell_1rw
* cell instance $30316 m0 *1 149.46,147.42
X$30316 490 622 491 644 645 cell_1rw
* cell instance $30317 r0 *1 149.46,147.42
X$30317 490 623 491 644 645 cell_1rw
* cell instance $30318 m0 *1 149.46,150.15
X$30318 490 624 491 644 645 cell_1rw
* cell instance $30319 m0 *1 149.46,152.88
X$30319 490 626 491 644 645 cell_1rw
* cell instance $30320 r0 *1 149.46,150.15
X$30320 490 625 491 644 645 cell_1rw
* cell instance $30321 r0 *1 149.46,152.88
X$30321 490 627 491 644 645 cell_1rw
* cell instance $30322 m0 *1 149.46,155.61
X$30322 490 628 491 644 645 cell_1rw
* cell instance $30323 r0 *1 149.46,155.61
X$30323 490 629 491 644 645 cell_1rw
* cell instance $30324 m0 *1 149.46,158.34
X$30324 490 630 491 644 645 cell_1rw
* cell instance $30325 r0 *1 149.46,158.34
X$30325 490 631 491 644 645 cell_1rw
* cell instance $30326 m0 *1 149.46,161.07
X$30326 490 632 491 644 645 cell_1rw
* cell instance $30327 r0 *1 149.46,161.07
X$30327 490 633 491 644 645 cell_1rw
* cell instance $30328 m0 *1 149.46,163.8
X$30328 490 634 491 644 645 cell_1rw
* cell instance $30329 m0 *1 149.46,166.53
X$30329 490 637 491 644 645 cell_1rw
* cell instance $30330 r0 *1 149.46,163.8
X$30330 490 635 491 644 645 cell_1rw
* cell instance $30331 r0 *1 149.46,166.53
X$30331 490 636 491 644 645 cell_1rw
* cell instance $30332 m0 *1 149.46,169.26
X$30332 490 639 491 644 645 cell_1rw
* cell instance $30333 r0 *1 149.46,169.26
X$30333 490 638 491 644 645 cell_1rw
* cell instance $30334 m0 *1 149.46,171.99
X$30334 490 640 491 644 645 cell_1rw
* cell instance $30335 r0 *1 149.46,171.99
X$30335 490 641 491 644 645 cell_1rw
* cell instance $30336 m0 *1 149.46,174.72
X$30336 490 642 491 644 645 cell_1rw
* cell instance $30337 r0 *1 149.46,174.72
X$30337 490 643 491 644 645 cell_1rw
* cell instance $30338 m0 *1 150.165,90.09
X$30338 492 581 493 644 645 cell_1rw
* cell instance $30339 r0 *1 150.165,90.09
X$30339 492 580 493 644 645 cell_1rw
* cell instance $30340 m0 *1 150.165,92.82
X$30340 492 583 493 644 645 cell_1rw
* cell instance $30341 r0 *1 150.165,92.82
X$30341 492 582 493 644 645 cell_1rw
* cell instance $30342 m0 *1 150.165,95.55
X$30342 492 584 493 644 645 cell_1rw
* cell instance $30343 r0 *1 150.165,95.55
X$30343 492 585 493 644 645 cell_1rw
* cell instance $30344 m0 *1 150.165,98.28
X$30344 492 586 493 644 645 cell_1rw
* cell instance $30345 r0 *1 150.165,98.28
X$30345 492 587 493 644 645 cell_1rw
* cell instance $30346 m0 *1 150.165,101.01
X$30346 492 588 493 644 645 cell_1rw
* cell instance $30347 r0 *1 150.165,101.01
X$30347 492 589 493 644 645 cell_1rw
* cell instance $30348 m0 *1 150.165,103.74
X$30348 492 590 493 644 645 cell_1rw
* cell instance $30349 m0 *1 150.165,106.47
X$30349 492 593 493 644 645 cell_1rw
* cell instance $30350 r0 *1 150.165,103.74
X$30350 492 591 493 644 645 cell_1rw
* cell instance $30351 r0 *1 150.165,106.47
X$30351 492 592 493 644 645 cell_1rw
* cell instance $30352 m0 *1 150.165,109.2
X$30352 492 594 493 644 645 cell_1rw
* cell instance $30353 r0 *1 150.165,109.2
X$30353 492 595 493 644 645 cell_1rw
* cell instance $30354 m0 *1 150.165,111.93
X$30354 492 597 493 644 645 cell_1rw
* cell instance $30355 r0 *1 150.165,111.93
X$30355 492 596 493 644 645 cell_1rw
* cell instance $30356 m0 *1 150.165,114.66
X$30356 492 598 493 644 645 cell_1rw
* cell instance $30357 r0 *1 150.165,114.66
X$30357 492 599 493 644 645 cell_1rw
* cell instance $30358 m0 *1 150.165,117.39
X$30358 492 600 493 644 645 cell_1rw
* cell instance $30359 r0 *1 150.165,117.39
X$30359 492 601 493 644 645 cell_1rw
* cell instance $30360 m0 *1 150.165,120.12
X$30360 492 602 493 644 645 cell_1rw
* cell instance $30361 r0 *1 150.165,120.12
X$30361 492 603 493 644 645 cell_1rw
* cell instance $30362 m0 *1 150.165,122.85
X$30362 492 604 493 644 645 cell_1rw
* cell instance $30363 r0 *1 150.165,122.85
X$30363 492 605 493 644 645 cell_1rw
* cell instance $30364 m0 *1 150.165,125.58
X$30364 492 606 493 644 645 cell_1rw
* cell instance $30365 r0 *1 150.165,125.58
X$30365 492 607 493 644 645 cell_1rw
* cell instance $30366 m0 *1 150.165,128.31
X$30366 492 609 493 644 645 cell_1rw
* cell instance $30367 r0 *1 150.165,128.31
X$30367 492 608 493 644 645 cell_1rw
* cell instance $30368 m0 *1 150.165,131.04
X$30368 492 610 493 644 645 cell_1rw
* cell instance $30369 r0 *1 150.165,131.04
X$30369 492 611 493 644 645 cell_1rw
* cell instance $30370 m0 *1 150.165,133.77
X$30370 492 612 493 644 645 cell_1rw
* cell instance $30371 r0 *1 150.165,133.77
X$30371 492 613 493 644 645 cell_1rw
* cell instance $30372 m0 *1 150.165,136.5
X$30372 492 615 493 644 645 cell_1rw
* cell instance $30373 r0 *1 150.165,136.5
X$30373 492 614 493 644 645 cell_1rw
* cell instance $30374 m0 *1 150.165,139.23
X$30374 492 617 493 644 645 cell_1rw
* cell instance $30375 r0 *1 150.165,139.23
X$30375 492 616 493 644 645 cell_1rw
* cell instance $30376 m0 *1 150.165,141.96
X$30376 492 618 493 644 645 cell_1rw
* cell instance $30377 r0 *1 150.165,141.96
X$30377 492 619 493 644 645 cell_1rw
* cell instance $30378 m0 *1 150.165,144.69
X$30378 492 620 493 644 645 cell_1rw
* cell instance $30379 r0 *1 150.165,144.69
X$30379 492 621 493 644 645 cell_1rw
* cell instance $30380 m0 *1 150.165,147.42
X$30380 492 622 493 644 645 cell_1rw
* cell instance $30381 r0 *1 150.165,147.42
X$30381 492 623 493 644 645 cell_1rw
* cell instance $30382 m0 *1 150.165,150.15
X$30382 492 624 493 644 645 cell_1rw
* cell instance $30383 m0 *1 150.165,152.88
X$30383 492 626 493 644 645 cell_1rw
* cell instance $30384 r0 *1 150.165,150.15
X$30384 492 625 493 644 645 cell_1rw
* cell instance $30385 r0 *1 150.165,152.88
X$30385 492 627 493 644 645 cell_1rw
* cell instance $30386 m0 *1 150.165,155.61
X$30386 492 628 493 644 645 cell_1rw
* cell instance $30387 r0 *1 150.165,155.61
X$30387 492 629 493 644 645 cell_1rw
* cell instance $30388 m0 *1 150.165,158.34
X$30388 492 630 493 644 645 cell_1rw
* cell instance $30389 r0 *1 150.165,158.34
X$30389 492 631 493 644 645 cell_1rw
* cell instance $30390 m0 *1 150.165,161.07
X$30390 492 632 493 644 645 cell_1rw
* cell instance $30391 r0 *1 150.165,161.07
X$30391 492 633 493 644 645 cell_1rw
* cell instance $30392 m0 *1 150.165,163.8
X$30392 492 634 493 644 645 cell_1rw
* cell instance $30393 r0 *1 150.165,163.8
X$30393 492 635 493 644 645 cell_1rw
* cell instance $30394 m0 *1 150.165,166.53
X$30394 492 637 493 644 645 cell_1rw
* cell instance $30395 r0 *1 150.165,166.53
X$30395 492 636 493 644 645 cell_1rw
* cell instance $30396 m0 *1 150.165,169.26
X$30396 492 639 493 644 645 cell_1rw
* cell instance $30397 r0 *1 150.165,169.26
X$30397 492 638 493 644 645 cell_1rw
* cell instance $30398 m0 *1 150.165,171.99
X$30398 492 640 493 644 645 cell_1rw
* cell instance $30399 r0 *1 150.165,171.99
X$30399 492 641 493 644 645 cell_1rw
* cell instance $30400 m0 *1 150.165,174.72
X$30400 492 642 493 644 645 cell_1rw
* cell instance $30401 r0 *1 150.165,174.72
X$30401 492 643 493 644 645 cell_1rw
* cell instance $30402 m0 *1 150.87,90.09
X$30402 494 581 495 644 645 cell_1rw
* cell instance $30403 r0 *1 150.87,90.09
X$30403 494 580 495 644 645 cell_1rw
* cell instance $30404 m0 *1 150.87,92.82
X$30404 494 583 495 644 645 cell_1rw
* cell instance $30405 m0 *1 150.87,95.55
X$30405 494 584 495 644 645 cell_1rw
* cell instance $30406 r0 *1 150.87,92.82
X$30406 494 582 495 644 645 cell_1rw
* cell instance $30407 r0 *1 150.87,95.55
X$30407 494 585 495 644 645 cell_1rw
* cell instance $30408 m0 *1 150.87,98.28
X$30408 494 586 495 644 645 cell_1rw
* cell instance $30409 r0 *1 150.87,98.28
X$30409 494 587 495 644 645 cell_1rw
* cell instance $30410 m0 *1 150.87,101.01
X$30410 494 588 495 644 645 cell_1rw
* cell instance $30411 r0 *1 150.87,101.01
X$30411 494 589 495 644 645 cell_1rw
* cell instance $30412 m0 *1 150.87,103.74
X$30412 494 590 495 644 645 cell_1rw
* cell instance $30413 r0 *1 150.87,103.74
X$30413 494 591 495 644 645 cell_1rw
* cell instance $30414 m0 *1 150.87,106.47
X$30414 494 593 495 644 645 cell_1rw
* cell instance $30415 r0 *1 150.87,106.47
X$30415 494 592 495 644 645 cell_1rw
* cell instance $30416 m0 *1 150.87,109.2
X$30416 494 594 495 644 645 cell_1rw
* cell instance $30417 r0 *1 150.87,109.2
X$30417 494 595 495 644 645 cell_1rw
* cell instance $30418 m0 *1 150.87,111.93
X$30418 494 597 495 644 645 cell_1rw
* cell instance $30419 m0 *1 150.87,114.66
X$30419 494 598 495 644 645 cell_1rw
* cell instance $30420 r0 *1 150.87,111.93
X$30420 494 596 495 644 645 cell_1rw
* cell instance $30421 r0 *1 150.87,114.66
X$30421 494 599 495 644 645 cell_1rw
* cell instance $30422 m0 *1 150.87,117.39
X$30422 494 600 495 644 645 cell_1rw
* cell instance $30423 r0 *1 150.87,117.39
X$30423 494 601 495 644 645 cell_1rw
* cell instance $30424 m0 *1 150.87,120.12
X$30424 494 602 495 644 645 cell_1rw
* cell instance $30425 r0 *1 150.87,120.12
X$30425 494 603 495 644 645 cell_1rw
* cell instance $30426 m0 *1 150.87,122.85
X$30426 494 604 495 644 645 cell_1rw
* cell instance $30427 r0 *1 150.87,122.85
X$30427 494 605 495 644 645 cell_1rw
* cell instance $30428 m0 *1 150.87,125.58
X$30428 494 606 495 644 645 cell_1rw
* cell instance $30429 r0 *1 150.87,125.58
X$30429 494 607 495 644 645 cell_1rw
* cell instance $30430 m0 *1 150.87,128.31
X$30430 494 609 495 644 645 cell_1rw
* cell instance $30431 m0 *1 150.87,131.04
X$30431 494 610 495 644 645 cell_1rw
* cell instance $30432 r0 *1 150.87,128.31
X$30432 494 608 495 644 645 cell_1rw
* cell instance $30433 m0 *1 150.87,133.77
X$30433 494 612 495 644 645 cell_1rw
* cell instance $30434 r0 *1 150.87,131.04
X$30434 494 611 495 644 645 cell_1rw
* cell instance $30435 r0 *1 150.87,133.77
X$30435 494 613 495 644 645 cell_1rw
* cell instance $30436 m0 *1 150.87,136.5
X$30436 494 615 495 644 645 cell_1rw
* cell instance $30437 r0 *1 150.87,136.5
X$30437 494 614 495 644 645 cell_1rw
* cell instance $30438 m0 *1 150.87,139.23
X$30438 494 617 495 644 645 cell_1rw
* cell instance $30439 r0 *1 150.87,139.23
X$30439 494 616 495 644 645 cell_1rw
* cell instance $30440 m0 *1 150.87,141.96
X$30440 494 618 495 644 645 cell_1rw
* cell instance $30441 r0 *1 150.87,141.96
X$30441 494 619 495 644 645 cell_1rw
* cell instance $30442 m0 *1 150.87,144.69
X$30442 494 620 495 644 645 cell_1rw
* cell instance $30443 r0 *1 150.87,144.69
X$30443 494 621 495 644 645 cell_1rw
* cell instance $30444 m0 *1 150.87,147.42
X$30444 494 622 495 644 645 cell_1rw
* cell instance $30445 m0 *1 150.87,150.15
X$30445 494 624 495 644 645 cell_1rw
* cell instance $30446 r0 *1 150.87,147.42
X$30446 494 623 495 644 645 cell_1rw
* cell instance $30447 r0 *1 150.87,150.15
X$30447 494 625 495 644 645 cell_1rw
* cell instance $30448 m0 *1 150.87,152.88
X$30448 494 626 495 644 645 cell_1rw
* cell instance $30449 r0 *1 150.87,152.88
X$30449 494 627 495 644 645 cell_1rw
* cell instance $30450 m0 *1 150.87,155.61
X$30450 494 628 495 644 645 cell_1rw
* cell instance $30451 r0 *1 150.87,155.61
X$30451 494 629 495 644 645 cell_1rw
* cell instance $30452 m0 *1 150.87,158.34
X$30452 494 630 495 644 645 cell_1rw
* cell instance $30453 r0 *1 150.87,158.34
X$30453 494 631 495 644 645 cell_1rw
* cell instance $30454 m0 *1 150.87,161.07
X$30454 494 632 495 644 645 cell_1rw
* cell instance $30455 r0 *1 150.87,161.07
X$30455 494 633 495 644 645 cell_1rw
* cell instance $30456 m0 *1 150.87,163.8
X$30456 494 634 495 644 645 cell_1rw
* cell instance $30457 r0 *1 150.87,163.8
X$30457 494 635 495 644 645 cell_1rw
* cell instance $30458 m0 *1 150.87,166.53
X$30458 494 637 495 644 645 cell_1rw
* cell instance $30459 r0 *1 150.87,166.53
X$30459 494 636 495 644 645 cell_1rw
* cell instance $30460 m0 *1 150.87,169.26
X$30460 494 639 495 644 645 cell_1rw
* cell instance $30461 m0 *1 150.87,171.99
X$30461 494 640 495 644 645 cell_1rw
* cell instance $30462 r0 *1 150.87,169.26
X$30462 494 638 495 644 645 cell_1rw
* cell instance $30463 r0 *1 150.87,171.99
X$30463 494 641 495 644 645 cell_1rw
* cell instance $30464 m0 *1 150.87,174.72
X$30464 494 642 495 644 645 cell_1rw
* cell instance $30465 r0 *1 150.87,174.72
X$30465 494 643 495 644 645 cell_1rw
* cell instance $30466 m0 *1 151.575,90.09
X$30466 496 581 497 644 645 cell_1rw
* cell instance $30467 r0 *1 151.575,90.09
X$30467 496 580 497 644 645 cell_1rw
* cell instance $30468 m0 *1 151.575,92.82
X$30468 496 583 497 644 645 cell_1rw
* cell instance $30469 r0 *1 151.575,92.82
X$30469 496 582 497 644 645 cell_1rw
* cell instance $30470 m0 *1 151.575,95.55
X$30470 496 584 497 644 645 cell_1rw
* cell instance $30471 r0 *1 151.575,95.55
X$30471 496 585 497 644 645 cell_1rw
* cell instance $30472 m0 *1 151.575,98.28
X$30472 496 586 497 644 645 cell_1rw
* cell instance $30473 r0 *1 151.575,98.28
X$30473 496 587 497 644 645 cell_1rw
* cell instance $30474 m0 *1 151.575,101.01
X$30474 496 588 497 644 645 cell_1rw
* cell instance $30475 r0 *1 151.575,101.01
X$30475 496 589 497 644 645 cell_1rw
* cell instance $30476 m0 *1 151.575,103.74
X$30476 496 590 497 644 645 cell_1rw
* cell instance $30477 r0 *1 151.575,103.74
X$30477 496 591 497 644 645 cell_1rw
* cell instance $30478 m0 *1 151.575,106.47
X$30478 496 593 497 644 645 cell_1rw
* cell instance $30479 r0 *1 151.575,106.47
X$30479 496 592 497 644 645 cell_1rw
* cell instance $30480 m0 *1 151.575,109.2
X$30480 496 594 497 644 645 cell_1rw
* cell instance $30481 r0 *1 151.575,109.2
X$30481 496 595 497 644 645 cell_1rw
* cell instance $30482 m0 *1 151.575,111.93
X$30482 496 597 497 644 645 cell_1rw
* cell instance $30483 r0 *1 151.575,111.93
X$30483 496 596 497 644 645 cell_1rw
* cell instance $30484 m0 *1 151.575,114.66
X$30484 496 598 497 644 645 cell_1rw
* cell instance $30485 r0 *1 151.575,114.66
X$30485 496 599 497 644 645 cell_1rw
* cell instance $30486 m0 *1 151.575,117.39
X$30486 496 600 497 644 645 cell_1rw
* cell instance $30487 r0 *1 151.575,117.39
X$30487 496 601 497 644 645 cell_1rw
* cell instance $30488 m0 *1 151.575,120.12
X$30488 496 602 497 644 645 cell_1rw
* cell instance $30489 r0 *1 151.575,120.12
X$30489 496 603 497 644 645 cell_1rw
* cell instance $30490 m0 *1 151.575,122.85
X$30490 496 604 497 644 645 cell_1rw
* cell instance $30491 m0 *1 151.575,125.58
X$30491 496 606 497 644 645 cell_1rw
* cell instance $30492 r0 *1 151.575,122.85
X$30492 496 605 497 644 645 cell_1rw
* cell instance $30493 r0 *1 151.575,125.58
X$30493 496 607 497 644 645 cell_1rw
* cell instance $30494 m0 *1 151.575,128.31
X$30494 496 609 497 644 645 cell_1rw
* cell instance $30495 r0 *1 151.575,128.31
X$30495 496 608 497 644 645 cell_1rw
* cell instance $30496 m0 *1 151.575,131.04
X$30496 496 610 497 644 645 cell_1rw
* cell instance $30497 r0 *1 151.575,131.04
X$30497 496 611 497 644 645 cell_1rw
* cell instance $30498 m0 *1 151.575,133.77
X$30498 496 612 497 644 645 cell_1rw
* cell instance $30499 m0 *1 151.575,136.5
X$30499 496 615 497 644 645 cell_1rw
* cell instance $30500 r0 *1 151.575,133.77
X$30500 496 613 497 644 645 cell_1rw
* cell instance $30501 r0 *1 151.575,136.5
X$30501 496 614 497 644 645 cell_1rw
* cell instance $30502 m0 *1 151.575,139.23
X$30502 496 617 497 644 645 cell_1rw
* cell instance $30503 r0 *1 151.575,139.23
X$30503 496 616 497 644 645 cell_1rw
* cell instance $30504 m0 *1 151.575,141.96
X$30504 496 618 497 644 645 cell_1rw
* cell instance $30505 m0 *1 151.575,144.69
X$30505 496 620 497 644 645 cell_1rw
* cell instance $30506 r0 *1 151.575,141.96
X$30506 496 619 497 644 645 cell_1rw
* cell instance $30507 m0 *1 151.575,147.42
X$30507 496 622 497 644 645 cell_1rw
* cell instance $30508 r0 *1 151.575,144.69
X$30508 496 621 497 644 645 cell_1rw
* cell instance $30509 r0 *1 151.575,147.42
X$30509 496 623 497 644 645 cell_1rw
* cell instance $30510 m0 *1 151.575,150.15
X$30510 496 624 497 644 645 cell_1rw
* cell instance $30511 r0 *1 151.575,150.15
X$30511 496 625 497 644 645 cell_1rw
* cell instance $30512 m0 *1 151.575,152.88
X$30512 496 626 497 644 645 cell_1rw
* cell instance $30513 r0 *1 151.575,152.88
X$30513 496 627 497 644 645 cell_1rw
* cell instance $30514 m0 *1 151.575,155.61
X$30514 496 628 497 644 645 cell_1rw
* cell instance $30515 m0 *1 151.575,158.34
X$30515 496 630 497 644 645 cell_1rw
* cell instance $30516 r0 *1 151.575,155.61
X$30516 496 629 497 644 645 cell_1rw
* cell instance $30517 r0 *1 151.575,158.34
X$30517 496 631 497 644 645 cell_1rw
* cell instance $30518 m0 *1 151.575,161.07
X$30518 496 632 497 644 645 cell_1rw
* cell instance $30519 r0 *1 151.575,161.07
X$30519 496 633 497 644 645 cell_1rw
* cell instance $30520 m0 *1 151.575,163.8
X$30520 496 634 497 644 645 cell_1rw
* cell instance $30521 r0 *1 151.575,163.8
X$30521 496 635 497 644 645 cell_1rw
* cell instance $30522 m0 *1 151.575,166.53
X$30522 496 637 497 644 645 cell_1rw
* cell instance $30523 r0 *1 151.575,166.53
X$30523 496 636 497 644 645 cell_1rw
* cell instance $30524 m0 *1 151.575,169.26
X$30524 496 639 497 644 645 cell_1rw
* cell instance $30525 r0 *1 151.575,169.26
X$30525 496 638 497 644 645 cell_1rw
* cell instance $30526 m0 *1 151.575,171.99
X$30526 496 640 497 644 645 cell_1rw
* cell instance $30527 m0 *1 151.575,174.72
X$30527 496 642 497 644 645 cell_1rw
* cell instance $30528 r0 *1 151.575,171.99
X$30528 496 641 497 644 645 cell_1rw
* cell instance $30529 r0 *1 151.575,174.72
X$30529 496 643 497 644 645 cell_1rw
* cell instance $30530 m0 *1 152.28,90.09
X$30530 498 581 499 644 645 cell_1rw
* cell instance $30531 r0 *1 152.28,90.09
X$30531 498 580 499 644 645 cell_1rw
* cell instance $30532 m0 *1 152.28,92.82
X$30532 498 583 499 644 645 cell_1rw
* cell instance $30533 r0 *1 152.28,92.82
X$30533 498 582 499 644 645 cell_1rw
* cell instance $30534 m0 *1 152.28,95.55
X$30534 498 584 499 644 645 cell_1rw
* cell instance $30535 r0 *1 152.28,95.55
X$30535 498 585 499 644 645 cell_1rw
* cell instance $30536 m0 *1 152.28,98.28
X$30536 498 586 499 644 645 cell_1rw
* cell instance $30537 m0 *1 152.28,101.01
X$30537 498 588 499 644 645 cell_1rw
* cell instance $30538 r0 *1 152.28,98.28
X$30538 498 587 499 644 645 cell_1rw
* cell instance $30539 r0 *1 152.28,101.01
X$30539 498 589 499 644 645 cell_1rw
* cell instance $30540 m0 *1 152.28,103.74
X$30540 498 590 499 644 645 cell_1rw
* cell instance $30541 r0 *1 152.28,103.74
X$30541 498 591 499 644 645 cell_1rw
* cell instance $30542 m0 *1 152.28,106.47
X$30542 498 593 499 644 645 cell_1rw
* cell instance $30543 r0 *1 152.28,106.47
X$30543 498 592 499 644 645 cell_1rw
* cell instance $30544 m0 *1 152.28,109.2
X$30544 498 594 499 644 645 cell_1rw
* cell instance $30545 r0 *1 152.28,109.2
X$30545 498 595 499 644 645 cell_1rw
* cell instance $30546 m0 *1 152.28,111.93
X$30546 498 597 499 644 645 cell_1rw
* cell instance $30547 m0 *1 152.28,114.66
X$30547 498 598 499 644 645 cell_1rw
* cell instance $30548 r0 *1 152.28,111.93
X$30548 498 596 499 644 645 cell_1rw
* cell instance $30549 r0 *1 152.28,114.66
X$30549 498 599 499 644 645 cell_1rw
* cell instance $30550 m0 *1 152.28,117.39
X$30550 498 600 499 644 645 cell_1rw
* cell instance $30551 r0 *1 152.28,117.39
X$30551 498 601 499 644 645 cell_1rw
* cell instance $30552 m0 *1 152.28,120.12
X$30552 498 602 499 644 645 cell_1rw
* cell instance $30553 r0 *1 152.28,120.12
X$30553 498 603 499 644 645 cell_1rw
* cell instance $30554 m0 *1 152.28,122.85
X$30554 498 604 499 644 645 cell_1rw
* cell instance $30555 r0 *1 152.28,122.85
X$30555 498 605 499 644 645 cell_1rw
* cell instance $30556 m0 *1 152.28,125.58
X$30556 498 606 499 644 645 cell_1rw
* cell instance $30557 m0 *1 152.28,128.31
X$30557 498 609 499 644 645 cell_1rw
* cell instance $30558 r0 *1 152.28,125.58
X$30558 498 607 499 644 645 cell_1rw
* cell instance $30559 r0 *1 152.28,128.31
X$30559 498 608 499 644 645 cell_1rw
* cell instance $30560 m0 *1 152.28,131.04
X$30560 498 610 499 644 645 cell_1rw
* cell instance $30561 r0 *1 152.28,131.04
X$30561 498 611 499 644 645 cell_1rw
* cell instance $30562 m0 *1 152.28,133.77
X$30562 498 612 499 644 645 cell_1rw
* cell instance $30563 r0 *1 152.28,133.77
X$30563 498 613 499 644 645 cell_1rw
* cell instance $30564 m0 *1 152.28,136.5
X$30564 498 615 499 644 645 cell_1rw
* cell instance $30565 r0 *1 152.28,136.5
X$30565 498 614 499 644 645 cell_1rw
* cell instance $30566 m0 *1 152.28,139.23
X$30566 498 617 499 644 645 cell_1rw
* cell instance $30567 r0 *1 152.28,139.23
X$30567 498 616 499 644 645 cell_1rw
* cell instance $30568 m0 *1 152.28,141.96
X$30568 498 618 499 644 645 cell_1rw
* cell instance $30569 r0 *1 152.28,141.96
X$30569 498 619 499 644 645 cell_1rw
* cell instance $30570 m0 *1 152.28,144.69
X$30570 498 620 499 644 645 cell_1rw
* cell instance $30571 r0 *1 152.28,144.69
X$30571 498 621 499 644 645 cell_1rw
* cell instance $30572 m0 *1 152.28,147.42
X$30572 498 622 499 644 645 cell_1rw
* cell instance $30573 r0 *1 152.28,147.42
X$30573 498 623 499 644 645 cell_1rw
* cell instance $30574 m0 *1 152.28,150.15
X$30574 498 624 499 644 645 cell_1rw
* cell instance $30575 r0 *1 152.28,150.15
X$30575 498 625 499 644 645 cell_1rw
* cell instance $30576 m0 *1 152.28,152.88
X$30576 498 626 499 644 645 cell_1rw
* cell instance $30577 r0 *1 152.28,152.88
X$30577 498 627 499 644 645 cell_1rw
* cell instance $30578 m0 *1 152.28,155.61
X$30578 498 628 499 644 645 cell_1rw
* cell instance $30579 r0 *1 152.28,155.61
X$30579 498 629 499 644 645 cell_1rw
* cell instance $30580 m0 *1 152.28,158.34
X$30580 498 630 499 644 645 cell_1rw
* cell instance $30581 r0 *1 152.28,158.34
X$30581 498 631 499 644 645 cell_1rw
* cell instance $30582 m0 *1 152.28,161.07
X$30582 498 632 499 644 645 cell_1rw
* cell instance $30583 r0 *1 152.28,161.07
X$30583 498 633 499 644 645 cell_1rw
* cell instance $30584 m0 *1 152.28,163.8
X$30584 498 634 499 644 645 cell_1rw
* cell instance $30585 r0 *1 152.28,163.8
X$30585 498 635 499 644 645 cell_1rw
* cell instance $30586 m0 *1 152.28,166.53
X$30586 498 637 499 644 645 cell_1rw
* cell instance $30587 r0 *1 152.28,166.53
X$30587 498 636 499 644 645 cell_1rw
* cell instance $30588 m0 *1 152.28,169.26
X$30588 498 639 499 644 645 cell_1rw
* cell instance $30589 m0 *1 152.28,171.99
X$30589 498 640 499 644 645 cell_1rw
* cell instance $30590 r0 *1 152.28,169.26
X$30590 498 638 499 644 645 cell_1rw
* cell instance $30591 m0 *1 152.28,174.72
X$30591 498 642 499 644 645 cell_1rw
* cell instance $30592 r0 *1 152.28,171.99
X$30592 498 641 499 644 645 cell_1rw
* cell instance $30593 r0 *1 152.28,174.72
X$30593 498 643 499 644 645 cell_1rw
* cell instance $30594 m0 *1 152.985,90.09
X$30594 500 581 501 644 645 cell_1rw
* cell instance $30595 r0 *1 152.985,90.09
X$30595 500 580 501 644 645 cell_1rw
* cell instance $30596 m0 *1 152.985,92.82
X$30596 500 583 501 644 645 cell_1rw
* cell instance $30597 m0 *1 152.985,95.55
X$30597 500 584 501 644 645 cell_1rw
* cell instance $30598 r0 *1 152.985,92.82
X$30598 500 582 501 644 645 cell_1rw
* cell instance $30599 r0 *1 152.985,95.55
X$30599 500 585 501 644 645 cell_1rw
* cell instance $30600 m0 *1 152.985,98.28
X$30600 500 586 501 644 645 cell_1rw
* cell instance $30601 r0 *1 152.985,98.28
X$30601 500 587 501 644 645 cell_1rw
* cell instance $30602 m0 *1 152.985,101.01
X$30602 500 588 501 644 645 cell_1rw
* cell instance $30603 r0 *1 152.985,101.01
X$30603 500 589 501 644 645 cell_1rw
* cell instance $30604 m0 *1 152.985,103.74
X$30604 500 590 501 644 645 cell_1rw
* cell instance $30605 r0 *1 152.985,103.74
X$30605 500 591 501 644 645 cell_1rw
* cell instance $30606 m0 *1 152.985,106.47
X$30606 500 593 501 644 645 cell_1rw
* cell instance $30607 r0 *1 152.985,106.47
X$30607 500 592 501 644 645 cell_1rw
* cell instance $30608 m0 *1 152.985,109.2
X$30608 500 594 501 644 645 cell_1rw
* cell instance $30609 r0 *1 152.985,109.2
X$30609 500 595 501 644 645 cell_1rw
* cell instance $30610 m0 *1 152.985,111.93
X$30610 500 597 501 644 645 cell_1rw
* cell instance $30611 m0 *1 152.985,114.66
X$30611 500 598 501 644 645 cell_1rw
* cell instance $30612 r0 *1 152.985,111.93
X$30612 500 596 501 644 645 cell_1rw
* cell instance $30613 r0 *1 152.985,114.66
X$30613 500 599 501 644 645 cell_1rw
* cell instance $30614 m0 *1 152.985,117.39
X$30614 500 600 501 644 645 cell_1rw
* cell instance $30615 m0 *1 152.985,120.12
X$30615 500 602 501 644 645 cell_1rw
* cell instance $30616 r0 *1 152.985,117.39
X$30616 500 601 501 644 645 cell_1rw
* cell instance $30617 r0 *1 152.985,120.12
X$30617 500 603 501 644 645 cell_1rw
* cell instance $30618 m0 *1 152.985,122.85
X$30618 500 604 501 644 645 cell_1rw
* cell instance $30619 r0 *1 152.985,122.85
X$30619 500 605 501 644 645 cell_1rw
* cell instance $30620 m0 *1 152.985,125.58
X$30620 500 606 501 644 645 cell_1rw
* cell instance $30621 m0 *1 152.985,128.31
X$30621 500 609 501 644 645 cell_1rw
* cell instance $30622 r0 *1 152.985,125.58
X$30622 500 607 501 644 645 cell_1rw
* cell instance $30623 r0 *1 152.985,128.31
X$30623 500 608 501 644 645 cell_1rw
* cell instance $30624 m0 *1 152.985,131.04
X$30624 500 610 501 644 645 cell_1rw
* cell instance $30625 m0 *1 152.985,133.77
X$30625 500 612 501 644 645 cell_1rw
* cell instance $30626 r0 *1 152.985,131.04
X$30626 500 611 501 644 645 cell_1rw
* cell instance $30627 r0 *1 152.985,133.77
X$30627 500 613 501 644 645 cell_1rw
* cell instance $30628 m0 *1 152.985,136.5
X$30628 500 615 501 644 645 cell_1rw
* cell instance $30629 m0 *1 152.985,139.23
X$30629 500 617 501 644 645 cell_1rw
* cell instance $30630 r0 *1 152.985,136.5
X$30630 500 614 501 644 645 cell_1rw
* cell instance $30631 r0 *1 152.985,139.23
X$30631 500 616 501 644 645 cell_1rw
* cell instance $30632 m0 *1 152.985,141.96
X$30632 500 618 501 644 645 cell_1rw
* cell instance $30633 r0 *1 152.985,141.96
X$30633 500 619 501 644 645 cell_1rw
* cell instance $30634 m0 *1 152.985,144.69
X$30634 500 620 501 644 645 cell_1rw
* cell instance $30635 r0 *1 152.985,144.69
X$30635 500 621 501 644 645 cell_1rw
* cell instance $30636 m0 *1 152.985,147.42
X$30636 500 622 501 644 645 cell_1rw
* cell instance $30637 r0 *1 152.985,147.42
X$30637 500 623 501 644 645 cell_1rw
* cell instance $30638 m0 *1 152.985,150.15
X$30638 500 624 501 644 645 cell_1rw
* cell instance $30639 r0 *1 152.985,150.15
X$30639 500 625 501 644 645 cell_1rw
* cell instance $30640 m0 *1 152.985,152.88
X$30640 500 626 501 644 645 cell_1rw
* cell instance $30641 r0 *1 152.985,152.88
X$30641 500 627 501 644 645 cell_1rw
* cell instance $30642 m0 *1 152.985,155.61
X$30642 500 628 501 644 645 cell_1rw
* cell instance $30643 r0 *1 152.985,155.61
X$30643 500 629 501 644 645 cell_1rw
* cell instance $30644 m0 *1 152.985,158.34
X$30644 500 630 501 644 645 cell_1rw
* cell instance $30645 m0 *1 152.985,161.07
X$30645 500 632 501 644 645 cell_1rw
* cell instance $30646 r0 *1 152.985,158.34
X$30646 500 631 501 644 645 cell_1rw
* cell instance $30647 r0 *1 152.985,161.07
X$30647 500 633 501 644 645 cell_1rw
* cell instance $30648 m0 *1 152.985,163.8
X$30648 500 634 501 644 645 cell_1rw
* cell instance $30649 r0 *1 152.985,163.8
X$30649 500 635 501 644 645 cell_1rw
* cell instance $30650 m0 *1 152.985,166.53
X$30650 500 637 501 644 645 cell_1rw
* cell instance $30651 r0 *1 152.985,166.53
X$30651 500 636 501 644 645 cell_1rw
* cell instance $30652 m0 *1 152.985,169.26
X$30652 500 639 501 644 645 cell_1rw
* cell instance $30653 r0 *1 152.985,169.26
X$30653 500 638 501 644 645 cell_1rw
* cell instance $30654 m0 *1 152.985,171.99
X$30654 500 640 501 644 645 cell_1rw
* cell instance $30655 r0 *1 152.985,171.99
X$30655 500 641 501 644 645 cell_1rw
* cell instance $30656 m0 *1 152.985,174.72
X$30656 500 642 501 644 645 cell_1rw
* cell instance $30657 r0 *1 152.985,174.72
X$30657 500 643 501 644 645 cell_1rw
* cell instance $30658 m0 *1 153.69,90.09
X$30658 502 581 503 644 645 cell_1rw
* cell instance $30659 r0 *1 153.69,90.09
X$30659 502 580 503 644 645 cell_1rw
* cell instance $30660 m0 *1 153.69,92.82
X$30660 502 583 503 644 645 cell_1rw
* cell instance $30661 r0 *1 153.69,92.82
X$30661 502 582 503 644 645 cell_1rw
* cell instance $30662 m0 *1 153.69,95.55
X$30662 502 584 503 644 645 cell_1rw
* cell instance $30663 r0 *1 153.69,95.55
X$30663 502 585 503 644 645 cell_1rw
* cell instance $30664 m0 *1 153.69,98.28
X$30664 502 586 503 644 645 cell_1rw
* cell instance $30665 m0 *1 153.69,101.01
X$30665 502 588 503 644 645 cell_1rw
* cell instance $30666 r0 *1 153.69,98.28
X$30666 502 587 503 644 645 cell_1rw
* cell instance $30667 r0 *1 153.69,101.01
X$30667 502 589 503 644 645 cell_1rw
* cell instance $30668 m0 *1 153.69,103.74
X$30668 502 590 503 644 645 cell_1rw
* cell instance $30669 r0 *1 153.69,103.74
X$30669 502 591 503 644 645 cell_1rw
* cell instance $30670 m0 *1 153.69,106.47
X$30670 502 593 503 644 645 cell_1rw
* cell instance $30671 m0 *1 153.69,109.2
X$30671 502 594 503 644 645 cell_1rw
* cell instance $30672 r0 *1 153.69,106.47
X$30672 502 592 503 644 645 cell_1rw
* cell instance $30673 r0 *1 153.69,109.2
X$30673 502 595 503 644 645 cell_1rw
* cell instance $30674 m0 *1 153.69,111.93
X$30674 502 597 503 644 645 cell_1rw
* cell instance $30675 r0 *1 153.69,111.93
X$30675 502 596 503 644 645 cell_1rw
* cell instance $30676 m0 *1 153.69,114.66
X$30676 502 598 503 644 645 cell_1rw
* cell instance $30677 r0 *1 153.69,114.66
X$30677 502 599 503 644 645 cell_1rw
* cell instance $30678 m0 *1 153.69,117.39
X$30678 502 600 503 644 645 cell_1rw
* cell instance $30679 r0 *1 153.69,117.39
X$30679 502 601 503 644 645 cell_1rw
* cell instance $30680 m0 *1 153.69,120.12
X$30680 502 602 503 644 645 cell_1rw
* cell instance $30681 r0 *1 153.69,120.12
X$30681 502 603 503 644 645 cell_1rw
* cell instance $30682 m0 *1 153.69,122.85
X$30682 502 604 503 644 645 cell_1rw
* cell instance $30683 r0 *1 153.69,122.85
X$30683 502 605 503 644 645 cell_1rw
* cell instance $30684 m0 *1 153.69,125.58
X$30684 502 606 503 644 645 cell_1rw
* cell instance $30685 r0 *1 153.69,125.58
X$30685 502 607 503 644 645 cell_1rw
* cell instance $30686 m0 *1 153.69,128.31
X$30686 502 609 503 644 645 cell_1rw
* cell instance $30687 r0 *1 153.69,128.31
X$30687 502 608 503 644 645 cell_1rw
* cell instance $30688 m0 *1 153.69,131.04
X$30688 502 610 503 644 645 cell_1rw
* cell instance $30689 r0 *1 153.69,131.04
X$30689 502 611 503 644 645 cell_1rw
* cell instance $30690 m0 *1 153.69,133.77
X$30690 502 612 503 644 645 cell_1rw
* cell instance $30691 m0 *1 153.69,136.5
X$30691 502 615 503 644 645 cell_1rw
* cell instance $30692 r0 *1 153.69,133.77
X$30692 502 613 503 644 645 cell_1rw
* cell instance $30693 m0 *1 153.69,139.23
X$30693 502 617 503 644 645 cell_1rw
* cell instance $30694 r0 *1 153.69,136.5
X$30694 502 614 503 644 645 cell_1rw
* cell instance $30695 r0 *1 153.69,139.23
X$30695 502 616 503 644 645 cell_1rw
* cell instance $30696 m0 *1 153.69,141.96
X$30696 502 618 503 644 645 cell_1rw
* cell instance $30697 r0 *1 153.69,141.96
X$30697 502 619 503 644 645 cell_1rw
* cell instance $30698 m0 *1 153.69,144.69
X$30698 502 620 503 644 645 cell_1rw
* cell instance $30699 r0 *1 153.69,144.69
X$30699 502 621 503 644 645 cell_1rw
* cell instance $30700 m0 *1 153.69,147.42
X$30700 502 622 503 644 645 cell_1rw
* cell instance $30701 r0 *1 153.69,147.42
X$30701 502 623 503 644 645 cell_1rw
* cell instance $30702 m0 *1 153.69,150.15
X$30702 502 624 503 644 645 cell_1rw
* cell instance $30703 r0 *1 153.69,150.15
X$30703 502 625 503 644 645 cell_1rw
* cell instance $30704 m0 *1 153.69,152.88
X$30704 502 626 503 644 645 cell_1rw
* cell instance $30705 r0 *1 153.69,152.88
X$30705 502 627 503 644 645 cell_1rw
* cell instance $30706 m0 *1 153.69,155.61
X$30706 502 628 503 644 645 cell_1rw
* cell instance $30707 m0 *1 153.69,158.34
X$30707 502 630 503 644 645 cell_1rw
* cell instance $30708 r0 *1 153.69,155.61
X$30708 502 629 503 644 645 cell_1rw
* cell instance $30709 r0 *1 153.69,158.34
X$30709 502 631 503 644 645 cell_1rw
* cell instance $30710 m0 *1 153.69,161.07
X$30710 502 632 503 644 645 cell_1rw
* cell instance $30711 m0 *1 153.69,163.8
X$30711 502 634 503 644 645 cell_1rw
* cell instance $30712 r0 *1 153.69,161.07
X$30712 502 633 503 644 645 cell_1rw
* cell instance $30713 r0 *1 153.69,163.8
X$30713 502 635 503 644 645 cell_1rw
* cell instance $30714 m0 *1 153.69,166.53
X$30714 502 637 503 644 645 cell_1rw
* cell instance $30715 r0 *1 153.69,166.53
X$30715 502 636 503 644 645 cell_1rw
* cell instance $30716 m0 *1 153.69,169.26
X$30716 502 639 503 644 645 cell_1rw
* cell instance $30717 r0 *1 153.69,169.26
X$30717 502 638 503 644 645 cell_1rw
* cell instance $30718 m0 *1 153.69,171.99
X$30718 502 640 503 644 645 cell_1rw
* cell instance $30719 m0 *1 153.69,174.72
X$30719 502 642 503 644 645 cell_1rw
* cell instance $30720 r0 *1 153.69,171.99
X$30720 502 641 503 644 645 cell_1rw
* cell instance $30721 r0 *1 153.69,174.72
X$30721 502 643 503 644 645 cell_1rw
* cell instance $30722 m0 *1 154.395,90.09
X$30722 504 581 505 644 645 cell_1rw
* cell instance $30723 r0 *1 154.395,90.09
X$30723 504 580 505 644 645 cell_1rw
* cell instance $30724 m0 *1 154.395,92.82
X$30724 504 583 505 644 645 cell_1rw
* cell instance $30725 r0 *1 154.395,92.82
X$30725 504 582 505 644 645 cell_1rw
* cell instance $30726 m0 *1 154.395,95.55
X$30726 504 584 505 644 645 cell_1rw
* cell instance $30727 m0 *1 154.395,98.28
X$30727 504 586 505 644 645 cell_1rw
* cell instance $30728 r0 *1 154.395,95.55
X$30728 504 585 505 644 645 cell_1rw
* cell instance $30729 r0 *1 154.395,98.28
X$30729 504 587 505 644 645 cell_1rw
* cell instance $30730 m0 *1 154.395,101.01
X$30730 504 588 505 644 645 cell_1rw
* cell instance $30731 r0 *1 154.395,101.01
X$30731 504 589 505 644 645 cell_1rw
* cell instance $30732 m0 *1 154.395,103.74
X$30732 504 590 505 644 645 cell_1rw
* cell instance $30733 m0 *1 154.395,106.47
X$30733 504 593 505 644 645 cell_1rw
* cell instance $30734 r0 *1 154.395,103.74
X$30734 504 591 505 644 645 cell_1rw
* cell instance $30735 r0 *1 154.395,106.47
X$30735 504 592 505 644 645 cell_1rw
* cell instance $30736 m0 *1 154.395,109.2
X$30736 504 594 505 644 645 cell_1rw
* cell instance $30737 r0 *1 154.395,109.2
X$30737 504 595 505 644 645 cell_1rw
* cell instance $30738 m0 *1 154.395,111.93
X$30738 504 597 505 644 645 cell_1rw
* cell instance $30739 r0 *1 154.395,111.93
X$30739 504 596 505 644 645 cell_1rw
* cell instance $30740 m0 *1 154.395,114.66
X$30740 504 598 505 644 645 cell_1rw
* cell instance $30741 m0 *1 154.395,117.39
X$30741 504 600 505 644 645 cell_1rw
* cell instance $30742 r0 *1 154.395,114.66
X$30742 504 599 505 644 645 cell_1rw
* cell instance $30743 r0 *1 154.395,117.39
X$30743 504 601 505 644 645 cell_1rw
* cell instance $30744 m0 *1 154.395,120.12
X$30744 504 602 505 644 645 cell_1rw
* cell instance $30745 r0 *1 154.395,120.12
X$30745 504 603 505 644 645 cell_1rw
* cell instance $30746 m0 *1 154.395,122.85
X$30746 504 604 505 644 645 cell_1rw
* cell instance $30747 r0 *1 154.395,122.85
X$30747 504 605 505 644 645 cell_1rw
* cell instance $30748 m0 *1 154.395,125.58
X$30748 504 606 505 644 645 cell_1rw
* cell instance $30749 m0 *1 154.395,128.31
X$30749 504 609 505 644 645 cell_1rw
* cell instance $30750 r0 *1 154.395,125.58
X$30750 504 607 505 644 645 cell_1rw
* cell instance $30751 r0 *1 154.395,128.31
X$30751 504 608 505 644 645 cell_1rw
* cell instance $30752 m0 *1 154.395,131.04
X$30752 504 610 505 644 645 cell_1rw
* cell instance $30753 r0 *1 154.395,131.04
X$30753 504 611 505 644 645 cell_1rw
* cell instance $30754 m0 *1 154.395,133.77
X$30754 504 612 505 644 645 cell_1rw
* cell instance $30755 r0 *1 154.395,133.77
X$30755 504 613 505 644 645 cell_1rw
* cell instance $30756 m0 *1 154.395,136.5
X$30756 504 615 505 644 645 cell_1rw
* cell instance $30757 r0 *1 154.395,136.5
X$30757 504 614 505 644 645 cell_1rw
* cell instance $30758 m0 *1 154.395,139.23
X$30758 504 617 505 644 645 cell_1rw
* cell instance $30759 r0 *1 154.395,139.23
X$30759 504 616 505 644 645 cell_1rw
* cell instance $30760 m0 *1 154.395,141.96
X$30760 504 618 505 644 645 cell_1rw
* cell instance $30761 r0 *1 154.395,141.96
X$30761 504 619 505 644 645 cell_1rw
* cell instance $30762 m0 *1 154.395,144.69
X$30762 504 620 505 644 645 cell_1rw
* cell instance $30763 r0 *1 154.395,144.69
X$30763 504 621 505 644 645 cell_1rw
* cell instance $30764 m0 *1 154.395,147.42
X$30764 504 622 505 644 645 cell_1rw
* cell instance $30765 r0 *1 154.395,147.42
X$30765 504 623 505 644 645 cell_1rw
* cell instance $30766 m0 *1 154.395,150.15
X$30766 504 624 505 644 645 cell_1rw
* cell instance $30767 r0 *1 154.395,150.15
X$30767 504 625 505 644 645 cell_1rw
* cell instance $30768 m0 *1 154.395,152.88
X$30768 504 626 505 644 645 cell_1rw
* cell instance $30769 r0 *1 154.395,152.88
X$30769 504 627 505 644 645 cell_1rw
* cell instance $30770 m0 *1 154.395,155.61
X$30770 504 628 505 644 645 cell_1rw
* cell instance $30771 m0 *1 154.395,158.34
X$30771 504 630 505 644 645 cell_1rw
* cell instance $30772 r0 *1 154.395,155.61
X$30772 504 629 505 644 645 cell_1rw
* cell instance $30773 r0 *1 154.395,158.34
X$30773 504 631 505 644 645 cell_1rw
* cell instance $30774 m0 *1 154.395,161.07
X$30774 504 632 505 644 645 cell_1rw
* cell instance $30775 r0 *1 154.395,161.07
X$30775 504 633 505 644 645 cell_1rw
* cell instance $30776 m0 *1 154.395,163.8
X$30776 504 634 505 644 645 cell_1rw
* cell instance $30777 r0 *1 154.395,163.8
X$30777 504 635 505 644 645 cell_1rw
* cell instance $30778 m0 *1 154.395,166.53
X$30778 504 637 505 644 645 cell_1rw
* cell instance $30779 r0 *1 154.395,166.53
X$30779 504 636 505 644 645 cell_1rw
* cell instance $30780 m0 *1 154.395,169.26
X$30780 504 639 505 644 645 cell_1rw
* cell instance $30781 r0 *1 154.395,169.26
X$30781 504 638 505 644 645 cell_1rw
* cell instance $30782 m0 *1 154.395,171.99
X$30782 504 640 505 644 645 cell_1rw
* cell instance $30783 r0 *1 154.395,171.99
X$30783 504 641 505 644 645 cell_1rw
* cell instance $30784 m0 *1 154.395,174.72
X$30784 504 642 505 644 645 cell_1rw
* cell instance $30785 r0 *1 154.395,174.72
X$30785 504 643 505 644 645 cell_1rw
* cell instance $30786 m0 *1 155.1,90.09
X$30786 506 581 507 644 645 cell_1rw
* cell instance $30787 r0 *1 155.1,90.09
X$30787 506 580 507 644 645 cell_1rw
* cell instance $30788 m0 *1 155.1,92.82
X$30788 506 583 507 644 645 cell_1rw
* cell instance $30789 r0 *1 155.1,92.82
X$30789 506 582 507 644 645 cell_1rw
* cell instance $30790 m0 *1 155.1,95.55
X$30790 506 584 507 644 645 cell_1rw
* cell instance $30791 r0 *1 155.1,95.55
X$30791 506 585 507 644 645 cell_1rw
* cell instance $30792 m0 *1 155.1,98.28
X$30792 506 586 507 644 645 cell_1rw
* cell instance $30793 r0 *1 155.1,98.28
X$30793 506 587 507 644 645 cell_1rw
* cell instance $30794 m0 *1 155.1,101.01
X$30794 506 588 507 644 645 cell_1rw
* cell instance $30795 r0 *1 155.1,101.01
X$30795 506 589 507 644 645 cell_1rw
* cell instance $30796 m0 *1 155.1,103.74
X$30796 506 590 507 644 645 cell_1rw
* cell instance $30797 r0 *1 155.1,103.74
X$30797 506 591 507 644 645 cell_1rw
* cell instance $30798 m0 *1 155.1,106.47
X$30798 506 593 507 644 645 cell_1rw
* cell instance $30799 r0 *1 155.1,106.47
X$30799 506 592 507 644 645 cell_1rw
* cell instance $30800 m0 *1 155.1,109.2
X$30800 506 594 507 644 645 cell_1rw
* cell instance $30801 r0 *1 155.1,109.2
X$30801 506 595 507 644 645 cell_1rw
* cell instance $30802 m0 *1 155.1,111.93
X$30802 506 597 507 644 645 cell_1rw
* cell instance $30803 m0 *1 155.1,114.66
X$30803 506 598 507 644 645 cell_1rw
* cell instance $30804 r0 *1 155.1,111.93
X$30804 506 596 507 644 645 cell_1rw
* cell instance $30805 r0 *1 155.1,114.66
X$30805 506 599 507 644 645 cell_1rw
* cell instance $30806 m0 *1 155.1,117.39
X$30806 506 600 507 644 645 cell_1rw
* cell instance $30807 m0 *1 155.1,120.12
X$30807 506 602 507 644 645 cell_1rw
* cell instance $30808 r0 *1 155.1,117.39
X$30808 506 601 507 644 645 cell_1rw
* cell instance $30809 m0 *1 155.1,122.85
X$30809 506 604 507 644 645 cell_1rw
* cell instance $30810 r0 *1 155.1,120.12
X$30810 506 603 507 644 645 cell_1rw
* cell instance $30811 r0 *1 155.1,122.85
X$30811 506 605 507 644 645 cell_1rw
* cell instance $30812 m0 *1 155.1,125.58
X$30812 506 606 507 644 645 cell_1rw
* cell instance $30813 r0 *1 155.1,125.58
X$30813 506 607 507 644 645 cell_1rw
* cell instance $30814 m0 *1 155.1,128.31
X$30814 506 609 507 644 645 cell_1rw
* cell instance $30815 m0 *1 155.1,131.04
X$30815 506 610 507 644 645 cell_1rw
* cell instance $30816 r0 *1 155.1,128.31
X$30816 506 608 507 644 645 cell_1rw
* cell instance $30817 r0 *1 155.1,131.04
X$30817 506 611 507 644 645 cell_1rw
* cell instance $30818 m0 *1 155.1,133.77
X$30818 506 612 507 644 645 cell_1rw
* cell instance $30819 r0 *1 155.1,133.77
X$30819 506 613 507 644 645 cell_1rw
* cell instance $30820 m0 *1 155.1,136.5
X$30820 506 615 507 644 645 cell_1rw
* cell instance $30821 r0 *1 155.1,136.5
X$30821 506 614 507 644 645 cell_1rw
* cell instance $30822 m0 *1 155.1,139.23
X$30822 506 617 507 644 645 cell_1rw
* cell instance $30823 r0 *1 155.1,139.23
X$30823 506 616 507 644 645 cell_1rw
* cell instance $30824 m0 *1 155.1,141.96
X$30824 506 618 507 644 645 cell_1rw
* cell instance $30825 r0 *1 155.1,141.96
X$30825 506 619 507 644 645 cell_1rw
* cell instance $30826 m0 *1 155.1,144.69
X$30826 506 620 507 644 645 cell_1rw
* cell instance $30827 r0 *1 155.1,144.69
X$30827 506 621 507 644 645 cell_1rw
* cell instance $30828 m0 *1 155.1,147.42
X$30828 506 622 507 644 645 cell_1rw
* cell instance $30829 r0 *1 155.1,147.42
X$30829 506 623 507 644 645 cell_1rw
* cell instance $30830 m0 *1 155.1,150.15
X$30830 506 624 507 644 645 cell_1rw
* cell instance $30831 m0 *1 155.1,152.88
X$30831 506 626 507 644 645 cell_1rw
* cell instance $30832 r0 *1 155.1,150.15
X$30832 506 625 507 644 645 cell_1rw
* cell instance $30833 r0 *1 155.1,152.88
X$30833 506 627 507 644 645 cell_1rw
* cell instance $30834 m0 *1 155.1,155.61
X$30834 506 628 507 644 645 cell_1rw
* cell instance $30835 m0 *1 155.1,158.34
X$30835 506 630 507 644 645 cell_1rw
* cell instance $30836 r0 *1 155.1,155.61
X$30836 506 629 507 644 645 cell_1rw
* cell instance $30837 r0 *1 155.1,158.34
X$30837 506 631 507 644 645 cell_1rw
* cell instance $30838 m0 *1 155.1,161.07
X$30838 506 632 507 644 645 cell_1rw
* cell instance $30839 r0 *1 155.1,161.07
X$30839 506 633 507 644 645 cell_1rw
* cell instance $30840 m0 *1 155.1,163.8
X$30840 506 634 507 644 645 cell_1rw
* cell instance $30841 r0 *1 155.1,163.8
X$30841 506 635 507 644 645 cell_1rw
* cell instance $30842 m0 *1 155.1,166.53
X$30842 506 637 507 644 645 cell_1rw
* cell instance $30843 r0 *1 155.1,166.53
X$30843 506 636 507 644 645 cell_1rw
* cell instance $30844 m0 *1 155.1,169.26
X$30844 506 639 507 644 645 cell_1rw
* cell instance $30845 r0 *1 155.1,169.26
X$30845 506 638 507 644 645 cell_1rw
* cell instance $30846 m0 *1 155.1,171.99
X$30846 506 640 507 644 645 cell_1rw
* cell instance $30847 r0 *1 155.1,171.99
X$30847 506 641 507 644 645 cell_1rw
* cell instance $30848 m0 *1 155.1,174.72
X$30848 506 642 507 644 645 cell_1rw
* cell instance $30849 r0 *1 155.1,174.72
X$30849 506 643 507 644 645 cell_1rw
* cell instance $30850 m0 *1 155.805,90.09
X$30850 508 581 509 644 645 cell_1rw
* cell instance $30851 r0 *1 155.805,90.09
X$30851 508 580 509 644 645 cell_1rw
* cell instance $30852 m0 *1 155.805,92.82
X$30852 508 583 509 644 645 cell_1rw
* cell instance $30853 r0 *1 155.805,92.82
X$30853 508 582 509 644 645 cell_1rw
* cell instance $30854 m0 *1 155.805,95.55
X$30854 508 584 509 644 645 cell_1rw
* cell instance $30855 r0 *1 155.805,95.55
X$30855 508 585 509 644 645 cell_1rw
* cell instance $30856 m0 *1 155.805,98.28
X$30856 508 586 509 644 645 cell_1rw
* cell instance $30857 r0 *1 155.805,98.28
X$30857 508 587 509 644 645 cell_1rw
* cell instance $30858 m0 *1 155.805,101.01
X$30858 508 588 509 644 645 cell_1rw
* cell instance $30859 r0 *1 155.805,101.01
X$30859 508 589 509 644 645 cell_1rw
* cell instance $30860 m0 *1 155.805,103.74
X$30860 508 590 509 644 645 cell_1rw
* cell instance $30861 r0 *1 155.805,103.74
X$30861 508 591 509 644 645 cell_1rw
* cell instance $30862 m0 *1 155.805,106.47
X$30862 508 593 509 644 645 cell_1rw
* cell instance $30863 r0 *1 155.805,106.47
X$30863 508 592 509 644 645 cell_1rw
* cell instance $30864 m0 *1 155.805,109.2
X$30864 508 594 509 644 645 cell_1rw
* cell instance $30865 r0 *1 155.805,109.2
X$30865 508 595 509 644 645 cell_1rw
* cell instance $30866 m0 *1 155.805,111.93
X$30866 508 597 509 644 645 cell_1rw
* cell instance $30867 m0 *1 155.805,114.66
X$30867 508 598 509 644 645 cell_1rw
* cell instance $30868 r0 *1 155.805,111.93
X$30868 508 596 509 644 645 cell_1rw
* cell instance $30869 r0 *1 155.805,114.66
X$30869 508 599 509 644 645 cell_1rw
* cell instance $30870 m0 *1 155.805,117.39
X$30870 508 600 509 644 645 cell_1rw
* cell instance $30871 m0 *1 155.805,120.12
X$30871 508 602 509 644 645 cell_1rw
* cell instance $30872 r0 *1 155.805,117.39
X$30872 508 601 509 644 645 cell_1rw
* cell instance $30873 r0 *1 155.805,120.12
X$30873 508 603 509 644 645 cell_1rw
* cell instance $30874 m0 *1 155.805,122.85
X$30874 508 604 509 644 645 cell_1rw
* cell instance $30875 r0 *1 155.805,122.85
X$30875 508 605 509 644 645 cell_1rw
* cell instance $30876 m0 *1 155.805,125.58
X$30876 508 606 509 644 645 cell_1rw
* cell instance $30877 r0 *1 155.805,125.58
X$30877 508 607 509 644 645 cell_1rw
* cell instance $30878 m0 *1 155.805,128.31
X$30878 508 609 509 644 645 cell_1rw
* cell instance $30879 r0 *1 155.805,128.31
X$30879 508 608 509 644 645 cell_1rw
* cell instance $30880 m0 *1 155.805,131.04
X$30880 508 610 509 644 645 cell_1rw
* cell instance $30881 r0 *1 155.805,131.04
X$30881 508 611 509 644 645 cell_1rw
* cell instance $30882 m0 *1 155.805,133.77
X$30882 508 612 509 644 645 cell_1rw
* cell instance $30883 r0 *1 155.805,133.77
X$30883 508 613 509 644 645 cell_1rw
* cell instance $30884 m0 *1 155.805,136.5
X$30884 508 615 509 644 645 cell_1rw
* cell instance $30885 r0 *1 155.805,136.5
X$30885 508 614 509 644 645 cell_1rw
* cell instance $30886 m0 *1 155.805,139.23
X$30886 508 617 509 644 645 cell_1rw
* cell instance $30887 r0 *1 155.805,139.23
X$30887 508 616 509 644 645 cell_1rw
* cell instance $30888 m0 *1 155.805,141.96
X$30888 508 618 509 644 645 cell_1rw
* cell instance $30889 r0 *1 155.805,141.96
X$30889 508 619 509 644 645 cell_1rw
* cell instance $30890 m0 *1 155.805,144.69
X$30890 508 620 509 644 645 cell_1rw
* cell instance $30891 r0 *1 155.805,144.69
X$30891 508 621 509 644 645 cell_1rw
* cell instance $30892 m0 *1 155.805,147.42
X$30892 508 622 509 644 645 cell_1rw
* cell instance $30893 r0 *1 155.805,147.42
X$30893 508 623 509 644 645 cell_1rw
* cell instance $30894 m0 *1 155.805,150.15
X$30894 508 624 509 644 645 cell_1rw
* cell instance $30895 r0 *1 155.805,150.15
X$30895 508 625 509 644 645 cell_1rw
* cell instance $30896 m0 *1 155.805,152.88
X$30896 508 626 509 644 645 cell_1rw
* cell instance $30897 r0 *1 155.805,152.88
X$30897 508 627 509 644 645 cell_1rw
* cell instance $30898 m0 *1 155.805,155.61
X$30898 508 628 509 644 645 cell_1rw
* cell instance $30899 m0 *1 155.805,158.34
X$30899 508 630 509 644 645 cell_1rw
* cell instance $30900 r0 *1 155.805,155.61
X$30900 508 629 509 644 645 cell_1rw
* cell instance $30901 r0 *1 155.805,158.34
X$30901 508 631 509 644 645 cell_1rw
* cell instance $30902 m0 *1 155.805,161.07
X$30902 508 632 509 644 645 cell_1rw
* cell instance $30903 m0 *1 155.805,163.8
X$30903 508 634 509 644 645 cell_1rw
* cell instance $30904 r0 *1 155.805,161.07
X$30904 508 633 509 644 645 cell_1rw
* cell instance $30905 r0 *1 155.805,163.8
X$30905 508 635 509 644 645 cell_1rw
* cell instance $30906 m0 *1 155.805,166.53
X$30906 508 637 509 644 645 cell_1rw
* cell instance $30907 r0 *1 155.805,166.53
X$30907 508 636 509 644 645 cell_1rw
* cell instance $30908 m0 *1 155.805,169.26
X$30908 508 639 509 644 645 cell_1rw
* cell instance $30909 r0 *1 155.805,169.26
X$30909 508 638 509 644 645 cell_1rw
* cell instance $30910 m0 *1 155.805,171.99
X$30910 508 640 509 644 645 cell_1rw
* cell instance $30911 r0 *1 155.805,171.99
X$30911 508 641 509 644 645 cell_1rw
* cell instance $30912 m0 *1 155.805,174.72
X$30912 508 642 509 644 645 cell_1rw
* cell instance $30913 r0 *1 155.805,174.72
X$30913 508 643 509 644 645 cell_1rw
* cell instance $30914 m0 *1 156.51,90.09
X$30914 510 581 511 644 645 cell_1rw
* cell instance $30915 m0 *1 156.51,92.82
X$30915 510 583 511 644 645 cell_1rw
* cell instance $30916 r0 *1 156.51,90.09
X$30916 510 580 511 644 645 cell_1rw
* cell instance $30917 r0 *1 156.51,92.82
X$30917 510 582 511 644 645 cell_1rw
* cell instance $30918 m0 *1 156.51,95.55
X$30918 510 584 511 644 645 cell_1rw
* cell instance $30919 r0 *1 156.51,95.55
X$30919 510 585 511 644 645 cell_1rw
* cell instance $30920 m0 *1 156.51,98.28
X$30920 510 586 511 644 645 cell_1rw
* cell instance $30921 r0 *1 156.51,98.28
X$30921 510 587 511 644 645 cell_1rw
* cell instance $30922 m0 *1 156.51,101.01
X$30922 510 588 511 644 645 cell_1rw
* cell instance $30923 r0 *1 156.51,101.01
X$30923 510 589 511 644 645 cell_1rw
* cell instance $30924 m0 *1 156.51,103.74
X$30924 510 590 511 644 645 cell_1rw
* cell instance $30925 r0 *1 156.51,103.74
X$30925 510 591 511 644 645 cell_1rw
* cell instance $30926 m0 *1 156.51,106.47
X$30926 510 593 511 644 645 cell_1rw
* cell instance $30927 r0 *1 156.51,106.47
X$30927 510 592 511 644 645 cell_1rw
* cell instance $30928 m0 *1 156.51,109.2
X$30928 510 594 511 644 645 cell_1rw
* cell instance $30929 r0 *1 156.51,109.2
X$30929 510 595 511 644 645 cell_1rw
* cell instance $30930 m0 *1 156.51,111.93
X$30930 510 597 511 644 645 cell_1rw
* cell instance $30931 r0 *1 156.51,111.93
X$30931 510 596 511 644 645 cell_1rw
* cell instance $30932 m0 *1 156.51,114.66
X$30932 510 598 511 644 645 cell_1rw
* cell instance $30933 r0 *1 156.51,114.66
X$30933 510 599 511 644 645 cell_1rw
* cell instance $30934 m0 *1 156.51,117.39
X$30934 510 600 511 644 645 cell_1rw
* cell instance $30935 r0 *1 156.51,117.39
X$30935 510 601 511 644 645 cell_1rw
* cell instance $30936 m0 *1 156.51,120.12
X$30936 510 602 511 644 645 cell_1rw
* cell instance $30937 r0 *1 156.51,120.12
X$30937 510 603 511 644 645 cell_1rw
* cell instance $30938 m0 *1 156.51,122.85
X$30938 510 604 511 644 645 cell_1rw
* cell instance $30939 r0 *1 156.51,122.85
X$30939 510 605 511 644 645 cell_1rw
* cell instance $30940 m0 *1 156.51,125.58
X$30940 510 606 511 644 645 cell_1rw
* cell instance $30941 r0 *1 156.51,125.58
X$30941 510 607 511 644 645 cell_1rw
* cell instance $30942 m0 *1 156.51,128.31
X$30942 510 609 511 644 645 cell_1rw
* cell instance $30943 r0 *1 156.51,128.31
X$30943 510 608 511 644 645 cell_1rw
* cell instance $30944 m0 *1 156.51,131.04
X$30944 510 610 511 644 645 cell_1rw
* cell instance $30945 r0 *1 156.51,131.04
X$30945 510 611 511 644 645 cell_1rw
* cell instance $30946 m0 *1 156.51,133.77
X$30946 510 612 511 644 645 cell_1rw
* cell instance $30947 r0 *1 156.51,133.77
X$30947 510 613 511 644 645 cell_1rw
* cell instance $30948 m0 *1 156.51,136.5
X$30948 510 615 511 644 645 cell_1rw
* cell instance $30949 r0 *1 156.51,136.5
X$30949 510 614 511 644 645 cell_1rw
* cell instance $30950 m0 *1 156.51,139.23
X$30950 510 617 511 644 645 cell_1rw
* cell instance $30951 r0 *1 156.51,139.23
X$30951 510 616 511 644 645 cell_1rw
* cell instance $30952 m0 *1 156.51,141.96
X$30952 510 618 511 644 645 cell_1rw
* cell instance $30953 r0 *1 156.51,141.96
X$30953 510 619 511 644 645 cell_1rw
* cell instance $30954 m0 *1 156.51,144.69
X$30954 510 620 511 644 645 cell_1rw
* cell instance $30955 r0 *1 156.51,144.69
X$30955 510 621 511 644 645 cell_1rw
* cell instance $30956 m0 *1 156.51,147.42
X$30956 510 622 511 644 645 cell_1rw
* cell instance $30957 r0 *1 156.51,147.42
X$30957 510 623 511 644 645 cell_1rw
* cell instance $30958 m0 *1 156.51,150.15
X$30958 510 624 511 644 645 cell_1rw
* cell instance $30959 r0 *1 156.51,150.15
X$30959 510 625 511 644 645 cell_1rw
* cell instance $30960 m0 *1 156.51,152.88
X$30960 510 626 511 644 645 cell_1rw
* cell instance $30961 r0 *1 156.51,152.88
X$30961 510 627 511 644 645 cell_1rw
* cell instance $30962 m0 *1 156.51,155.61
X$30962 510 628 511 644 645 cell_1rw
* cell instance $30963 r0 *1 156.51,155.61
X$30963 510 629 511 644 645 cell_1rw
* cell instance $30964 m0 *1 156.51,158.34
X$30964 510 630 511 644 645 cell_1rw
* cell instance $30965 r0 *1 156.51,158.34
X$30965 510 631 511 644 645 cell_1rw
* cell instance $30966 m0 *1 156.51,161.07
X$30966 510 632 511 644 645 cell_1rw
* cell instance $30967 r0 *1 156.51,161.07
X$30967 510 633 511 644 645 cell_1rw
* cell instance $30968 m0 *1 156.51,163.8
X$30968 510 634 511 644 645 cell_1rw
* cell instance $30969 m0 *1 156.51,166.53
X$30969 510 637 511 644 645 cell_1rw
* cell instance $30970 r0 *1 156.51,163.8
X$30970 510 635 511 644 645 cell_1rw
* cell instance $30971 r0 *1 156.51,166.53
X$30971 510 636 511 644 645 cell_1rw
* cell instance $30972 m0 *1 156.51,169.26
X$30972 510 639 511 644 645 cell_1rw
* cell instance $30973 r0 *1 156.51,169.26
X$30973 510 638 511 644 645 cell_1rw
* cell instance $30974 m0 *1 156.51,171.99
X$30974 510 640 511 644 645 cell_1rw
* cell instance $30975 r0 *1 156.51,171.99
X$30975 510 641 511 644 645 cell_1rw
* cell instance $30976 m0 *1 156.51,174.72
X$30976 510 642 511 644 645 cell_1rw
* cell instance $30977 r0 *1 156.51,174.72
X$30977 510 643 511 644 645 cell_1rw
* cell instance $30978 m0 *1 157.215,90.09
X$30978 512 581 513 644 645 cell_1rw
* cell instance $30979 r0 *1 157.215,90.09
X$30979 512 580 513 644 645 cell_1rw
* cell instance $30980 m0 *1 157.215,92.82
X$30980 512 583 513 644 645 cell_1rw
* cell instance $30981 r0 *1 157.215,92.82
X$30981 512 582 513 644 645 cell_1rw
* cell instance $30982 m0 *1 157.215,95.55
X$30982 512 584 513 644 645 cell_1rw
* cell instance $30983 r0 *1 157.215,95.55
X$30983 512 585 513 644 645 cell_1rw
* cell instance $30984 m0 *1 157.215,98.28
X$30984 512 586 513 644 645 cell_1rw
* cell instance $30985 r0 *1 157.215,98.28
X$30985 512 587 513 644 645 cell_1rw
* cell instance $30986 m0 *1 157.215,101.01
X$30986 512 588 513 644 645 cell_1rw
* cell instance $30987 r0 *1 157.215,101.01
X$30987 512 589 513 644 645 cell_1rw
* cell instance $30988 m0 *1 157.215,103.74
X$30988 512 590 513 644 645 cell_1rw
* cell instance $30989 r0 *1 157.215,103.74
X$30989 512 591 513 644 645 cell_1rw
* cell instance $30990 m0 *1 157.215,106.47
X$30990 512 593 513 644 645 cell_1rw
* cell instance $30991 r0 *1 157.215,106.47
X$30991 512 592 513 644 645 cell_1rw
* cell instance $30992 m0 *1 157.215,109.2
X$30992 512 594 513 644 645 cell_1rw
* cell instance $30993 r0 *1 157.215,109.2
X$30993 512 595 513 644 645 cell_1rw
* cell instance $30994 m0 *1 157.215,111.93
X$30994 512 597 513 644 645 cell_1rw
* cell instance $30995 r0 *1 157.215,111.93
X$30995 512 596 513 644 645 cell_1rw
* cell instance $30996 m0 *1 157.215,114.66
X$30996 512 598 513 644 645 cell_1rw
* cell instance $30997 r0 *1 157.215,114.66
X$30997 512 599 513 644 645 cell_1rw
* cell instance $30998 m0 *1 157.215,117.39
X$30998 512 600 513 644 645 cell_1rw
* cell instance $30999 r0 *1 157.215,117.39
X$30999 512 601 513 644 645 cell_1rw
* cell instance $31000 m0 *1 157.215,120.12
X$31000 512 602 513 644 645 cell_1rw
* cell instance $31001 r0 *1 157.215,120.12
X$31001 512 603 513 644 645 cell_1rw
* cell instance $31002 m0 *1 157.215,122.85
X$31002 512 604 513 644 645 cell_1rw
* cell instance $31003 r0 *1 157.215,122.85
X$31003 512 605 513 644 645 cell_1rw
* cell instance $31004 m0 *1 157.215,125.58
X$31004 512 606 513 644 645 cell_1rw
* cell instance $31005 r0 *1 157.215,125.58
X$31005 512 607 513 644 645 cell_1rw
* cell instance $31006 m0 *1 157.215,128.31
X$31006 512 609 513 644 645 cell_1rw
* cell instance $31007 r0 *1 157.215,128.31
X$31007 512 608 513 644 645 cell_1rw
* cell instance $31008 m0 *1 157.215,131.04
X$31008 512 610 513 644 645 cell_1rw
* cell instance $31009 r0 *1 157.215,131.04
X$31009 512 611 513 644 645 cell_1rw
* cell instance $31010 m0 *1 157.215,133.77
X$31010 512 612 513 644 645 cell_1rw
* cell instance $31011 r0 *1 157.215,133.77
X$31011 512 613 513 644 645 cell_1rw
* cell instance $31012 m0 *1 157.215,136.5
X$31012 512 615 513 644 645 cell_1rw
* cell instance $31013 r0 *1 157.215,136.5
X$31013 512 614 513 644 645 cell_1rw
* cell instance $31014 m0 *1 157.215,139.23
X$31014 512 617 513 644 645 cell_1rw
* cell instance $31015 r0 *1 157.215,139.23
X$31015 512 616 513 644 645 cell_1rw
* cell instance $31016 m0 *1 157.215,141.96
X$31016 512 618 513 644 645 cell_1rw
* cell instance $31017 r0 *1 157.215,141.96
X$31017 512 619 513 644 645 cell_1rw
* cell instance $31018 m0 *1 157.215,144.69
X$31018 512 620 513 644 645 cell_1rw
* cell instance $31019 r0 *1 157.215,144.69
X$31019 512 621 513 644 645 cell_1rw
* cell instance $31020 m0 *1 157.215,147.42
X$31020 512 622 513 644 645 cell_1rw
* cell instance $31021 r0 *1 157.215,147.42
X$31021 512 623 513 644 645 cell_1rw
* cell instance $31022 m0 *1 157.215,150.15
X$31022 512 624 513 644 645 cell_1rw
* cell instance $31023 r0 *1 157.215,150.15
X$31023 512 625 513 644 645 cell_1rw
* cell instance $31024 m0 *1 157.215,152.88
X$31024 512 626 513 644 645 cell_1rw
* cell instance $31025 m0 *1 157.215,155.61
X$31025 512 628 513 644 645 cell_1rw
* cell instance $31026 r0 *1 157.215,152.88
X$31026 512 627 513 644 645 cell_1rw
* cell instance $31027 r0 *1 157.215,155.61
X$31027 512 629 513 644 645 cell_1rw
* cell instance $31028 m0 *1 157.215,158.34
X$31028 512 630 513 644 645 cell_1rw
* cell instance $31029 r0 *1 157.215,158.34
X$31029 512 631 513 644 645 cell_1rw
* cell instance $31030 m0 *1 157.215,161.07
X$31030 512 632 513 644 645 cell_1rw
* cell instance $31031 r0 *1 157.215,161.07
X$31031 512 633 513 644 645 cell_1rw
* cell instance $31032 m0 *1 157.215,163.8
X$31032 512 634 513 644 645 cell_1rw
* cell instance $31033 r0 *1 157.215,163.8
X$31033 512 635 513 644 645 cell_1rw
* cell instance $31034 m0 *1 157.215,166.53
X$31034 512 637 513 644 645 cell_1rw
* cell instance $31035 r0 *1 157.215,166.53
X$31035 512 636 513 644 645 cell_1rw
* cell instance $31036 m0 *1 157.215,169.26
X$31036 512 639 513 644 645 cell_1rw
* cell instance $31037 r0 *1 157.215,169.26
X$31037 512 638 513 644 645 cell_1rw
* cell instance $31038 m0 *1 157.215,171.99
X$31038 512 640 513 644 645 cell_1rw
* cell instance $31039 m0 *1 157.215,174.72
X$31039 512 642 513 644 645 cell_1rw
* cell instance $31040 r0 *1 157.215,171.99
X$31040 512 641 513 644 645 cell_1rw
* cell instance $31041 r0 *1 157.215,174.72
X$31041 512 643 513 644 645 cell_1rw
* cell instance $31042 m0 *1 157.92,90.09
X$31042 514 581 515 644 645 cell_1rw
* cell instance $31043 r0 *1 157.92,90.09
X$31043 514 580 515 644 645 cell_1rw
* cell instance $31044 m0 *1 157.92,92.82
X$31044 514 583 515 644 645 cell_1rw
* cell instance $31045 r0 *1 157.92,92.82
X$31045 514 582 515 644 645 cell_1rw
* cell instance $31046 m0 *1 157.92,95.55
X$31046 514 584 515 644 645 cell_1rw
* cell instance $31047 r0 *1 157.92,95.55
X$31047 514 585 515 644 645 cell_1rw
* cell instance $31048 m0 *1 157.92,98.28
X$31048 514 586 515 644 645 cell_1rw
* cell instance $31049 m0 *1 157.92,101.01
X$31049 514 588 515 644 645 cell_1rw
* cell instance $31050 r0 *1 157.92,98.28
X$31050 514 587 515 644 645 cell_1rw
* cell instance $31051 m0 *1 157.92,103.74
X$31051 514 590 515 644 645 cell_1rw
* cell instance $31052 r0 *1 157.92,101.01
X$31052 514 589 515 644 645 cell_1rw
* cell instance $31053 r0 *1 157.92,103.74
X$31053 514 591 515 644 645 cell_1rw
* cell instance $31054 m0 *1 157.92,106.47
X$31054 514 593 515 644 645 cell_1rw
* cell instance $31055 r0 *1 157.92,106.47
X$31055 514 592 515 644 645 cell_1rw
* cell instance $31056 m0 *1 157.92,109.2
X$31056 514 594 515 644 645 cell_1rw
* cell instance $31057 r0 *1 157.92,109.2
X$31057 514 595 515 644 645 cell_1rw
* cell instance $31058 m0 *1 157.92,111.93
X$31058 514 597 515 644 645 cell_1rw
* cell instance $31059 m0 *1 157.92,114.66
X$31059 514 598 515 644 645 cell_1rw
* cell instance $31060 r0 *1 157.92,111.93
X$31060 514 596 515 644 645 cell_1rw
* cell instance $31061 r0 *1 157.92,114.66
X$31061 514 599 515 644 645 cell_1rw
* cell instance $31062 m0 *1 157.92,117.39
X$31062 514 600 515 644 645 cell_1rw
* cell instance $31063 r0 *1 157.92,117.39
X$31063 514 601 515 644 645 cell_1rw
* cell instance $31064 m0 *1 157.92,120.12
X$31064 514 602 515 644 645 cell_1rw
* cell instance $31065 r0 *1 157.92,120.12
X$31065 514 603 515 644 645 cell_1rw
* cell instance $31066 m0 *1 157.92,122.85
X$31066 514 604 515 644 645 cell_1rw
* cell instance $31067 r0 *1 157.92,122.85
X$31067 514 605 515 644 645 cell_1rw
* cell instance $31068 m0 *1 157.92,125.58
X$31068 514 606 515 644 645 cell_1rw
* cell instance $31069 m0 *1 157.92,128.31
X$31069 514 609 515 644 645 cell_1rw
* cell instance $31070 r0 *1 157.92,125.58
X$31070 514 607 515 644 645 cell_1rw
* cell instance $31071 m0 *1 157.92,131.04
X$31071 514 610 515 644 645 cell_1rw
* cell instance $31072 r0 *1 157.92,128.31
X$31072 514 608 515 644 645 cell_1rw
* cell instance $31073 r0 *1 157.92,131.04
X$31073 514 611 515 644 645 cell_1rw
* cell instance $31074 m0 *1 157.92,133.77
X$31074 514 612 515 644 645 cell_1rw
* cell instance $31075 r0 *1 157.92,133.77
X$31075 514 613 515 644 645 cell_1rw
* cell instance $31076 m0 *1 157.92,136.5
X$31076 514 615 515 644 645 cell_1rw
* cell instance $31077 r0 *1 157.92,136.5
X$31077 514 614 515 644 645 cell_1rw
* cell instance $31078 m0 *1 157.92,139.23
X$31078 514 617 515 644 645 cell_1rw
* cell instance $31079 r0 *1 157.92,139.23
X$31079 514 616 515 644 645 cell_1rw
* cell instance $31080 m0 *1 157.92,141.96
X$31080 514 618 515 644 645 cell_1rw
* cell instance $31081 r0 *1 157.92,141.96
X$31081 514 619 515 644 645 cell_1rw
* cell instance $31082 m0 *1 157.92,144.69
X$31082 514 620 515 644 645 cell_1rw
* cell instance $31083 r0 *1 157.92,144.69
X$31083 514 621 515 644 645 cell_1rw
* cell instance $31084 m0 *1 157.92,147.42
X$31084 514 622 515 644 645 cell_1rw
* cell instance $31085 r0 *1 157.92,147.42
X$31085 514 623 515 644 645 cell_1rw
* cell instance $31086 m0 *1 157.92,150.15
X$31086 514 624 515 644 645 cell_1rw
* cell instance $31087 r0 *1 157.92,150.15
X$31087 514 625 515 644 645 cell_1rw
* cell instance $31088 m0 *1 157.92,152.88
X$31088 514 626 515 644 645 cell_1rw
* cell instance $31089 r0 *1 157.92,152.88
X$31089 514 627 515 644 645 cell_1rw
* cell instance $31090 m0 *1 157.92,155.61
X$31090 514 628 515 644 645 cell_1rw
* cell instance $31091 r0 *1 157.92,155.61
X$31091 514 629 515 644 645 cell_1rw
* cell instance $31092 m0 *1 157.92,158.34
X$31092 514 630 515 644 645 cell_1rw
* cell instance $31093 r0 *1 157.92,158.34
X$31093 514 631 515 644 645 cell_1rw
* cell instance $31094 m0 *1 157.92,161.07
X$31094 514 632 515 644 645 cell_1rw
* cell instance $31095 r0 *1 157.92,161.07
X$31095 514 633 515 644 645 cell_1rw
* cell instance $31096 m0 *1 157.92,163.8
X$31096 514 634 515 644 645 cell_1rw
* cell instance $31097 m0 *1 157.92,166.53
X$31097 514 637 515 644 645 cell_1rw
* cell instance $31098 r0 *1 157.92,163.8
X$31098 514 635 515 644 645 cell_1rw
* cell instance $31099 r0 *1 157.92,166.53
X$31099 514 636 515 644 645 cell_1rw
* cell instance $31100 m0 *1 157.92,169.26
X$31100 514 639 515 644 645 cell_1rw
* cell instance $31101 r0 *1 157.92,169.26
X$31101 514 638 515 644 645 cell_1rw
* cell instance $31102 m0 *1 157.92,171.99
X$31102 514 640 515 644 645 cell_1rw
* cell instance $31103 m0 *1 157.92,174.72
X$31103 514 642 515 644 645 cell_1rw
* cell instance $31104 r0 *1 157.92,171.99
X$31104 514 641 515 644 645 cell_1rw
* cell instance $31105 r0 *1 157.92,174.72
X$31105 514 643 515 644 645 cell_1rw
* cell instance $31106 m0 *1 158.625,90.09
X$31106 516 581 517 644 645 cell_1rw
* cell instance $31107 r0 *1 158.625,90.09
X$31107 516 580 517 644 645 cell_1rw
* cell instance $31108 m0 *1 158.625,92.82
X$31108 516 583 517 644 645 cell_1rw
* cell instance $31109 r0 *1 158.625,92.82
X$31109 516 582 517 644 645 cell_1rw
* cell instance $31110 m0 *1 158.625,95.55
X$31110 516 584 517 644 645 cell_1rw
* cell instance $31111 r0 *1 158.625,95.55
X$31111 516 585 517 644 645 cell_1rw
* cell instance $31112 m0 *1 158.625,98.28
X$31112 516 586 517 644 645 cell_1rw
* cell instance $31113 r0 *1 158.625,98.28
X$31113 516 587 517 644 645 cell_1rw
* cell instance $31114 m0 *1 158.625,101.01
X$31114 516 588 517 644 645 cell_1rw
* cell instance $31115 r0 *1 158.625,101.01
X$31115 516 589 517 644 645 cell_1rw
* cell instance $31116 m0 *1 158.625,103.74
X$31116 516 590 517 644 645 cell_1rw
* cell instance $31117 r0 *1 158.625,103.74
X$31117 516 591 517 644 645 cell_1rw
* cell instance $31118 m0 *1 158.625,106.47
X$31118 516 593 517 644 645 cell_1rw
* cell instance $31119 m0 *1 158.625,109.2
X$31119 516 594 517 644 645 cell_1rw
* cell instance $31120 r0 *1 158.625,106.47
X$31120 516 592 517 644 645 cell_1rw
* cell instance $31121 r0 *1 158.625,109.2
X$31121 516 595 517 644 645 cell_1rw
* cell instance $31122 m0 *1 158.625,111.93
X$31122 516 597 517 644 645 cell_1rw
* cell instance $31123 r0 *1 158.625,111.93
X$31123 516 596 517 644 645 cell_1rw
* cell instance $31124 m0 *1 158.625,114.66
X$31124 516 598 517 644 645 cell_1rw
* cell instance $31125 r0 *1 158.625,114.66
X$31125 516 599 517 644 645 cell_1rw
* cell instance $31126 m0 *1 158.625,117.39
X$31126 516 600 517 644 645 cell_1rw
* cell instance $31127 r0 *1 158.625,117.39
X$31127 516 601 517 644 645 cell_1rw
* cell instance $31128 m0 *1 158.625,120.12
X$31128 516 602 517 644 645 cell_1rw
* cell instance $31129 r0 *1 158.625,120.12
X$31129 516 603 517 644 645 cell_1rw
* cell instance $31130 m0 *1 158.625,122.85
X$31130 516 604 517 644 645 cell_1rw
* cell instance $31131 r0 *1 158.625,122.85
X$31131 516 605 517 644 645 cell_1rw
* cell instance $31132 m0 *1 158.625,125.58
X$31132 516 606 517 644 645 cell_1rw
* cell instance $31133 r0 *1 158.625,125.58
X$31133 516 607 517 644 645 cell_1rw
* cell instance $31134 m0 *1 158.625,128.31
X$31134 516 609 517 644 645 cell_1rw
* cell instance $31135 r0 *1 158.625,128.31
X$31135 516 608 517 644 645 cell_1rw
* cell instance $31136 m0 *1 158.625,131.04
X$31136 516 610 517 644 645 cell_1rw
* cell instance $31137 r0 *1 158.625,131.04
X$31137 516 611 517 644 645 cell_1rw
* cell instance $31138 m0 *1 158.625,133.77
X$31138 516 612 517 644 645 cell_1rw
* cell instance $31139 r0 *1 158.625,133.77
X$31139 516 613 517 644 645 cell_1rw
* cell instance $31140 m0 *1 158.625,136.5
X$31140 516 615 517 644 645 cell_1rw
* cell instance $31141 r0 *1 158.625,136.5
X$31141 516 614 517 644 645 cell_1rw
* cell instance $31142 m0 *1 158.625,139.23
X$31142 516 617 517 644 645 cell_1rw
* cell instance $31143 r0 *1 158.625,139.23
X$31143 516 616 517 644 645 cell_1rw
* cell instance $31144 m0 *1 158.625,141.96
X$31144 516 618 517 644 645 cell_1rw
* cell instance $31145 r0 *1 158.625,141.96
X$31145 516 619 517 644 645 cell_1rw
* cell instance $31146 m0 *1 158.625,144.69
X$31146 516 620 517 644 645 cell_1rw
* cell instance $31147 r0 *1 158.625,144.69
X$31147 516 621 517 644 645 cell_1rw
* cell instance $31148 m0 *1 158.625,147.42
X$31148 516 622 517 644 645 cell_1rw
* cell instance $31149 r0 *1 158.625,147.42
X$31149 516 623 517 644 645 cell_1rw
* cell instance $31150 m0 *1 158.625,150.15
X$31150 516 624 517 644 645 cell_1rw
* cell instance $31151 r0 *1 158.625,150.15
X$31151 516 625 517 644 645 cell_1rw
* cell instance $31152 m0 *1 158.625,152.88
X$31152 516 626 517 644 645 cell_1rw
* cell instance $31153 r0 *1 158.625,152.88
X$31153 516 627 517 644 645 cell_1rw
* cell instance $31154 m0 *1 158.625,155.61
X$31154 516 628 517 644 645 cell_1rw
* cell instance $31155 r0 *1 158.625,155.61
X$31155 516 629 517 644 645 cell_1rw
* cell instance $31156 m0 *1 158.625,158.34
X$31156 516 630 517 644 645 cell_1rw
* cell instance $31157 r0 *1 158.625,158.34
X$31157 516 631 517 644 645 cell_1rw
* cell instance $31158 m0 *1 158.625,161.07
X$31158 516 632 517 644 645 cell_1rw
* cell instance $31159 m0 *1 158.625,163.8
X$31159 516 634 517 644 645 cell_1rw
* cell instance $31160 r0 *1 158.625,161.07
X$31160 516 633 517 644 645 cell_1rw
* cell instance $31161 r0 *1 158.625,163.8
X$31161 516 635 517 644 645 cell_1rw
* cell instance $31162 m0 *1 158.625,166.53
X$31162 516 637 517 644 645 cell_1rw
* cell instance $31163 r0 *1 158.625,166.53
X$31163 516 636 517 644 645 cell_1rw
* cell instance $31164 m0 *1 158.625,169.26
X$31164 516 639 517 644 645 cell_1rw
* cell instance $31165 r0 *1 158.625,169.26
X$31165 516 638 517 644 645 cell_1rw
* cell instance $31166 m0 *1 158.625,171.99
X$31166 516 640 517 644 645 cell_1rw
* cell instance $31167 r0 *1 158.625,171.99
X$31167 516 641 517 644 645 cell_1rw
* cell instance $31168 m0 *1 158.625,174.72
X$31168 516 642 517 644 645 cell_1rw
* cell instance $31169 r0 *1 158.625,174.72
X$31169 516 643 517 644 645 cell_1rw
* cell instance $31170 m0 *1 159.33,90.09
X$31170 518 581 519 644 645 cell_1rw
* cell instance $31171 r0 *1 159.33,90.09
X$31171 518 580 519 644 645 cell_1rw
* cell instance $31172 m0 *1 159.33,92.82
X$31172 518 583 519 644 645 cell_1rw
* cell instance $31173 r0 *1 159.33,92.82
X$31173 518 582 519 644 645 cell_1rw
* cell instance $31174 m0 *1 159.33,95.55
X$31174 518 584 519 644 645 cell_1rw
* cell instance $31175 r0 *1 159.33,95.55
X$31175 518 585 519 644 645 cell_1rw
* cell instance $31176 m0 *1 159.33,98.28
X$31176 518 586 519 644 645 cell_1rw
* cell instance $31177 r0 *1 159.33,98.28
X$31177 518 587 519 644 645 cell_1rw
* cell instance $31178 m0 *1 159.33,101.01
X$31178 518 588 519 644 645 cell_1rw
* cell instance $31179 r0 *1 159.33,101.01
X$31179 518 589 519 644 645 cell_1rw
* cell instance $31180 m0 *1 159.33,103.74
X$31180 518 590 519 644 645 cell_1rw
* cell instance $31181 r0 *1 159.33,103.74
X$31181 518 591 519 644 645 cell_1rw
* cell instance $31182 m0 *1 159.33,106.47
X$31182 518 593 519 644 645 cell_1rw
* cell instance $31183 m0 *1 159.33,109.2
X$31183 518 594 519 644 645 cell_1rw
* cell instance $31184 r0 *1 159.33,106.47
X$31184 518 592 519 644 645 cell_1rw
* cell instance $31185 m0 *1 159.33,111.93
X$31185 518 597 519 644 645 cell_1rw
* cell instance $31186 r0 *1 159.33,109.2
X$31186 518 595 519 644 645 cell_1rw
* cell instance $31187 r0 *1 159.33,111.93
X$31187 518 596 519 644 645 cell_1rw
* cell instance $31188 m0 *1 159.33,114.66
X$31188 518 598 519 644 645 cell_1rw
* cell instance $31189 r0 *1 159.33,114.66
X$31189 518 599 519 644 645 cell_1rw
* cell instance $31190 m0 *1 159.33,117.39
X$31190 518 600 519 644 645 cell_1rw
* cell instance $31191 m0 *1 159.33,120.12
X$31191 518 602 519 644 645 cell_1rw
* cell instance $31192 r0 *1 159.33,117.39
X$31192 518 601 519 644 645 cell_1rw
* cell instance $31193 r0 *1 159.33,120.12
X$31193 518 603 519 644 645 cell_1rw
* cell instance $31194 m0 *1 159.33,122.85
X$31194 518 604 519 644 645 cell_1rw
* cell instance $31195 r0 *1 159.33,122.85
X$31195 518 605 519 644 645 cell_1rw
* cell instance $31196 m0 *1 159.33,125.58
X$31196 518 606 519 644 645 cell_1rw
* cell instance $31197 r0 *1 159.33,125.58
X$31197 518 607 519 644 645 cell_1rw
* cell instance $31198 m0 *1 159.33,128.31
X$31198 518 609 519 644 645 cell_1rw
* cell instance $31199 r0 *1 159.33,128.31
X$31199 518 608 519 644 645 cell_1rw
* cell instance $31200 m0 *1 159.33,131.04
X$31200 518 610 519 644 645 cell_1rw
* cell instance $31201 r0 *1 159.33,131.04
X$31201 518 611 519 644 645 cell_1rw
* cell instance $31202 m0 *1 159.33,133.77
X$31202 518 612 519 644 645 cell_1rw
* cell instance $31203 r0 *1 159.33,133.77
X$31203 518 613 519 644 645 cell_1rw
* cell instance $31204 m0 *1 159.33,136.5
X$31204 518 615 519 644 645 cell_1rw
* cell instance $31205 r0 *1 159.33,136.5
X$31205 518 614 519 644 645 cell_1rw
* cell instance $31206 m0 *1 159.33,139.23
X$31206 518 617 519 644 645 cell_1rw
* cell instance $31207 m0 *1 159.33,141.96
X$31207 518 618 519 644 645 cell_1rw
* cell instance $31208 r0 *1 159.33,139.23
X$31208 518 616 519 644 645 cell_1rw
* cell instance $31209 r0 *1 159.33,141.96
X$31209 518 619 519 644 645 cell_1rw
* cell instance $31210 m0 *1 159.33,144.69
X$31210 518 620 519 644 645 cell_1rw
* cell instance $31211 r0 *1 159.33,144.69
X$31211 518 621 519 644 645 cell_1rw
* cell instance $31212 m0 *1 159.33,147.42
X$31212 518 622 519 644 645 cell_1rw
* cell instance $31213 m0 *1 159.33,150.15
X$31213 518 624 519 644 645 cell_1rw
* cell instance $31214 r0 *1 159.33,147.42
X$31214 518 623 519 644 645 cell_1rw
* cell instance $31215 r0 *1 159.33,150.15
X$31215 518 625 519 644 645 cell_1rw
* cell instance $31216 m0 *1 159.33,152.88
X$31216 518 626 519 644 645 cell_1rw
* cell instance $31217 r0 *1 159.33,152.88
X$31217 518 627 519 644 645 cell_1rw
* cell instance $31218 m0 *1 159.33,155.61
X$31218 518 628 519 644 645 cell_1rw
* cell instance $31219 m0 *1 159.33,158.34
X$31219 518 630 519 644 645 cell_1rw
* cell instance $31220 r0 *1 159.33,155.61
X$31220 518 629 519 644 645 cell_1rw
* cell instance $31221 r0 *1 159.33,158.34
X$31221 518 631 519 644 645 cell_1rw
* cell instance $31222 m0 *1 159.33,161.07
X$31222 518 632 519 644 645 cell_1rw
* cell instance $31223 r0 *1 159.33,161.07
X$31223 518 633 519 644 645 cell_1rw
* cell instance $31224 m0 *1 159.33,163.8
X$31224 518 634 519 644 645 cell_1rw
* cell instance $31225 r0 *1 159.33,163.8
X$31225 518 635 519 644 645 cell_1rw
* cell instance $31226 m0 *1 159.33,166.53
X$31226 518 637 519 644 645 cell_1rw
* cell instance $31227 r0 *1 159.33,166.53
X$31227 518 636 519 644 645 cell_1rw
* cell instance $31228 m0 *1 159.33,169.26
X$31228 518 639 519 644 645 cell_1rw
* cell instance $31229 r0 *1 159.33,169.26
X$31229 518 638 519 644 645 cell_1rw
* cell instance $31230 m0 *1 159.33,171.99
X$31230 518 640 519 644 645 cell_1rw
* cell instance $31231 r0 *1 159.33,171.99
X$31231 518 641 519 644 645 cell_1rw
* cell instance $31232 m0 *1 159.33,174.72
X$31232 518 642 519 644 645 cell_1rw
* cell instance $31233 r0 *1 159.33,174.72
X$31233 518 643 519 644 645 cell_1rw
* cell instance $31234 m0 *1 160.035,90.09
X$31234 520 581 521 644 645 cell_1rw
* cell instance $31235 m0 *1 160.035,92.82
X$31235 520 583 521 644 645 cell_1rw
* cell instance $31236 r0 *1 160.035,90.09
X$31236 520 580 521 644 645 cell_1rw
* cell instance $31237 r0 *1 160.035,92.82
X$31237 520 582 521 644 645 cell_1rw
* cell instance $31238 m0 *1 160.035,95.55
X$31238 520 584 521 644 645 cell_1rw
* cell instance $31239 r0 *1 160.035,95.55
X$31239 520 585 521 644 645 cell_1rw
* cell instance $31240 m0 *1 160.035,98.28
X$31240 520 586 521 644 645 cell_1rw
* cell instance $31241 m0 *1 160.035,101.01
X$31241 520 588 521 644 645 cell_1rw
* cell instance $31242 r0 *1 160.035,98.28
X$31242 520 587 521 644 645 cell_1rw
* cell instance $31243 m0 *1 160.035,103.74
X$31243 520 590 521 644 645 cell_1rw
* cell instance $31244 r0 *1 160.035,101.01
X$31244 520 589 521 644 645 cell_1rw
* cell instance $31245 r0 *1 160.035,103.74
X$31245 520 591 521 644 645 cell_1rw
* cell instance $31246 m0 *1 160.035,106.47
X$31246 520 593 521 644 645 cell_1rw
* cell instance $31247 r0 *1 160.035,106.47
X$31247 520 592 521 644 645 cell_1rw
* cell instance $31248 m0 *1 160.035,109.2
X$31248 520 594 521 644 645 cell_1rw
* cell instance $31249 r0 *1 160.035,109.2
X$31249 520 595 521 644 645 cell_1rw
* cell instance $31250 m0 *1 160.035,111.93
X$31250 520 597 521 644 645 cell_1rw
* cell instance $31251 m0 *1 160.035,114.66
X$31251 520 598 521 644 645 cell_1rw
* cell instance $31252 r0 *1 160.035,111.93
X$31252 520 596 521 644 645 cell_1rw
* cell instance $31253 r0 *1 160.035,114.66
X$31253 520 599 521 644 645 cell_1rw
* cell instance $31254 m0 *1 160.035,117.39
X$31254 520 600 521 644 645 cell_1rw
* cell instance $31255 m0 *1 160.035,120.12
X$31255 520 602 521 644 645 cell_1rw
* cell instance $31256 r0 *1 160.035,117.39
X$31256 520 601 521 644 645 cell_1rw
* cell instance $31257 r0 *1 160.035,120.12
X$31257 520 603 521 644 645 cell_1rw
* cell instance $31258 m0 *1 160.035,122.85
X$31258 520 604 521 644 645 cell_1rw
* cell instance $31259 r0 *1 160.035,122.85
X$31259 520 605 521 644 645 cell_1rw
* cell instance $31260 m0 *1 160.035,125.58
X$31260 520 606 521 644 645 cell_1rw
* cell instance $31261 m0 *1 160.035,128.31
X$31261 520 609 521 644 645 cell_1rw
* cell instance $31262 r0 *1 160.035,125.58
X$31262 520 607 521 644 645 cell_1rw
* cell instance $31263 r0 *1 160.035,128.31
X$31263 520 608 521 644 645 cell_1rw
* cell instance $31264 m0 *1 160.035,131.04
X$31264 520 610 521 644 645 cell_1rw
* cell instance $31265 m0 *1 160.035,133.77
X$31265 520 612 521 644 645 cell_1rw
* cell instance $31266 r0 *1 160.035,131.04
X$31266 520 611 521 644 645 cell_1rw
* cell instance $31267 r0 *1 160.035,133.77
X$31267 520 613 521 644 645 cell_1rw
* cell instance $31268 m0 *1 160.035,136.5
X$31268 520 615 521 644 645 cell_1rw
* cell instance $31269 r0 *1 160.035,136.5
X$31269 520 614 521 644 645 cell_1rw
* cell instance $31270 m0 *1 160.035,139.23
X$31270 520 617 521 644 645 cell_1rw
* cell instance $31271 r0 *1 160.035,139.23
X$31271 520 616 521 644 645 cell_1rw
* cell instance $31272 m0 *1 160.035,141.96
X$31272 520 618 521 644 645 cell_1rw
* cell instance $31273 r0 *1 160.035,141.96
X$31273 520 619 521 644 645 cell_1rw
* cell instance $31274 m0 *1 160.035,144.69
X$31274 520 620 521 644 645 cell_1rw
* cell instance $31275 r0 *1 160.035,144.69
X$31275 520 621 521 644 645 cell_1rw
* cell instance $31276 m0 *1 160.035,147.42
X$31276 520 622 521 644 645 cell_1rw
* cell instance $31277 r0 *1 160.035,147.42
X$31277 520 623 521 644 645 cell_1rw
* cell instance $31278 m0 *1 160.035,150.15
X$31278 520 624 521 644 645 cell_1rw
* cell instance $31279 r0 *1 160.035,150.15
X$31279 520 625 521 644 645 cell_1rw
* cell instance $31280 m0 *1 160.035,152.88
X$31280 520 626 521 644 645 cell_1rw
* cell instance $31281 r0 *1 160.035,152.88
X$31281 520 627 521 644 645 cell_1rw
* cell instance $31282 m0 *1 160.035,155.61
X$31282 520 628 521 644 645 cell_1rw
* cell instance $31283 r0 *1 160.035,155.61
X$31283 520 629 521 644 645 cell_1rw
* cell instance $31284 m0 *1 160.035,158.34
X$31284 520 630 521 644 645 cell_1rw
* cell instance $31285 r0 *1 160.035,158.34
X$31285 520 631 521 644 645 cell_1rw
* cell instance $31286 m0 *1 160.035,161.07
X$31286 520 632 521 644 645 cell_1rw
* cell instance $31287 r0 *1 160.035,161.07
X$31287 520 633 521 644 645 cell_1rw
* cell instance $31288 m0 *1 160.035,163.8
X$31288 520 634 521 644 645 cell_1rw
* cell instance $31289 r0 *1 160.035,163.8
X$31289 520 635 521 644 645 cell_1rw
* cell instance $31290 m0 *1 160.035,166.53
X$31290 520 637 521 644 645 cell_1rw
* cell instance $31291 r0 *1 160.035,166.53
X$31291 520 636 521 644 645 cell_1rw
* cell instance $31292 m0 *1 160.035,169.26
X$31292 520 639 521 644 645 cell_1rw
* cell instance $31293 r0 *1 160.035,169.26
X$31293 520 638 521 644 645 cell_1rw
* cell instance $31294 m0 *1 160.035,171.99
X$31294 520 640 521 644 645 cell_1rw
* cell instance $31295 r0 *1 160.035,171.99
X$31295 520 641 521 644 645 cell_1rw
* cell instance $31296 m0 *1 160.035,174.72
X$31296 520 642 521 644 645 cell_1rw
* cell instance $31297 r0 *1 160.035,174.72
X$31297 520 643 521 644 645 cell_1rw
* cell instance $31298 m0 *1 160.74,90.09
X$31298 522 581 523 644 645 cell_1rw
* cell instance $31299 r0 *1 160.74,90.09
X$31299 522 580 523 644 645 cell_1rw
* cell instance $31300 m0 *1 160.74,92.82
X$31300 522 583 523 644 645 cell_1rw
* cell instance $31301 r0 *1 160.74,92.82
X$31301 522 582 523 644 645 cell_1rw
* cell instance $31302 m0 *1 160.74,95.55
X$31302 522 584 523 644 645 cell_1rw
* cell instance $31303 r0 *1 160.74,95.55
X$31303 522 585 523 644 645 cell_1rw
* cell instance $31304 m0 *1 160.74,98.28
X$31304 522 586 523 644 645 cell_1rw
* cell instance $31305 r0 *1 160.74,98.28
X$31305 522 587 523 644 645 cell_1rw
* cell instance $31306 m0 *1 160.74,101.01
X$31306 522 588 523 644 645 cell_1rw
* cell instance $31307 r0 *1 160.74,101.01
X$31307 522 589 523 644 645 cell_1rw
* cell instance $31308 m0 *1 160.74,103.74
X$31308 522 590 523 644 645 cell_1rw
* cell instance $31309 r0 *1 160.74,103.74
X$31309 522 591 523 644 645 cell_1rw
* cell instance $31310 m0 *1 160.74,106.47
X$31310 522 593 523 644 645 cell_1rw
* cell instance $31311 r0 *1 160.74,106.47
X$31311 522 592 523 644 645 cell_1rw
* cell instance $31312 m0 *1 160.74,109.2
X$31312 522 594 523 644 645 cell_1rw
* cell instance $31313 r0 *1 160.74,109.2
X$31313 522 595 523 644 645 cell_1rw
* cell instance $31314 m0 *1 160.74,111.93
X$31314 522 597 523 644 645 cell_1rw
* cell instance $31315 r0 *1 160.74,111.93
X$31315 522 596 523 644 645 cell_1rw
* cell instance $31316 m0 *1 160.74,114.66
X$31316 522 598 523 644 645 cell_1rw
* cell instance $31317 r0 *1 160.74,114.66
X$31317 522 599 523 644 645 cell_1rw
* cell instance $31318 m0 *1 160.74,117.39
X$31318 522 600 523 644 645 cell_1rw
* cell instance $31319 r0 *1 160.74,117.39
X$31319 522 601 523 644 645 cell_1rw
* cell instance $31320 m0 *1 160.74,120.12
X$31320 522 602 523 644 645 cell_1rw
* cell instance $31321 r0 *1 160.74,120.12
X$31321 522 603 523 644 645 cell_1rw
* cell instance $31322 m0 *1 160.74,122.85
X$31322 522 604 523 644 645 cell_1rw
* cell instance $31323 r0 *1 160.74,122.85
X$31323 522 605 523 644 645 cell_1rw
* cell instance $31324 m0 *1 160.74,125.58
X$31324 522 606 523 644 645 cell_1rw
* cell instance $31325 r0 *1 160.74,125.58
X$31325 522 607 523 644 645 cell_1rw
* cell instance $31326 m0 *1 160.74,128.31
X$31326 522 609 523 644 645 cell_1rw
* cell instance $31327 r0 *1 160.74,128.31
X$31327 522 608 523 644 645 cell_1rw
* cell instance $31328 m0 *1 160.74,131.04
X$31328 522 610 523 644 645 cell_1rw
* cell instance $31329 m0 *1 160.74,133.77
X$31329 522 612 523 644 645 cell_1rw
* cell instance $31330 r0 *1 160.74,131.04
X$31330 522 611 523 644 645 cell_1rw
* cell instance $31331 r0 *1 160.74,133.77
X$31331 522 613 523 644 645 cell_1rw
* cell instance $31332 m0 *1 160.74,136.5
X$31332 522 615 523 644 645 cell_1rw
* cell instance $31333 r0 *1 160.74,136.5
X$31333 522 614 523 644 645 cell_1rw
* cell instance $31334 m0 *1 160.74,139.23
X$31334 522 617 523 644 645 cell_1rw
* cell instance $31335 r0 *1 160.74,139.23
X$31335 522 616 523 644 645 cell_1rw
* cell instance $31336 m0 *1 160.74,141.96
X$31336 522 618 523 644 645 cell_1rw
* cell instance $31337 r0 *1 160.74,141.96
X$31337 522 619 523 644 645 cell_1rw
* cell instance $31338 m0 *1 160.74,144.69
X$31338 522 620 523 644 645 cell_1rw
* cell instance $31339 r0 *1 160.74,144.69
X$31339 522 621 523 644 645 cell_1rw
* cell instance $31340 m0 *1 160.74,147.42
X$31340 522 622 523 644 645 cell_1rw
* cell instance $31341 m0 *1 160.74,150.15
X$31341 522 624 523 644 645 cell_1rw
* cell instance $31342 r0 *1 160.74,147.42
X$31342 522 623 523 644 645 cell_1rw
* cell instance $31343 r0 *1 160.74,150.15
X$31343 522 625 523 644 645 cell_1rw
* cell instance $31344 m0 *1 160.74,152.88
X$31344 522 626 523 644 645 cell_1rw
* cell instance $31345 r0 *1 160.74,152.88
X$31345 522 627 523 644 645 cell_1rw
* cell instance $31346 m0 *1 160.74,155.61
X$31346 522 628 523 644 645 cell_1rw
* cell instance $31347 r0 *1 160.74,155.61
X$31347 522 629 523 644 645 cell_1rw
* cell instance $31348 m0 *1 160.74,158.34
X$31348 522 630 523 644 645 cell_1rw
* cell instance $31349 r0 *1 160.74,158.34
X$31349 522 631 523 644 645 cell_1rw
* cell instance $31350 m0 *1 160.74,161.07
X$31350 522 632 523 644 645 cell_1rw
* cell instance $31351 r0 *1 160.74,161.07
X$31351 522 633 523 644 645 cell_1rw
* cell instance $31352 m0 *1 160.74,163.8
X$31352 522 634 523 644 645 cell_1rw
* cell instance $31353 r0 *1 160.74,163.8
X$31353 522 635 523 644 645 cell_1rw
* cell instance $31354 m0 *1 160.74,166.53
X$31354 522 637 523 644 645 cell_1rw
* cell instance $31355 r0 *1 160.74,166.53
X$31355 522 636 523 644 645 cell_1rw
* cell instance $31356 m0 *1 160.74,169.26
X$31356 522 639 523 644 645 cell_1rw
* cell instance $31357 r0 *1 160.74,169.26
X$31357 522 638 523 644 645 cell_1rw
* cell instance $31358 m0 *1 160.74,171.99
X$31358 522 640 523 644 645 cell_1rw
* cell instance $31359 m0 *1 160.74,174.72
X$31359 522 642 523 644 645 cell_1rw
* cell instance $31360 r0 *1 160.74,171.99
X$31360 522 641 523 644 645 cell_1rw
* cell instance $31361 r0 *1 160.74,174.72
X$31361 522 643 523 644 645 cell_1rw
* cell instance $31362 m0 *1 161.445,90.09
X$31362 524 581 525 644 645 cell_1rw
* cell instance $31363 r0 *1 161.445,90.09
X$31363 524 580 525 644 645 cell_1rw
* cell instance $31364 m0 *1 161.445,92.82
X$31364 524 583 525 644 645 cell_1rw
* cell instance $31365 r0 *1 161.445,92.82
X$31365 524 582 525 644 645 cell_1rw
* cell instance $31366 m0 *1 161.445,95.55
X$31366 524 584 525 644 645 cell_1rw
* cell instance $31367 r0 *1 161.445,95.55
X$31367 524 585 525 644 645 cell_1rw
* cell instance $31368 m0 *1 161.445,98.28
X$31368 524 586 525 644 645 cell_1rw
* cell instance $31369 r0 *1 161.445,98.28
X$31369 524 587 525 644 645 cell_1rw
* cell instance $31370 m0 *1 161.445,101.01
X$31370 524 588 525 644 645 cell_1rw
* cell instance $31371 m0 *1 161.445,103.74
X$31371 524 590 525 644 645 cell_1rw
* cell instance $31372 r0 *1 161.445,101.01
X$31372 524 589 525 644 645 cell_1rw
* cell instance $31373 r0 *1 161.445,103.74
X$31373 524 591 525 644 645 cell_1rw
* cell instance $31374 m0 *1 161.445,106.47
X$31374 524 593 525 644 645 cell_1rw
* cell instance $31375 r0 *1 161.445,106.47
X$31375 524 592 525 644 645 cell_1rw
* cell instance $31376 m0 *1 161.445,109.2
X$31376 524 594 525 644 645 cell_1rw
* cell instance $31377 r0 *1 161.445,109.2
X$31377 524 595 525 644 645 cell_1rw
* cell instance $31378 m0 *1 161.445,111.93
X$31378 524 597 525 644 645 cell_1rw
* cell instance $31379 r0 *1 161.445,111.93
X$31379 524 596 525 644 645 cell_1rw
* cell instance $31380 m0 *1 161.445,114.66
X$31380 524 598 525 644 645 cell_1rw
* cell instance $31381 r0 *1 161.445,114.66
X$31381 524 599 525 644 645 cell_1rw
* cell instance $31382 m0 *1 161.445,117.39
X$31382 524 600 525 644 645 cell_1rw
* cell instance $31383 r0 *1 161.445,117.39
X$31383 524 601 525 644 645 cell_1rw
* cell instance $31384 m0 *1 161.445,120.12
X$31384 524 602 525 644 645 cell_1rw
* cell instance $31385 r0 *1 161.445,120.12
X$31385 524 603 525 644 645 cell_1rw
* cell instance $31386 m0 *1 161.445,122.85
X$31386 524 604 525 644 645 cell_1rw
* cell instance $31387 r0 *1 161.445,122.85
X$31387 524 605 525 644 645 cell_1rw
* cell instance $31388 m0 *1 161.445,125.58
X$31388 524 606 525 644 645 cell_1rw
* cell instance $31389 m0 *1 161.445,128.31
X$31389 524 609 525 644 645 cell_1rw
* cell instance $31390 r0 *1 161.445,125.58
X$31390 524 607 525 644 645 cell_1rw
* cell instance $31391 r0 *1 161.445,128.31
X$31391 524 608 525 644 645 cell_1rw
* cell instance $31392 m0 *1 161.445,131.04
X$31392 524 610 525 644 645 cell_1rw
* cell instance $31393 r0 *1 161.445,131.04
X$31393 524 611 525 644 645 cell_1rw
* cell instance $31394 m0 *1 161.445,133.77
X$31394 524 612 525 644 645 cell_1rw
* cell instance $31395 r0 *1 161.445,133.77
X$31395 524 613 525 644 645 cell_1rw
* cell instance $31396 m0 *1 161.445,136.5
X$31396 524 615 525 644 645 cell_1rw
* cell instance $31397 r0 *1 161.445,136.5
X$31397 524 614 525 644 645 cell_1rw
* cell instance $31398 m0 *1 161.445,139.23
X$31398 524 617 525 644 645 cell_1rw
* cell instance $31399 m0 *1 161.445,141.96
X$31399 524 618 525 644 645 cell_1rw
* cell instance $31400 r0 *1 161.445,139.23
X$31400 524 616 525 644 645 cell_1rw
* cell instance $31401 r0 *1 161.445,141.96
X$31401 524 619 525 644 645 cell_1rw
* cell instance $31402 m0 *1 161.445,144.69
X$31402 524 620 525 644 645 cell_1rw
* cell instance $31403 m0 *1 161.445,147.42
X$31403 524 622 525 644 645 cell_1rw
* cell instance $31404 r0 *1 161.445,144.69
X$31404 524 621 525 644 645 cell_1rw
* cell instance $31405 r0 *1 161.445,147.42
X$31405 524 623 525 644 645 cell_1rw
* cell instance $31406 m0 *1 161.445,150.15
X$31406 524 624 525 644 645 cell_1rw
* cell instance $31407 r0 *1 161.445,150.15
X$31407 524 625 525 644 645 cell_1rw
* cell instance $31408 m0 *1 161.445,152.88
X$31408 524 626 525 644 645 cell_1rw
* cell instance $31409 r0 *1 161.445,152.88
X$31409 524 627 525 644 645 cell_1rw
* cell instance $31410 m0 *1 161.445,155.61
X$31410 524 628 525 644 645 cell_1rw
* cell instance $31411 r0 *1 161.445,155.61
X$31411 524 629 525 644 645 cell_1rw
* cell instance $31412 m0 *1 161.445,158.34
X$31412 524 630 525 644 645 cell_1rw
* cell instance $31413 m0 *1 161.445,161.07
X$31413 524 632 525 644 645 cell_1rw
* cell instance $31414 r0 *1 161.445,158.34
X$31414 524 631 525 644 645 cell_1rw
* cell instance $31415 r0 *1 161.445,161.07
X$31415 524 633 525 644 645 cell_1rw
* cell instance $31416 m0 *1 161.445,163.8
X$31416 524 634 525 644 645 cell_1rw
* cell instance $31417 r0 *1 161.445,163.8
X$31417 524 635 525 644 645 cell_1rw
* cell instance $31418 m0 *1 161.445,166.53
X$31418 524 637 525 644 645 cell_1rw
* cell instance $31419 r0 *1 161.445,166.53
X$31419 524 636 525 644 645 cell_1rw
* cell instance $31420 m0 *1 161.445,169.26
X$31420 524 639 525 644 645 cell_1rw
* cell instance $31421 r0 *1 161.445,169.26
X$31421 524 638 525 644 645 cell_1rw
* cell instance $31422 m0 *1 161.445,171.99
X$31422 524 640 525 644 645 cell_1rw
* cell instance $31423 r0 *1 161.445,171.99
X$31423 524 641 525 644 645 cell_1rw
* cell instance $31424 m0 *1 161.445,174.72
X$31424 524 642 525 644 645 cell_1rw
* cell instance $31425 r0 *1 161.445,174.72
X$31425 524 643 525 644 645 cell_1rw
* cell instance $31426 m0 *1 162.15,90.09
X$31426 526 581 527 644 645 cell_1rw
* cell instance $31427 r0 *1 162.15,90.09
X$31427 526 580 527 644 645 cell_1rw
* cell instance $31428 m0 *1 162.15,92.82
X$31428 526 583 527 644 645 cell_1rw
* cell instance $31429 r0 *1 162.15,92.82
X$31429 526 582 527 644 645 cell_1rw
* cell instance $31430 m0 *1 162.15,95.55
X$31430 526 584 527 644 645 cell_1rw
* cell instance $31431 r0 *1 162.15,95.55
X$31431 526 585 527 644 645 cell_1rw
* cell instance $31432 m0 *1 162.15,98.28
X$31432 526 586 527 644 645 cell_1rw
* cell instance $31433 m0 *1 162.15,101.01
X$31433 526 588 527 644 645 cell_1rw
* cell instance $31434 r0 *1 162.15,98.28
X$31434 526 587 527 644 645 cell_1rw
* cell instance $31435 r0 *1 162.15,101.01
X$31435 526 589 527 644 645 cell_1rw
* cell instance $31436 m0 *1 162.15,103.74
X$31436 526 590 527 644 645 cell_1rw
* cell instance $31437 r0 *1 162.15,103.74
X$31437 526 591 527 644 645 cell_1rw
* cell instance $31438 m0 *1 162.15,106.47
X$31438 526 593 527 644 645 cell_1rw
* cell instance $31439 r0 *1 162.15,106.47
X$31439 526 592 527 644 645 cell_1rw
* cell instance $31440 m0 *1 162.15,109.2
X$31440 526 594 527 644 645 cell_1rw
* cell instance $31441 r0 *1 162.15,109.2
X$31441 526 595 527 644 645 cell_1rw
* cell instance $31442 m0 *1 162.15,111.93
X$31442 526 597 527 644 645 cell_1rw
* cell instance $31443 r0 *1 162.15,111.93
X$31443 526 596 527 644 645 cell_1rw
* cell instance $31444 m0 *1 162.15,114.66
X$31444 526 598 527 644 645 cell_1rw
* cell instance $31445 r0 *1 162.15,114.66
X$31445 526 599 527 644 645 cell_1rw
* cell instance $31446 m0 *1 162.15,117.39
X$31446 526 600 527 644 645 cell_1rw
* cell instance $31447 r0 *1 162.15,117.39
X$31447 526 601 527 644 645 cell_1rw
* cell instance $31448 m0 *1 162.15,120.12
X$31448 526 602 527 644 645 cell_1rw
* cell instance $31449 r0 *1 162.15,120.12
X$31449 526 603 527 644 645 cell_1rw
* cell instance $31450 m0 *1 162.15,122.85
X$31450 526 604 527 644 645 cell_1rw
* cell instance $31451 r0 *1 162.15,122.85
X$31451 526 605 527 644 645 cell_1rw
* cell instance $31452 m0 *1 162.15,125.58
X$31452 526 606 527 644 645 cell_1rw
* cell instance $31453 r0 *1 162.15,125.58
X$31453 526 607 527 644 645 cell_1rw
* cell instance $31454 m0 *1 162.15,128.31
X$31454 526 609 527 644 645 cell_1rw
* cell instance $31455 r0 *1 162.15,128.31
X$31455 526 608 527 644 645 cell_1rw
* cell instance $31456 m0 *1 162.15,131.04
X$31456 526 610 527 644 645 cell_1rw
* cell instance $31457 r0 *1 162.15,131.04
X$31457 526 611 527 644 645 cell_1rw
* cell instance $31458 m0 *1 162.15,133.77
X$31458 526 612 527 644 645 cell_1rw
* cell instance $31459 r0 *1 162.15,133.77
X$31459 526 613 527 644 645 cell_1rw
* cell instance $31460 m0 *1 162.15,136.5
X$31460 526 615 527 644 645 cell_1rw
* cell instance $31461 m0 *1 162.15,139.23
X$31461 526 617 527 644 645 cell_1rw
* cell instance $31462 r0 *1 162.15,136.5
X$31462 526 614 527 644 645 cell_1rw
* cell instance $31463 r0 *1 162.15,139.23
X$31463 526 616 527 644 645 cell_1rw
* cell instance $31464 m0 *1 162.15,141.96
X$31464 526 618 527 644 645 cell_1rw
* cell instance $31465 r0 *1 162.15,141.96
X$31465 526 619 527 644 645 cell_1rw
* cell instance $31466 m0 *1 162.15,144.69
X$31466 526 620 527 644 645 cell_1rw
* cell instance $31467 r0 *1 162.15,144.69
X$31467 526 621 527 644 645 cell_1rw
* cell instance $31468 m0 *1 162.15,147.42
X$31468 526 622 527 644 645 cell_1rw
* cell instance $31469 m0 *1 162.15,150.15
X$31469 526 624 527 644 645 cell_1rw
* cell instance $31470 r0 *1 162.15,147.42
X$31470 526 623 527 644 645 cell_1rw
* cell instance $31471 r0 *1 162.15,150.15
X$31471 526 625 527 644 645 cell_1rw
* cell instance $31472 m0 *1 162.15,152.88
X$31472 526 626 527 644 645 cell_1rw
* cell instance $31473 m0 *1 162.15,155.61
X$31473 526 628 527 644 645 cell_1rw
* cell instance $31474 r0 *1 162.15,152.88
X$31474 526 627 527 644 645 cell_1rw
* cell instance $31475 r0 *1 162.15,155.61
X$31475 526 629 527 644 645 cell_1rw
* cell instance $31476 m0 *1 162.15,158.34
X$31476 526 630 527 644 645 cell_1rw
* cell instance $31477 m0 *1 162.15,161.07
X$31477 526 632 527 644 645 cell_1rw
* cell instance $31478 r0 *1 162.15,158.34
X$31478 526 631 527 644 645 cell_1rw
* cell instance $31479 r0 *1 162.15,161.07
X$31479 526 633 527 644 645 cell_1rw
* cell instance $31480 m0 *1 162.15,163.8
X$31480 526 634 527 644 645 cell_1rw
* cell instance $31481 m0 *1 162.15,166.53
X$31481 526 637 527 644 645 cell_1rw
* cell instance $31482 r0 *1 162.15,163.8
X$31482 526 635 527 644 645 cell_1rw
* cell instance $31483 r0 *1 162.15,166.53
X$31483 526 636 527 644 645 cell_1rw
* cell instance $31484 m0 *1 162.15,169.26
X$31484 526 639 527 644 645 cell_1rw
* cell instance $31485 r0 *1 162.15,169.26
X$31485 526 638 527 644 645 cell_1rw
* cell instance $31486 m0 *1 162.15,171.99
X$31486 526 640 527 644 645 cell_1rw
* cell instance $31487 r0 *1 162.15,171.99
X$31487 526 641 527 644 645 cell_1rw
* cell instance $31488 m0 *1 162.15,174.72
X$31488 526 642 527 644 645 cell_1rw
* cell instance $31489 r0 *1 162.15,174.72
X$31489 526 643 527 644 645 cell_1rw
* cell instance $31490 m0 *1 162.855,90.09
X$31490 528 581 529 644 645 cell_1rw
* cell instance $31491 r0 *1 162.855,90.09
X$31491 528 580 529 644 645 cell_1rw
* cell instance $31492 m0 *1 162.855,92.82
X$31492 528 583 529 644 645 cell_1rw
* cell instance $31493 r0 *1 162.855,92.82
X$31493 528 582 529 644 645 cell_1rw
* cell instance $31494 m0 *1 162.855,95.55
X$31494 528 584 529 644 645 cell_1rw
* cell instance $31495 r0 *1 162.855,95.55
X$31495 528 585 529 644 645 cell_1rw
* cell instance $31496 m0 *1 162.855,98.28
X$31496 528 586 529 644 645 cell_1rw
* cell instance $31497 r0 *1 162.855,98.28
X$31497 528 587 529 644 645 cell_1rw
* cell instance $31498 m0 *1 162.855,101.01
X$31498 528 588 529 644 645 cell_1rw
* cell instance $31499 r0 *1 162.855,101.01
X$31499 528 589 529 644 645 cell_1rw
* cell instance $31500 m0 *1 162.855,103.74
X$31500 528 590 529 644 645 cell_1rw
* cell instance $31501 r0 *1 162.855,103.74
X$31501 528 591 529 644 645 cell_1rw
* cell instance $31502 m0 *1 162.855,106.47
X$31502 528 593 529 644 645 cell_1rw
* cell instance $31503 m0 *1 162.855,109.2
X$31503 528 594 529 644 645 cell_1rw
* cell instance $31504 r0 *1 162.855,106.47
X$31504 528 592 529 644 645 cell_1rw
* cell instance $31505 r0 *1 162.855,109.2
X$31505 528 595 529 644 645 cell_1rw
* cell instance $31506 m0 *1 162.855,111.93
X$31506 528 597 529 644 645 cell_1rw
* cell instance $31507 m0 *1 162.855,114.66
X$31507 528 598 529 644 645 cell_1rw
* cell instance $31508 r0 *1 162.855,111.93
X$31508 528 596 529 644 645 cell_1rw
* cell instance $31509 r0 *1 162.855,114.66
X$31509 528 599 529 644 645 cell_1rw
* cell instance $31510 m0 *1 162.855,117.39
X$31510 528 600 529 644 645 cell_1rw
* cell instance $31511 r0 *1 162.855,117.39
X$31511 528 601 529 644 645 cell_1rw
* cell instance $31512 m0 *1 162.855,120.12
X$31512 528 602 529 644 645 cell_1rw
* cell instance $31513 r0 *1 162.855,120.12
X$31513 528 603 529 644 645 cell_1rw
* cell instance $31514 m0 *1 162.855,122.85
X$31514 528 604 529 644 645 cell_1rw
* cell instance $31515 r0 *1 162.855,122.85
X$31515 528 605 529 644 645 cell_1rw
* cell instance $31516 m0 *1 162.855,125.58
X$31516 528 606 529 644 645 cell_1rw
* cell instance $31517 r0 *1 162.855,125.58
X$31517 528 607 529 644 645 cell_1rw
* cell instance $31518 m0 *1 162.855,128.31
X$31518 528 609 529 644 645 cell_1rw
* cell instance $31519 r0 *1 162.855,128.31
X$31519 528 608 529 644 645 cell_1rw
* cell instance $31520 m0 *1 162.855,131.04
X$31520 528 610 529 644 645 cell_1rw
* cell instance $31521 r0 *1 162.855,131.04
X$31521 528 611 529 644 645 cell_1rw
* cell instance $31522 m0 *1 162.855,133.77
X$31522 528 612 529 644 645 cell_1rw
* cell instance $31523 r0 *1 162.855,133.77
X$31523 528 613 529 644 645 cell_1rw
* cell instance $31524 m0 *1 162.855,136.5
X$31524 528 615 529 644 645 cell_1rw
* cell instance $31525 m0 *1 162.855,139.23
X$31525 528 617 529 644 645 cell_1rw
* cell instance $31526 r0 *1 162.855,136.5
X$31526 528 614 529 644 645 cell_1rw
* cell instance $31527 r0 *1 162.855,139.23
X$31527 528 616 529 644 645 cell_1rw
* cell instance $31528 m0 *1 162.855,141.96
X$31528 528 618 529 644 645 cell_1rw
* cell instance $31529 r0 *1 162.855,141.96
X$31529 528 619 529 644 645 cell_1rw
* cell instance $31530 m0 *1 162.855,144.69
X$31530 528 620 529 644 645 cell_1rw
* cell instance $31531 r0 *1 162.855,144.69
X$31531 528 621 529 644 645 cell_1rw
* cell instance $31532 m0 *1 162.855,147.42
X$31532 528 622 529 644 645 cell_1rw
* cell instance $31533 r0 *1 162.855,147.42
X$31533 528 623 529 644 645 cell_1rw
* cell instance $31534 m0 *1 162.855,150.15
X$31534 528 624 529 644 645 cell_1rw
* cell instance $31535 r0 *1 162.855,150.15
X$31535 528 625 529 644 645 cell_1rw
* cell instance $31536 m0 *1 162.855,152.88
X$31536 528 626 529 644 645 cell_1rw
* cell instance $31537 m0 *1 162.855,155.61
X$31537 528 628 529 644 645 cell_1rw
* cell instance $31538 r0 *1 162.855,152.88
X$31538 528 627 529 644 645 cell_1rw
* cell instance $31539 r0 *1 162.855,155.61
X$31539 528 629 529 644 645 cell_1rw
* cell instance $31540 m0 *1 162.855,158.34
X$31540 528 630 529 644 645 cell_1rw
* cell instance $31541 r0 *1 162.855,158.34
X$31541 528 631 529 644 645 cell_1rw
* cell instance $31542 m0 *1 162.855,161.07
X$31542 528 632 529 644 645 cell_1rw
* cell instance $31543 r0 *1 162.855,161.07
X$31543 528 633 529 644 645 cell_1rw
* cell instance $31544 m0 *1 162.855,163.8
X$31544 528 634 529 644 645 cell_1rw
* cell instance $31545 r0 *1 162.855,163.8
X$31545 528 635 529 644 645 cell_1rw
* cell instance $31546 m0 *1 162.855,166.53
X$31546 528 637 529 644 645 cell_1rw
* cell instance $31547 r0 *1 162.855,166.53
X$31547 528 636 529 644 645 cell_1rw
* cell instance $31548 m0 *1 162.855,169.26
X$31548 528 639 529 644 645 cell_1rw
* cell instance $31549 r0 *1 162.855,169.26
X$31549 528 638 529 644 645 cell_1rw
* cell instance $31550 m0 *1 162.855,171.99
X$31550 528 640 529 644 645 cell_1rw
* cell instance $31551 r0 *1 162.855,171.99
X$31551 528 641 529 644 645 cell_1rw
* cell instance $31552 m0 *1 162.855,174.72
X$31552 528 642 529 644 645 cell_1rw
* cell instance $31553 r0 *1 162.855,174.72
X$31553 528 643 529 644 645 cell_1rw
* cell instance $31554 m0 *1 163.56,90.09
X$31554 530 581 531 644 645 cell_1rw
* cell instance $31555 r0 *1 163.56,90.09
X$31555 530 580 531 644 645 cell_1rw
* cell instance $31556 m0 *1 163.56,92.82
X$31556 530 583 531 644 645 cell_1rw
* cell instance $31557 r0 *1 163.56,92.82
X$31557 530 582 531 644 645 cell_1rw
* cell instance $31558 m0 *1 163.56,95.55
X$31558 530 584 531 644 645 cell_1rw
* cell instance $31559 r0 *1 163.56,95.55
X$31559 530 585 531 644 645 cell_1rw
* cell instance $31560 m0 *1 163.56,98.28
X$31560 530 586 531 644 645 cell_1rw
* cell instance $31561 m0 *1 163.56,101.01
X$31561 530 588 531 644 645 cell_1rw
* cell instance $31562 r0 *1 163.56,98.28
X$31562 530 587 531 644 645 cell_1rw
* cell instance $31563 r0 *1 163.56,101.01
X$31563 530 589 531 644 645 cell_1rw
* cell instance $31564 m0 *1 163.56,103.74
X$31564 530 590 531 644 645 cell_1rw
* cell instance $31565 r0 *1 163.56,103.74
X$31565 530 591 531 644 645 cell_1rw
* cell instance $31566 m0 *1 163.56,106.47
X$31566 530 593 531 644 645 cell_1rw
* cell instance $31567 r0 *1 163.56,106.47
X$31567 530 592 531 644 645 cell_1rw
* cell instance $31568 m0 *1 163.56,109.2
X$31568 530 594 531 644 645 cell_1rw
* cell instance $31569 r0 *1 163.56,109.2
X$31569 530 595 531 644 645 cell_1rw
* cell instance $31570 m0 *1 163.56,111.93
X$31570 530 597 531 644 645 cell_1rw
* cell instance $31571 r0 *1 163.56,111.93
X$31571 530 596 531 644 645 cell_1rw
* cell instance $31572 m0 *1 163.56,114.66
X$31572 530 598 531 644 645 cell_1rw
* cell instance $31573 r0 *1 163.56,114.66
X$31573 530 599 531 644 645 cell_1rw
* cell instance $31574 m0 *1 163.56,117.39
X$31574 530 600 531 644 645 cell_1rw
* cell instance $31575 r0 *1 163.56,117.39
X$31575 530 601 531 644 645 cell_1rw
* cell instance $31576 m0 *1 163.56,120.12
X$31576 530 602 531 644 645 cell_1rw
* cell instance $31577 m0 *1 163.56,122.85
X$31577 530 604 531 644 645 cell_1rw
* cell instance $31578 r0 *1 163.56,120.12
X$31578 530 603 531 644 645 cell_1rw
* cell instance $31579 r0 *1 163.56,122.85
X$31579 530 605 531 644 645 cell_1rw
* cell instance $31580 m0 *1 163.56,125.58
X$31580 530 606 531 644 645 cell_1rw
* cell instance $31581 r0 *1 163.56,125.58
X$31581 530 607 531 644 645 cell_1rw
* cell instance $31582 m0 *1 163.56,128.31
X$31582 530 609 531 644 645 cell_1rw
* cell instance $31583 m0 *1 163.56,131.04
X$31583 530 610 531 644 645 cell_1rw
* cell instance $31584 r0 *1 163.56,128.31
X$31584 530 608 531 644 645 cell_1rw
* cell instance $31585 r0 *1 163.56,131.04
X$31585 530 611 531 644 645 cell_1rw
* cell instance $31586 m0 *1 163.56,133.77
X$31586 530 612 531 644 645 cell_1rw
* cell instance $31587 r0 *1 163.56,133.77
X$31587 530 613 531 644 645 cell_1rw
* cell instance $31588 m0 *1 163.56,136.5
X$31588 530 615 531 644 645 cell_1rw
* cell instance $31589 r0 *1 163.56,136.5
X$31589 530 614 531 644 645 cell_1rw
* cell instance $31590 m0 *1 163.56,139.23
X$31590 530 617 531 644 645 cell_1rw
* cell instance $31591 m0 *1 163.56,141.96
X$31591 530 618 531 644 645 cell_1rw
* cell instance $31592 r0 *1 163.56,139.23
X$31592 530 616 531 644 645 cell_1rw
* cell instance $31593 r0 *1 163.56,141.96
X$31593 530 619 531 644 645 cell_1rw
* cell instance $31594 m0 *1 163.56,144.69
X$31594 530 620 531 644 645 cell_1rw
* cell instance $31595 r0 *1 163.56,144.69
X$31595 530 621 531 644 645 cell_1rw
* cell instance $31596 m0 *1 163.56,147.42
X$31596 530 622 531 644 645 cell_1rw
* cell instance $31597 r0 *1 163.56,147.42
X$31597 530 623 531 644 645 cell_1rw
* cell instance $31598 m0 *1 163.56,150.15
X$31598 530 624 531 644 645 cell_1rw
* cell instance $31599 r0 *1 163.56,150.15
X$31599 530 625 531 644 645 cell_1rw
* cell instance $31600 m0 *1 163.56,152.88
X$31600 530 626 531 644 645 cell_1rw
* cell instance $31601 r0 *1 163.56,152.88
X$31601 530 627 531 644 645 cell_1rw
* cell instance $31602 m0 *1 163.56,155.61
X$31602 530 628 531 644 645 cell_1rw
* cell instance $31603 r0 *1 163.56,155.61
X$31603 530 629 531 644 645 cell_1rw
* cell instance $31604 m0 *1 163.56,158.34
X$31604 530 630 531 644 645 cell_1rw
* cell instance $31605 m0 *1 163.56,161.07
X$31605 530 632 531 644 645 cell_1rw
* cell instance $31606 r0 *1 163.56,158.34
X$31606 530 631 531 644 645 cell_1rw
* cell instance $31607 r0 *1 163.56,161.07
X$31607 530 633 531 644 645 cell_1rw
* cell instance $31608 m0 *1 163.56,163.8
X$31608 530 634 531 644 645 cell_1rw
* cell instance $31609 r0 *1 163.56,163.8
X$31609 530 635 531 644 645 cell_1rw
* cell instance $31610 m0 *1 163.56,166.53
X$31610 530 637 531 644 645 cell_1rw
* cell instance $31611 r0 *1 163.56,166.53
X$31611 530 636 531 644 645 cell_1rw
* cell instance $31612 m0 *1 163.56,169.26
X$31612 530 639 531 644 645 cell_1rw
* cell instance $31613 r0 *1 163.56,169.26
X$31613 530 638 531 644 645 cell_1rw
* cell instance $31614 m0 *1 163.56,171.99
X$31614 530 640 531 644 645 cell_1rw
* cell instance $31615 r0 *1 163.56,171.99
X$31615 530 641 531 644 645 cell_1rw
* cell instance $31616 m0 *1 163.56,174.72
X$31616 530 642 531 644 645 cell_1rw
* cell instance $31617 r0 *1 163.56,174.72
X$31617 530 643 531 644 645 cell_1rw
* cell instance $31618 m0 *1 164.265,90.09
X$31618 532 581 533 644 645 cell_1rw
* cell instance $31619 r0 *1 164.265,90.09
X$31619 532 580 533 644 645 cell_1rw
* cell instance $31620 m0 *1 164.265,92.82
X$31620 532 583 533 644 645 cell_1rw
* cell instance $31621 r0 *1 164.265,92.82
X$31621 532 582 533 644 645 cell_1rw
* cell instance $31622 m0 *1 164.265,95.55
X$31622 532 584 533 644 645 cell_1rw
* cell instance $31623 r0 *1 164.265,95.55
X$31623 532 585 533 644 645 cell_1rw
* cell instance $31624 m0 *1 164.265,98.28
X$31624 532 586 533 644 645 cell_1rw
* cell instance $31625 r0 *1 164.265,98.28
X$31625 532 587 533 644 645 cell_1rw
* cell instance $31626 m0 *1 164.265,101.01
X$31626 532 588 533 644 645 cell_1rw
* cell instance $31627 r0 *1 164.265,101.01
X$31627 532 589 533 644 645 cell_1rw
* cell instance $31628 m0 *1 164.265,103.74
X$31628 532 590 533 644 645 cell_1rw
* cell instance $31629 m0 *1 164.265,106.47
X$31629 532 593 533 644 645 cell_1rw
* cell instance $31630 r0 *1 164.265,103.74
X$31630 532 591 533 644 645 cell_1rw
* cell instance $31631 r0 *1 164.265,106.47
X$31631 532 592 533 644 645 cell_1rw
* cell instance $31632 m0 *1 164.265,109.2
X$31632 532 594 533 644 645 cell_1rw
* cell instance $31633 r0 *1 164.265,109.2
X$31633 532 595 533 644 645 cell_1rw
* cell instance $31634 m0 *1 164.265,111.93
X$31634 532 597 533 644 645 cell_1rw
* cell instance $31635 r0 *1 164.265,111.93
X$31635 532 596 533 644 645 cell_1rw
* cell instance $31636 m0 *1 164.265,114.66
X$31636 532 598 533 644 645 cell_1rw
* cell instance $31637 r0 *1 164.265,114.66
X$31637 532 599 533 644 645 cell_1rw
* cell instance $31638 m0 *1 164.265,117.39
X$31638 532 600 533 644 645 cell_1rw
* cell instance $31639 r0 *1 164.265,117.39
X$31639 532 601 533 644 645 cell_1rw
* cell instance $31640 m0 *1 164.265,120.12
X$31640 532 602 533 644 645 cell_1rw
* cell instance $31641 r0 *1 164.265,120.12
X$31641 532 603 533 644 645 cell_1rw
* cell instance $31642 m0 *1 164.265,122.85
X$31642 532 604 533 644 645 cell_1rw
* cell instance $31643 r0 *1 164.265,122.85
X$31643 532 605 533 644 645 cell_1rw
* cell instance $31644 m0 *1 164.265,125.58
X$31644 532 606 533 644 645 cell_1rw
* cell instance $31645 r0 *1 164.265,125.58
X$31645 532 607 533 644 645 cell_1rw
* cell instance $31646 m0 *1 164.265,128.31
X$31646 532 609 533 644 645 cell_1rw
* cell instance $31647 r0 *1 164.265,128.31
X$31647 532 608 533 644 645 cell_1rw
* cell instance $31648 m0 *1 164.265,131.04
X$31648 532 610 533 644 645 cell_1rw
* cell instance $31649 r0 *1 164.265,131.04
X$31649 532 611 533 644 645 cell_1rw
* cell instance $31650 m0 *1 164.265,133.77
X$31650 532 612 533 644 645 cell_1rw
* cell instance $31651 m0 *1 164.265,136.5
X$31651 532 615 533 644 645 cell_1rw
* cell instance $31652 r0 *1 164.265,133.77
X$31652 532 613 533 644 645 cell_1rw
* cell instance $31653 m0 *1 164.265,139.23
X$31653 532 617 533 644 645 cell_1rw
* cell instance $31654 r0 *1 164.265,136.5
X$31654 532 614 533 644 645 cell_1rw
* cell instance $31655 r0 *1 164.265,139.23
X$31655 532 616 533 644 645 cell_1rw
* cell instance $31656 m0 *1 164.265,141.96
X$31656 532 618 533 644 645 cell_1rw
* cell instance $31657 r0 *1 164.265,141.96
X$31657 532 619 533 644 645 cell_1rw
* cell instance $31658 m0 *1 164.265,144.69
X$31658 532 620 533 644 645 cell_1rw
* cell instance $31659 m0 *1 164.265,147.42
X$31659 532 622 533 644 645 cell_1rw
* cell instance $31660 r0 *1 164.265,144.69
X$31660 532 621 533 644 645 cell_1rw
* cell instance $31661 m0 *1 164.265,150.15
X$31661 532 624 533 644 645 cell_1rw
* cell instance $31662 r0 *1 164.265,147.42
X$31662 532 623 533 644 645 cell_1rw
* cell instance $31663 r0 *1 164.265,150.15
X$31663 532 625 533 644 645 cell_1rw
* cell instance $31664 m0 *1 164.265,152.88
X$31664 532 626 533 644 645 cell_1rw
* cell instance $31665 r0 *1 164.265,152.88
X$31665 532 627 533 644 645 cell_1rw
* cell instance $31666 m0 *1 164.265,155.61
X$31666 532 628 533 644 645 cell_1rw
* cell instance $31667 m0 *1 164.265,158.34
X$31667 532 630 533 644 645 cell_1rw
* cell instance $31668 r0 *1 164.265,155.61
X$31668 532 629 533 644 645 cell_1rw
* cell instance $31669 r0 *1 164.265,158.34
X$31669 532 631 533 644 645 cell_1rw
* cell instance $31670 m0 *1 164.265,161.07
X$31670 532 632 533 644 645 cell_1rw
* cell instance $31671 r0 *1 164.265,161.07
X$31671 532 633 533 644 645 cell_1rw
* cell instance $31672 m0 *1 164.265,163.8
X$31672 532 634 533 644 645 cell_1rw
* cell instance $31673 r0 *1 164.265,163.8
X$31673 532 635 533 644 645 cell_1rw
* cell instance $31674 m0 *1 164.265,166.53
X$31674 532 637 533 644 645 cell_1rw
* cell instance $31675 r0 *1 164.265,166.53
X$31675 532 636 533 644 645 cell_1rw
* cell instance $31676 m0 *1 164.265,169.26
X$31676 532 639 533 644 645 cell_1rw
* cell instance $31677 r0 *1 164.265,169.26
X$31677 532 638 533 644 645 cell_1rw
* cell instance $31678 m0 *1 164.265,171.99
X$31678 532 640 533 644 645 cell_1rw
* cell instance $31679 m0 *1 164.265,174.72
X$31679 532 642 533 644 645 cell_1rw
* cell instance $31680 r0 *1 164.265,171.99
X$31680 532 641 533 644 645 cell_1rw
* cell instance $31681 r0 *1 164.265,174.72
X$31681 532 643 533 644 645 cell_1rw
* cell instance $31682 m0 *1 164.97,90.09
X$31682 534 581 535 644 645 cell_1rw
* cell instance $31683 r0 *1 164.97,90.09
X$31683 534 580 535 644 645 cell_1rw
* cell instance $31684 m0 *1 164.97,92.82
X$31684 534 583 535 644 645 cell_1rw
* cell instance $31685 r0 *1 164.97,92.82
X$31685 534 582 535 644 645 cell_1rw
* cell instance $31686 m0 *1 164.97,95.55
X$31686 534 584 535 644 645 cell_1rw
* cell instance $31687 r0 *1 164.97,95.55
X$31687 534 585 535 644 645 cell_1rw
* cell instance $31688 m0 *1 164.97,98.28
X$31688 534 586 535 644 645 cell_1rw
* cell instance $31689 r0 *1 164.97,98.28
X$31689 534 587 535 644 645 cell_1rw
* cell instance $31690 m0 *1 164.97,101.01
X$31690 534 588 535 644 645 cell_1rw
* cell instance $31691 r0 *1 164.97,101.01
X$31691 534 589 535 644 645 cell_1rw
* cell instance $31692 m0 *1 164.97,103.74
X$31692 534 590 535 644 645 cell_1rw
* cell instance $31693 r0 *1 164.97,103.74
X$31693 534 591 535 644 645 cell_1rw
* cell instance $31694 m0 *1 164.97,106.47
X$31694 534 593 535 644 645 cell_1rw
* cell instance $31695 r0 *1 164.97,106.47
X$31695 534 592 535 644 645 cell_1rw
* cell instance $31696 m0 *1 164.97,109.2
X$31696 534 594 535 644 645 cell_1rw
* cell instance $31697 m0 *1 164.97,111.93
X$31697 534 597 535 644 645 cell_1rw
* cell instance $31698 r0 *1 164.97,109.2
X$31698 534 595 535 644 645 cell_1rw
* cell instance $31699 r0 *1 164.97,111.93
X$31699 534 596 535 644 645 cell_1rw
* cell instance $31700 m0 *1 164.97,114.66
X$31700 534 598 535 644 645 cell_1rw
* cell instance $31701 r0 *1 164.97,114.66
X$31701 534 599 535 644 645 cell_1rw
* cell instance $31702 m0 *1 164.97,117.39
X$31702 534 600 535 644 645 cell_1rw
* cell instance $31703 r0 *1 164.97,117.39
X$31703 534 601 535 644 645 cell_1rw
* cell instance $31704 m0 *1 164.97,120.12
X$31704 534 602 535 644 645 cell_1rw
* cell instance $31705 r0 *1 164.97,120.12
X$31705 534 603 535 644 645 cell_1rw
* cell instance $31706 m0 *1 164.97,122.85
X$31706 534 604 535 644 645 cell_1rw
* cell instance $31707 m0 *1 164.97,125.58
X$31707 534 606 535 644 645 cell_1rw
* cell instance $31708 r0 *1 164.97,122.85
X$31708 534 605 535 644 645 cell_1rw
* cell instance $31709 r0 *1 164.97,125.58
X$31709 534 607 535 644 645 cell_1rw
* cell instance $31710 m0 *1 164.97,128.31
X$31710 534 609 535 644 645 cell_1rw
* cell instance $31711 r0 *1 164.97,128.31
X$31711 534 608 535 644 645 cell_1rw
* cell instance $31712 m0 *1 164.97,131.04
X$31712 534 610 535 644 645 cell_1rw
* cell instance $31713 r0 *1 164.97,131.04
X$31713 534 611 535 644 645 cell_1rw
* cell instance $31714 m0 *1 164.97,133.77
X$31714 534 612 535 644 645 cell_1rw
* cell instance $31715 r0 *1 164.97,133.77
X$31715 534 613 535 644 645 cell_1rw
* cell instance $31716 m0 *1 164.97,136.5
X$31716 534 615 535 644 645 cell_1rw
* cell instance $31717 r0 *1 164.97,136.5
X$31717 534 614 535 644 645 cell_1rw
* cell instance $31718 m0 *1 164.97,139.23
X$31718 534 617 535 644 645 cell_1rw
* cell instance $31719 r0 *1 164.97,139.23
X$31719 534 616 535 644 645 cell_1rw
* cell instance $31720 m0 *1 164.97,141.96
X$31720 534 618 535 644 645 cell_1rw
* cell instance $31721 m0 *1 164.97,144.69
X$31721 534 620 535 644 645 cell_1rw
* cell instance $31722 r0 *1 164.97,141.96
X$31722 534 619 535 644 645 cell_1rw
* cell instance $31723 m0 *1 164.97,147.42
X$31723 534 622 535 644 645 cell_1rw
* cell instance $31724 r0 *1 164.97,144.69
X$31724 534 621 535 644 645 cell_1rw
* cell instance $31725 r0 *1 164.97,147.42
X$31725 534 623 535 644 645 cell_1rw
* cell instance $31726 m0 *1 164.97,150.15
X$31726 534 624 535 644 645 cell_1rw
* cell instance $31727 r0 *1 164.97,150.15
X$31727 534 625 535 644 645 cell_1rw
* cell instance $31728 m0 *1 164.97,152.88
X$31728 534 626 535 644 645 cell_1rw
* cell instance $31729 r0 *1 164.97,152.88
X$31729 534 627 535 644 645 cell_1rw
* cell instance $31730 m0 *1 164.97,155.61
X$31730 534 628 535 644 645 cell_1rw
* cell instance $31731 r0 *1 164.97,155.61
X$31731 534 629 535 644 645 cell_1rw
* cell instance $31732 m0 *1 164.97,158.34
X$31732 534 630 535 644 645 cell_1rw
* cell instance $31733 r0 *1 164.97,158.34
X$31733 534 631 535 644 645 cell_1rw
* cell instance $31734 m0 *1 164.97,161.07
X$31734 534 632 535 644 645 cell_1rw
* cell instance $31735 r0 *1 164.97,161.07
X$31735 534 633 535 644 645 cell_1rw
* cell instance $31736 m0 *1 164.97,163.8
X$31736 534 634 535 644 645 cell_1rw
* cell instance $31737 m0 *1 164.97,166.53
X$31737 534 637 535 644 645 cell_1rw
* cell instance $31738 r0 *1 164.97,163.8
X$31738 534 635 535 644 645 cell_1rw
* cell instance $31739 r0 *1 164.97,166.53
X$31739 534 636 535 644 645 cell_1rw
* cell instance $31740 m0 *1 164.97,169.26
X$31740 534 639 535 644 645 cell_1rw
* cell instance $31741 r0 *1 164.97,169.26
X$31741 534 638 535 644 645 cell_1rw
* cell instance $31742 m0 *1 164.97,171.99
X$31742 534 640 535 644 645 cell_1rw
* cell instance $31743 r0 *1 164.97,171.99
X$31743 534 641 535 644 645 cell_1rw
* cell instance $31744 m0 *1 164.97,174.72
X$31744 534 642 535 644 645 cell_1rw
* cell instance $31745 r0 *1 164.97,174.72
X$31745 534 643 535 644 645 cell_1rw
* cell instance $31746 m0 *1 165.675,90.09
X$31746 536 581 537 644 645 cell_1rw
* cell instance $31747 r0 *1 165.675,90.09
X$31747 536 580 537 644 645 cell_1rw
* cell instance $31748 m0 *1 165.675,92.82
X$31748 536 583 537 644 645 cell_1rw
* cell instance $31749 r0 *1 165.675,92.82
X$31749 536 582 537 644 645 cell_1rw
* cell instance $31750 m0 *1 165.675,95.55
X$31750 536 584 537 644 645 cell_1rw
* cell instance $31751 r0 *1 165.675,95.55
X$31751 536 585 537 644 645 cell_1rw
* cell instance $31752 m0 *1 165.675,98.28
X$31752 536 586 537 644 645 cell_1rw
* cell instance $31753 r0 *1 165.675,98.28
X$31753 536 587 537 644 645 cell_1rw
* cell instance $31754 m0 *1 165.675,101.01
X$31754 536 588 537 644 645 cell_1rw
* cell instance $31755 r0 *1 165.675,101.01
X$31755 536 589 537 644 645 cell_1rw
* cell instance $31756 m0 *1 165.675,103.74
X$31756 536 590 537 644 645 cell_1rw
* cell instance $31757 r0 *1 165.675,103.74
X$31757 536 591 537 644 645 cell_1rw
* cell instance $31758 m0 *1 165.675,106.47
X$31758 536 593 537 644 645 cell_1rw
* cell instance $31759 r0 *1 165.675,106.47
X$31759 536 592 537 644 645 cell_1rw
* cell instance $31760 m0 *1 165.675,109.2
X$31760 536 594 537 644 645 cell_1rw
* cell instance $31761 m0 *1 165.675,111.93
X$31761 536 597 537 644 645 cell_1rw
* cell instance $31762 r0 *1 165.675,109.2
X$31762 536 595 537 644 645 cell_1rw
* cell instance $31763 r0 *1 165.675,111.93
X$31763 536 596 537 644 645 cell_1rw
* cell instance $31764 m0 *1 165.675,114.66
X$31764 536 598 537 644 645 cell_1rw
* cell instance $31765 r0 *1 165.675,114.66
X$31765 536 599 537 644 645 cell_1rw
* cell instance $31766 m0 *1 165.675,117.39
X$31766 536 600 537 644 645 cell_1rw
* cell instance $31767 r0 *1 165.675,117.39
X$31767 536 601 537 644 645 cell_1rw
* cell instance $31768 m0 *1 165.675,120.12
X$31768 536 602 537 644 645 cell_1rw
* cell instance $31769 r0 *1 165.675,120.12
X$31769 536 603 537 644 645 cell_1rw
* cell instance $31770 m0 *1 165.675,122.85
X$31770 536 604 537 644 645 cell_1rw
* cell instance $31771 r0 *1 165.675,122.85
X$31771 536 605 537 644 645 cell_1rw
* cell instance $31772 m0 *1 165.675,125.58
X$31772 536 606 537 644 645 cell_1rw
* cell instance $31773 r0 *1 165.675,125.58
X$31773 536 607 537 644 645 cell_1rw
* cell instance $31774 m0 *1 165.675,128.31
X$31774 536 609 537 644 645 cell_1rw
* cell instance $31775 r0 *1 165.675,128.31
X$31775 536 608 537 644 645 cell_1rw
* cell instance $31776 m0 *1 165.675,131.04
X$31776 536 610 537 644 645 cell_1rw
* cell instance $31777 r0 *1 165.675,131.04
X$31777 536 611 537 644 645 cell_1rw
* cell instance $31778 m0 *1 165.675,133.77
X$31778 536 612 537 644 645 cell_1rw
* cell instance $31779 r0 *1 165.675,133.77
X$31779 536 613 537 644 645 cell_1rw
* cell instance $31780 m0 *1 165.675,136.5
X$31780 536 615 537 644 645 cell_1rw
* cell instance $31781 r0 *1 165.675,136.5
X$31781 536 614 537 644 645 cell_1rw
* cell instance $31782 m0 *1 165.675,139.23
X$31782 536 617 537 644 645 cell_1rw
* cell instance $31783 r0 *1 165.675,139.23
X$31783 536 616 537 644 645 cell_1rw
* cell instance $31784 m0 *1 165.675,141.96
X$31784 536 618 537 644 645 cell_1rw
* cell instance $31785 r0 *1 165.675,141.96
X$31785 536 619 537 644 645 cell_1rw
* cell instance $31786 m0 *1 165.675,144.69
X$31786 536 620 537 644 645 cell_1rw
* cell instance $31787 r0 *1 165.675,144.69
X$31787 536 621 537 644 645 cell_1rw
* cell instance $31788 m0 *1 165.675,147.42
X$31788 536 622 537 644 645 cell_1rw
* cell instance $31789 r0 *1 165.675,147.42
X$31789 536 623 537 644 645 cell_1rw
* cell instance $31790 m0 *1 165.675,150.15
X$31790 536 624 537 644 645 cell_1rw
* cell instance $31791 m0 *1 165.675,152.88
X$31791 536 626 537 644 645 cell_1rw
* cell instance $31792 r0 *1 165.675,150.15
X$31792 536 625 537 644 645 cell_1rw
* cell instance $31793 r0 *1 165.675,152.88
X$31793 536 627 537 644 645 cell_1rw
* cell instance $31794 m0 *1 165.675,155.61
X$31794 536 628 537 644 645 cell_1rw
* cell instance $31795 r0 *1 165.675,155.61
X$31795 536 629 537 644 645 cell_1rw
* cell instance $31796 m0 *1 165.675,158.34
X$31796 536 630 537 644 645 cell_1rw
* cell instance $31797 r0 *1 165.675,158.34
X$31797 536 631 537 644 645 cell_1rw
* cell instance $31798 m0 *1 165.675,161.07
X$31798 536 632 537 644 645 cell_1rw
* cell instance $31799 r0 *1 165.675,161.07
X$31799 536 633 537 644 645 cell_1rw
* cell instance $31800 m0 *1 165.675,163.8
X$31800 536 634 537 644 645 cell_1rw
* cell instance $31801 r0 *1 165.675,163.8
X$31801 536 635 537 644 645 cell_1rw
* cell instance $31802 m0 *1 165.675,166.53
X$31802 536 637 537 644 645 cell_1rw
* cell instance $31803 r0 *1 165.675,166.53
X$31803 536 636 537 644 645 cell_1rw
* cell instance $31804 m0 *1 165.675,169.26
X$31804 536 639 537 644 645 cell_1rw
* cell instance $31805 r0 *1 165.675,169.26
X$31805 536 638 537 644 645 cell_1rw
* cell instance $31806 m0 *1 165.675,171.99
X$31806 536 640 537 644 645 cell_1rw
* cell instance $31807 r0 *1 165.675,171.99
X$31807 536 641 537 644 645 cell_1rw
* cell instance $31808 m0 *1 165.675,174.72
X$31808 536 642 537 644 645 cell_1rw
* cell instance $31809 r0 *1 165.675,174.72
X$31809 536 643 537 644 645 cell_1rw
* cell instance $31810 m0 *1 166.38,90.09
X$31810 538 581 539 644 645 cell_1rw
* cell instance $31811 r0 *1 166.38,90.09
X$31811 538 580 539 644 645 cell_1rw
* cell instance $31812 m0 *1 166.38,92.82
X$31812 538 583 539 644 645 cell_1rw
* cell instance $31813 r0 *1 166.38,92.82
X$31813 538 582 539 644 645 cell_1rw
* cell instance $31814 m0 *1 166.38,95.55
X$31814 538 584 539 644 645 cell_1rw
* cell instance $31815 r0 *1 166.38,95.55
X$31815 538 585 539 644 645 cell_1rw
* cell instance $31816 m0 *1 166.38,98.28
X$31816 538 586 539 644 645 cell_1rw
* cell instance $31817 r0 *1 166.38,98.28
X$31817 538 587 539 644 645 cell_1rw
* cell instance $31818 m0 *1 166.38,101.01
X$31818 538 588 539 644 645 cell_1rw
* cell instance $31819 m0 *1 166.38,103.74
X$31819 538 590 539 644 645 cell_1rw
* cell instance $31820 r0 *1 166.38,101.01
X$31820 538 589 539 644 645 cell_1rw
* cell instance $31821 r0 *1 166.38,103.74
X$31821 538 591 539 644 645 cell_1rw
* cell instance $31822 m0 *1 166.38,106.47
X$31822 538 593 539 644 645 cell_1rw
* cell instance $31823 r0 *1 166.38,106.47
X$31823 538 592 539 644 645 cell_1rw
* cell instance $31824 m0 *1 166.38,109.2
X$31824 538 594 539 644 645 cell_1rw
* cell instance $31825 r0 *1 166.38,109.2
X$31825 538 595 539 644 645 cell_1rw
* cell instance $31826 m0 *1 166.38,111.93
X$31826 538 597 539 644 645 cell_1rw
* cell instance $31827 r0 *1 166.38,111.93
X$31827 538 596 539 644 645 cell_1rw
* cell instance $31828 m0 *1 166.38,114.66
X$31828 538 598 539 644 645 cell_1rw
* cell instance $31829 r0 *1 166.38,114.66
X$31829 538 599 539 644 645 cell_1rw
* cell instance $31830 m0 *1 166.38,117.39
X$31830 538 600 539 644 645 cell_1rw
* cell instance $31831 m0 *1 166.38,120.12
X$31831 538 602 539 644 645 cell_1rw
* cell instance $31832 r0 *1 166.38,117.39
X$31832 538 601 539 644 645 cell_1rw
* cell instance $31833 r0 *1 166.38,120.12
X$31833 538 603 539 644 645 cell_1rw
* cell instance $31834 m0 *1 166.38,122.85
X$31834 538 604 539 644 645 cell_1rw
* cell instance $31835 r0 *1 166.38,122.85
X$31835 538 605 539 644 645 cell_1rw
* cell instance $31836 m0 *1 166.38,125.58
X$31836 538 606 539 644 645 cell_1rw
* cell instance $31837 r0 *1 166.38,125.58
X$31837 538 607 539 644 645 cell_1rw
* cell instance $31838 m0 *1 166.38,128.31
X$31838 538 609 539 644 645 cell_1rw
* cell instance $31839 m0 *1 166.38,131.04
X$31839 538 610 539 644 645 cell_1rw
* cell instance $31840 r0 *1 166.38,128.31
X$31840 538 608 539 644 645 cell_1rw
* cell instance $31841 r0 *1 166.38,131.04
X$31841 538 611 539 644 645 cell_1rw
* cell instance $31842 m0 *1 166.38,133.77
X$31842 538 612 539 644 645 cell_1rw
* cell instance $31843 r0 *1 166.38,133.77
X$31843 538 613 539 644 645 cell_1rw
* cell instance $31844 m0 *1 166.38,136.5
X$31844 538 615 539 644 645 cell_1rw
* cell instance $31845 r0 *1 166.38,136.5
X$31845 538 614 539 644 645 cell_1rw
* cell instance $31846 m0 *1 166.38,139.23
X$31846 538 617 539 644 645 cell_1rw
* cell instance $31847 r0 *1 166.38,139.23
X$31847 538 616 539 644 645 cell_1rw
* cell instance $31848 m0 *1 166.38,141.96
X$31848 538 618 539 644 645 cell_1rw
* cell instance $31849 r0 *1 166.38,141.96
X$31849 538 619 539 644 645 cell_1rw
* cell instance $31850 m0 *1 166.38,144.69
X$31850 538 620 539 644 645 cell_1rw
* cell instance $31851 r0 *1 166.38,144.69
X$31851 538 621 539 644 645 cell_1rw
* cell instance $31852 m0 *1 166.38,147.42
X$31852 538 622 539 644 645 cell_1rw
* cell instance $31853 r0 *1 166.38,147.42
X$31853 538 623 539 644 645 cell_1rw
* cell instance $31854 m0 *1 166.38,150.15
X$31854 538 624 539 644 645 cell_1rw
* cell instance $31855 r0 *1 166.38,150.15
X$31855 538 625 539 644 645 cell_1rw
* cell instance $31856 m0 *1 166.38,152.88
X$31856 538 626 539 644 645 cell_1rw
* cell instance $31857 r0 *1 166.38,152.88
X$31857 538 627 539 644 645 cell_1rw
* cell instance $31858 m0 *1 166.38,155.61
X$31858 538 628 539 644 645 cell_1rw
* cell instance $31859 r0 *1 166.38,155.61
X$31859 538 629 539 644 645 cell_1rw
* cell instance $31860 m0 *1 166.38,158.34
X$31860 538 630 539 644 645 cell_1rw
* cell instance $31861 r0 *1 166.38,158.34
X$31861 538 631 539 644 645 cell_1rw
* cell instance $31862 m0 *1 166.38,161.07
X$31862 538 632 539 644 645 cell_1rw
* cell instance $31863 r0 *1 166.38,161.07
X$31863 538 633 539 644 645 cell_1rw
* cell instance $31864 m0 *1 166.38,163.8
X$31864 538 634 539 644 645 cell_1rw
* cell instance $31865 r0 *1 166.38,163.8
X$31865 538 635 539 644 645 cell_1rw
* cell instance $31866 m0 *1 166.38,166.53
X$31866 538 637 539 644 645 cell_1rw
* cell instance $31867 r0 *1 166.38,166.53
X$31867 538 636 539 644 645 cell_1rw
* cell instance $31868 m0 *1 166.38,169.26
X$31868 538 639 539 644 645 cell_1rw
* cell instance $31869 r0 *1 166.38,169.26
X$31869 538 638 539 644 645 cell_1rw
* cell instance $31870 m0 *1 166.38,171.99
X$31870 538 640 539 644 645 cell_1rw
* cell instance $31871 r0 *1 166.38,171.99
X$31871 538 641 539 644 645 cell_1rw
* cell instance $31872 m0 *1 166.38,174.72
X$31872 538 642 539 644 645 cell_1rw
* cell instance $31873 r0 *1 166.38,174.72
X$31873 538 643 539 644 645 cell_1rw
* cell instance $31874 m0 *1 167.085,90.09
X$31874 540 581 541 644 645 cell_1rw
* cell instance $31875 m0 *1 167.085,92.82
X$31875 540 583 541 644 645 cell_1rw
* cell instance $31876 r0 *1 167.085,90.09
X$31876 540 580 541 644 645 cell_1rw
* cell instance $31877 m0 *1 167.085,95.55
X$31877 540 584 541 644 645 cell_1rw
* cell instance $31878 r0 *1 167.085,92.82
X$31878 540 582 541 644 645 cell_1rw
* cell instance $31879 r0 *1 167.085,95.55
X$31879 540 585 541 644 645 cell_1rw
* cell instance $31880 m0 *1 167.085,98.28
X$31880 540 586 541 644 645 cell_1rw
* cell instance $31881 m0 *1 167.085,101.01
X$31881 540 588 541 644 645 cell_1rw
* cell instance $31882 r0 *1 167.085,98.28
X$31882 540 587 541 644 645 cell_1rw
* cell instance $31883 r0 *1 167.085,101.01
X$31883 540 589 541 644 645 cell_1rw
* cell instance $31884 m0 *1 167.085,103.74
X$31884 540 590 541 644 645 cell_1rw
* cell instance $31885 r0 *1 167.085,103.74
X$31885 540 591 541 644 645 cell_1rw
* cell instance $31886 m0 *1 167.085,106.47
X$31886 540 593 541 644 645 cell_1rw
* cell instance $31887 r0 *1 167.085,106.47
X$31887 540 592 541 644 645 cell_1rw
* cell instance $31888 m0 *1 167.085,109.2
X$31888 540 594 541 644 645 cell_1rw
* cell instance $31889 r0 *1 167.085,109.2
X$31889 540 595 541 644 645 cell_1rw
* cell instance $31890 m0 *1 167.085,111.93
X$31890 540 597 541 644 645 cell_1rw
* cell instance $31891 r0 *1 167.085,111.93
X$31891 540 596 541 644 645 cell_1rw
* cell instance $31892 m0 *1 167.085,114.66
X$31892 540 598 541 644 645 cell_1rw
* cell instance $31893 r0 *1 167.085,114.66
X$31893 540 599 541 644 645 cell_1rw
* cell instance $31894 m0 *1 167.085,117.39
X$31894 540 600 541 644 645 cell_1rw
* cell instance $31895 r0 *1 167.085,117.39
X$31895 540 601 541 644 645 cell_1rw
* cell instance $31896 m0 *1 167.085,120.12
X$31896 540 602 541 644 645 cell_1rw
* cell instance $31897 r0 *1 167.085,120.12
X$31897 540 603 541 644 645 cell_1rw
* cell instance $31898 m0 *1 167.085,122.85
X$31898 540 604 541 644 645 cell_1rw
* cell instance $31899 r0 *1 167.085,122.85
X$31899 540 605 541 644 645 cell_1rw
* cell instance $31900 m0 *1 167.085,125.58
X$31900 540 606 541 644 645 cell_1rw
* cell instance $31901 r0 *1 167.085,125.58
X$31901 540 607 541 644 645 cell_1rw
* cell instance $31902 m0 *1 167.085,128.31
X$31902 540 609 541 644 645 cell_1rw
* cell instance $31903 r0 *1 167.085,128.31
X$31903 540 608 541 644 645 cell_1rw
* cell instance $31904 m0 *1 167.085,131.04
X$31904 540 610 541 644 645 cell_1rw
* cell instance $31905 m0 *1 167.085,133.77
X$31905 540 612 541 644 645 cell_1rw
* cell instance $31906 r0 *1 167.085,131.04
X$31906 540 611 541 644 645 cell_1rw
* cell instance $31907 m0 *1 167.085,136.5
X$31907 540 615 541 644 645 cell_1rw
* cell instance $31908 r0 *1 167.085,133.77
X$31908 540 613 541 644 645 cell_1rw
* cell instance $31909 r0 *1 167.085,136.5
X$31909 540 614 541 644 645 cell_1rw
* cell instance $31910 m0 *1 167.085,139.23
X$31910 540 617 541 644 645 cell_1rw
* cell instance $31911 r0 *1 167.085,139.23
X$31911 540 616 541 644 645 cell_1rw
* cell instance $31912 m0 *1 167.085,141.96
X$31912 540 618 541 644 645 cell_1rw
* cell instance $31913 m0 *1 167.085,144.69
X$31913 540 620 541 644 645 cell_1rw
* cell instance $31914 r0 *1 167.085,141.96
X$31914 540 619 541 644 645 cell_1rw
* cell instance $31915 r0 *1 167.085,144.69
X$31915 540 621 541 644 645 cell_1rw
* cell instance $31916 m0 *1 167.085,147.42
X$31916 540 622 541 644 645 cell_1rw
* cell instance $31917 r0 *1 167.085,147.42
X$31917 540 623 541 644 645 cell_1rw
* cell instance $31918 m0 *1 167.085,150.15
X$31918 540 624 541 644 645 cell_1rw
* cell instance $31919 r0 *1 167.085,150.15
X$31919 540 625 541 644 645 cell_1rw
* cell instance $31920 m0 *1 167.085,152.88
X$31920 540 626 541 644 645 cell_1rw
* cell instance $31921 r0 *1 167.085,152.88
X$31921 540 627 541 644 645 cell_1rw
* cell instance $31922 m0 *1 167.085,155.61
X$31922 540 628 541 644 645 cell_1rw
* cell instance $31923 r0 *1 167.085,155.61
X$31923 540 629 541 644 645 cell_1rw
* cell instance $31924 m0 *1 167.085,158.34
X$31924 540 630 541 644 645 cell_1rw
* cell instance $31925 r0 *1 167.085,158.34
X$31925 540 631 541 644 645 cell_1rw
* cell instance $31926 m0 *1 167.085,161.07
X$31926 540 632 541 644 645 cell_1rw
* cell instance $31927 m0 *1 167.085,163.8
X$31927 540 634 541 644 645 cell_1rw
* cell instance $31928 r0 *1 167.085,161.07
X$31928 540 633 541 644 645 cell_1rw
* cell instance $31929 m0 *1 167.085,166.53
X$31929 540 637 541 644 645 cell_1rw
* cell instance $31930 r0 *1 167.085,163.8
X$31930 540 635 541 644 645 cell_1rw
* cell instance $31931 r0 *1 167.085,166.53
X$31931 540 636 541 644 645 cell_1rw
* cell instance $31932 m0 *1 167.085,169.26
X$31932 540 639 541 644 645 cell_1rw
* cell instance $31933 r0 *1 167.085,169.26
X$31933 540 638 541 644 645 cell_1rw
* cell instance $31934 m0 *1 167.085,171.99
X$31934 540 640 541 644 645 cell_1rw
* cell instance $31935 r0 *1 167.085,171.99
X$31935 540 641 541 644 645 cell_1rw
* cell instance $31936 m0 *1 167.085,174.72
X$31936 540 642 541 644 645 cell_1rw
* cell instance $31937 r0 *1 167.085,174.72
X$31937 540 643 541 644 645 cell_1rw
* cell instance $31938 m0 *1 167.79,90.09
X$31938 542 581 543 644 645 cell_1rw
* cell instance $31939 r0 *1 167.79,90.09
X$31939 542 580 543 644 645 cell_1rw
* cell instance $31940 m0 *1 167.79,92.82
X$31940 542 583 543 644 645 cell_1rw
* cell instance $31941 m0 *1 167.79,95.55
X$31941 542 584 543 644 645 cell_1rw
* cell instance $31942 r0 *1 167.79,92.82
X$31942 542 582 543 644 645 cell_1rw
* cell instance $31943 m0 *1 167.79,98.28
X$31943 542 586 543 644 645 cell_1rw
* cell instance $31944 r0 *1 167.79,95.55
X$31944 542 585 543 644 645 cell_1rw
* cell instance $31945 r0 *1 167.79,98.28
X$31945 542 587 543 644 645 cell_1rw
* cell instance $31946 m0 *1 167.79,101.01
X$31946 542 588 543 644 645 cell_1rw
* cell instance $31947 r0 *1 167.79,101.01
X$31947 542 589 543 644 645 cell_1rw
* cell instance $31948 m0 *1 167.79,103.74
X$31948 542 590 543 644 645 cell_1rw
* cell instance $31949 m0 *1 167.79,106.47
X$31949 542 593 543 644 645 cell_1rw
* cell instance $31950 r0 *1 167.79,103.74
X$31950 542 591 543 644 645 cell_1rw
* cell instance $31951 r0 *1 167.79,106.47
X$31951 542 592 543 644 645 cell_1rw
* cell instance $31952 m0 *1 167.79,109.2
X$31952 542 594 543 644 645 cell_1rw
* cell instance $31953 r0 *1 167.79,109.2
X$31953 542 595 543 644 645 cell_1rw
* cell instance $31954 m0 *1 167.79,111.93
X$31954 542 597 543 644 645 cell_1rw
* cell instance $31955 r0 *1 167.79,111.93
X$31955 542 596 543 644 645 cell_1rw
* cell instance $31956 m0 *1 167.79,114.66
X$31956 542 598 543 644 645 cell_1rw
* cell instance $31957 r0 *1 167.79,114.66
X$31957 542 599 543 644 645 cell_1rw
* cell instance $31958 m0 *1 167.79,117.39
X$31958 542 600 543 644 645 cell_1rw
* cell instance $31959 r0 *1 167.79,117.39
X$31959 542 601 543 644 645 cell_1rw
* cell instance $31960 m0 *1 167.79,120.12
X$31960 542 602 543 644 645 cell_1rw
* cell instance $31961 r0 *1 167.79,120.12
X$31961 542 603 543 644 645 cell_1rw
* cell instance $31962 m0 *1 167.79,122.85
X$31962 542 604 543 644 645 cell_1rw
* cell instance $31963 r0 *1 167.79,122.85
X$31963 542 605 543 644 645 cell_1rw
* cell instance $31964 m0 *1 167.79,125.58
X$31964 542 606 543 644 645 cell_1rw
* cell instance $31965 m0 *1 167.79,128.31
X$31965 542 609 543 644 645 cell_1rw
* cell instance $31966 r0 *1 167.79,125.58
X$31966 542 607 543 644 645 cell_1rw
* cell instance $31967 r0 *1 167.79,128.31
X$31967 542 608 543 644 645 cell_1rw
* cell instance $31968 m0 *1 167.79,131.04
X$31968 542 610 543 644 645 cell_1rw
* cell instance $31969 m0 *1 167.79,133.77
X$31969 542 612 543 644 645 cell_1rw
* cell instance $31970 r0 *1 167.79,131.04
X$31970 542 611 543 644 645 cell_1rw
* cell instance $31971 r0 *1 167.79,133.77
X$31971 542 613 543 644 645 cell_1rw
* cell instance $31972 m0 *1 167.79,136.5
X$31972 542 615 543 644 645 cell_1rw
* cell instance $31973 r0 *1 167.79,136.5
X$31973 542 614 543 644 645 cell_1rw
* cell instance $31974 m0 *1 167.79,139.23
X$31974 542 617 543 644 645 cell_1rw
* cell instance $31975 r0 *1 167.79,139.23
X$31975 542 616 543 644 645 cell_1rw
* cell instance $31976 m0 *1 167.79,141.96
X$31976 542 618 543 644 645 cell_1rw
* cell instance $31977 r0 *1 167.79,141.96
X$31977 542 619 543 644 645 cell_1rw
* cell instance $31978 m0 *1 167.79,144.69
X$31978 542 620 543 644 645 cell_1rw
* cell instance $31979 m0 *1 167.79,147.42
X$31979 542 622 543 644 645 cell_1rw
* cell instance $31980 r0 *1 167.79,144.69
X$31980 542 621 543 644 645 cell_1rw
* cell instance $31981 r0 *1 167.79,147.42
X$31981 542 623 543 644 645 cell_1rw
* cell instance $31982 m0 *1 167.79,150.15
X$31982 542 624 543 644 645 cell_1rw
* cell instance $31983 r0 *1 167.79,150.15
X$31983 542 625 543 644 645 cell_1rw
* cell instance $31984 m0 *1 167.79,152.88
X$31984 542 626 543 644 645 cell_1rw
* cell instance $31985 r0 *1 167.79,152.88
X$31985 542 627 543 644 645 cell_1rw
* cell instance $31986 m0 *1 167.79,155.61
X$31986 542 628 543 644 645 cell_1rw
* cell instance $31987 r0 *1 167.79,155.61
X$31987 542 629 543 644 645 cell_1rw
* cell instance $31988 m0 *1 167.79,158.34
X$31988 542 630 543 644 645 cell_1rw
* cell instance $31989 m0 *1 167.79,161.07
X$31989 542 632 543 644 645 cell_1rw
* cell instance $31990 r0 *1 167.79,158.34
X$31990 542 631 543 644 645 cell_1rw
* cell instance $31991 r0 *1 167.79,161.07
X$31991 542 633 543 644 645 cell_1rw
* cell instance $31992 m0 *1 167.79,163.8
X$31992 542 634 543 644 645 cell_1rw
* cell instance $31993 r0 *1 167.79,163.8
X$31993 542 635 543 644 645 cell_1rw
* cell instance $31994 m0 *1 167.79,166.53
X$31994 542 637 543 644 645 cell_1rw
* cell instance $31995 r0 *1 167.79,166.53
X$31995 542 636 543 644 645 cell_1rw
* cell instance $31996 m0 *1 167.79,169.26
X$31996 542 639 543 644 645 cell_1rw
* cell instance $31997 r0 *1 167.79,169.26
X$31997 542 638 543 644 645 cell_1rw
* cell instance $31998 m0 *1 167.79,171.99
X$31998 542 640 543 644 645 cell_1rw
* cell instance $31999 m0 *1 167.79,174.72
X$31999 542 642 543 644 645 cell_1rw
* cell instance $32000 r0 *1 167.79,171.99
X$32000 542 641 543 644 645 cell_1rw
* cell instance $32001 r0 *1 167.79,174.72
X$32001 542 643 543 644 645 cell_1rw
* cell instance $32002 m0 *1 168.495,90.09
X$32002 544 581 545 644 645 cell_1rw
* cell instance $32003 r0 *1 168.495,90.09
X$32003 544 580 545 644 645 cell_1rw
* cell instance $32004 m0 *1 168.495,92.82
X$32004 544 583 545 644 645 cell_1rw
* cell instance $32005 r0 *1 168.495,92.82
X$32005 544 582 545 644 645 cell_1rw
* cell instance $32006 m0 *1 168.495,95.55
X$32006 544 584 545 644 645 cell_1rw
* cell instance $32007 r0 *1 168.495,95.55
X$32007 544 585 545 644 645 cell_1rw
* cell instance $32008 m0 *1 168.495,98.28
X$32008 544 586 545 644 645 cell_1rw
* cell instance $32009 r0 *1 168.495,98.28
X$32009 544 587 545 644 645 cell_1rw
* cell instance $32010 m0 *1 168.495,101.01
X$32010 544 588 545 644 645 cell_1rw
* cell instance $32011 r0 *1 168.495,101.01
X$32011 544 589 545 644 645 cell_1rw
* cell instance $32012 m0 *1 168.495,103.74
X$32012 544 590 545 644 645 cell_1rw
* cell instance $32013 r0 *1 168.495,103.74
X$32013 544 591 545 644 645 cell_1rw
* cell instance $32014 m0 *1 168.495,106.47
X$32014 544 593 545 644 645 cell_1rw
* cell instance $32015 r0 *1 168.495,106.47
X$32015 544 592 545 644 645 cell_1rw
* cell instance $32016 m0 *1 168.495,109.2
X$32016 544 594 545 644 645 cell_1rw
* cell instance $32017 r0 *1 168.495,109.2
X$32017 544 595 545 644 645 cell_1rw
* cell instance $32018 m0 *1 168.495,111.93
X$32018 544 597 545 644 645 cell_1rw
* cell instance $32019 m0 *1 168.495,114.66
X$32019 544 598 545 644 645 cell_1rw
* cell instance $32020 r0 *1 168.495,111.93
X$32020 544 596 545 644 645 cell_1rw
* cell instance $32021 r0 *1 168.495,114.66
X$32021 544 599 545 644 645 cell_1rw
* cell instance $32022 m0 *1 168.495,117.39
X$32022 544 600 545 644 645 cell_1rw
* cell instance $32023 r0 *1 168.495,117.39
X$32023 544 601 545 644 645 cell_1rw
* cell instance $32024 m0 *1 168.495,120.12
X$32024 544 602 545 644 645 cell_1rw
* cell instance $32025 m0 *1 168.495,122.85
X$32025 544 604 545 644 645 cell_1rw
* cell instance $32026 r0 *1 168.495,120.12
X$32026 544 603 545 644 645 cell_1rw
* cell instance $32027 r0 *1 168.495,122.85
X$32027 544 605 545 644 645 cell_1rw
* cell instance $32028 m0 *1 168.495,125.58
X$32028 544 606 545 644 645 cell_1rw
* cell instance $32029 r0 *1 168.495,125.58
X$32029 544 607 545 644 645 cell_1rw
* cell instance $32030 m0 *1 168.495,128.31
X$32030 544 609 545 644 645 cell_1rw
* cell instance $32031 m0 *1 168.495,131.04
X$32031 544 610 545 644 645 cell_1rw
* cell instance $32032 r0 *1 168.495,128.31
X$32032 544 608 545 644 645 cell_1rw
* cell instance $32033 m0 *1 168.495,133.77
X$32033 544 612 545 644 645 cell_1rw
* cell instance $32034 r0 *1 168.495,131.04
X$32034 544 611 545 644 645 cell_1rw
* cell instance $32035 r0 *1 168.495,133.77
X$32035 544 613 545 644 645 cell_1rw
* cell instance $32036 m0 *1 168.495,136.5
X$32036 544 615 545 644 645 cell_1rw
* cell instance $32037 m0 *1 168.495,139.23
X$32037 544 617 545 644 645 cell_1rw
* cell instance $32038 r0 *1 168.495,136.5
X$32038 544 614 545 644 645 cell_1rw
* cell instance $32039 m0 *1 168.495,141.96
X$32039 544 618 545 644 645 cell_1rw
* cell instance $32040 r0 *1 168.495,139.23
X$32040 544 616 545 644 645 cell_1rw
* cell instance $32041 r0 *1 168.495,141.96
X$32041 544 619 545 644 645 cell_1rw
* cell instance $32042 m0 *1 168.495,144.69
X$32042 544 620 545 644 645 cell_1rw
* cell instance $32043 r0 *1 168.495,144.69
X$32043 544 621 545 644 645 cell_1rw
* cell instance $32044 m0 *1 168.495,147.42
X$32044 544 622 545 644 645 cell_1rw
* cell instance $32045 r0 *1 168.495,147.42
X$32045 544 623 545 644 645 cell_1rw
* cell instance $32046 m0 *1 168.495,150.15
X$32046 544 624 545 644 645 cell_1rw
* cell instance $32047 r0 *1 168.495,150.15
X$32047 544 625 545 644 645 cell_1rw
* cell instance $32048 m0 *1 168.495,152.88
X$32048 544 626 545 644 645 cell_1rw
* cell instance $32049 m0 *1 168.495,155.61
X$32049 544 628 545 644 645 cell_1rw
* cell instance $32050 r0 *1 168.495,152.88
X$32050 544 627 545 644 645 cell_1rw
* cell instance $32051 r0 *1 168.495,155.61
X$32051 544 629 545 644 645 cell_1rw
* cell instance $32052 m0 *1 168.495,158.34
X$32052 544 630 545 644 645 cell_1rw
* cell instance $32053 m0 *1 168.495,161.07
X$32053 544 632 545 644 645 cell_1rw
* cell instance $32054 r0 *1 168.495,158.34
X$32054 544 631 545 644 645 cell_1rw
* cell instance $32055 r0 *1 168.495,161.07
X$32055 544 633 545 644 645 cell_1rw
* cell instance $32056 m0 *1 168.495,163.8
X$32056 544 634 545 644 645 cell_1rw
* cell instance $32057 m0 *1 168.495,166.53
X$32057 544 637 545 644 645 cell_1rw
* cell instance $32058 r0 *1 168.495,163.8
X$32058 544 635 545 644 645 cell_1rw
* cell instance $32059 r0 *1 168.495,166.53
X$32059 544 636 545 644 645 cell_1rw
* cell instance $32060 m0 *1 168.495,169.26
X$32060 544 639 545 644 645 cell_1rw
* cell instance $32061 r0 *1 168.495,169.26
X$32061 544 638 545 644 645 cell_1rw
* cell instance $32062 m0 *1 168.495,171.99
X$32062 544 640 545 644 645 cell_1rw
* cell instance $32063 r0 *1 168.495,171.99
X$32063 544 641 545 644 645 cell_1rw
* cell instance $32064 m0 *1 168.495,174.72
X$32064 544 642 545 644 645 cell_1rw
* cell instance $32065 r0 *1 168.495,174.72
X$32065 544 643 545 644 645 cell_1rw
* cell instance $32066 m0 *1 169.2,90.09
X$32066 546 581 547 644 645 cell_1rw
* cell instance $32067 r0 *1 169.2,90.09
X$32067 546 580 547 644 645 cell_1rw
* cell instance $32068 m0 *1 169.2,92.82
X$32068 546 583 547 644 645 cell_1rw
* cell instance $32069 r0 *1 169.2,92.82
X$32069 546 582 547 644 645 cell_1rw
* cell instance $32070 m0 *1 169.2,95.55
X$32070 546 584 547 644 645 cell_1rw
* cell instance $32071 r0 *1 169.2,95.55
X$32071 546 585 547 644 645 cell_1rw
* cell instance $32072 m0 *1 169.2,98.28
X$32072 546 586 547 644 645 cell_1rw
* cell instance $32073 m0 *1 169.2,101.01
X$32073 546 588 547 644 645 cell_1rw
* cell instance $32074 r0 *1 169.2,98.28
X$32074 546 587 547 644 645 cell_1rw
* cell instance $32075 r0 *1 169.2,101.01
X$32075 546 589 547 644 645 cell_1rw
* cell instance $32076 m0 *1 169.2,103.74
X$32076 546 590 547 644 645 cell_1rw
* cell instance $32077 r0 *1 169.2,103.74
X$32077 546 591 547 644 645 cell_1rw
* cell instance $32078 m0 *1 169.2,106.47
X$32078 546 593 547 644 645 cell_1rw
* cell instance $32079 r0 *1 169.2,106.47
X$32079 546 592 547 644 645 cell_1rw
* cell instance $32080 m0 *1 169.2,109.2
X$32080 546 594 547 644 645 cell_1rw
* cell instance $32081 r0 *1 169.2,109.2
X$32081 546 595 547 644 645 cell_1rw
* cell instance $32082 m0 *1 169.2,111.93
X$32082 546 597 547 644 645 cell_1rw
* cell instance $32083 r0 *1 169.2,111.93
X$32083 546 596 547 644 645 cell_1rw
* cell instance $32084 m0 *1 169.2,114.66
X$32084 546 598 547 644 645 cell_1rw
* cell instance $32085 r0 *1 169.2,114.66
X$32085 546 599 547 644 645 cell_1rw
* cell instance $32086 m0 *1 169.2,117.39
X$32086 546 600 547 644 645 cell_1rw
* cell instance $32087 m0 *1 169.2,120.12
X$32087 546 602 547 644 645 cell_1rw
* cell instance $32088 r0 *1 169.2,117.39
X$32088 546 601 547 644 645 cell_1rw
* cell instance $32089 r0 *1 169.2,120.12
X$32089 546 603 547 644 645 cell_1rw
* cell instance $32090 m0 *1 169.2,122.85
X$32090 546 604 547 644 645 cell_1rw
* cell instance $32091 r0 *1 169.2,122.85
X$32091 546 605 547 644 645 cell_1rw
* cell instance $32092 m0 *1 169.2,125.58
X$32092 546 606 547 644 645 cell_1rw
* cell instance $32093 r0 *1 169.2,125.58
X$32093 546 607 547 644 645 cell_1rw
* cell instance $32094 m0 *1 169.2,128.31
X$32094 546 609 547 644 645 cell_1rw
* cell instance $32095 r0 *1 169.2,128.31
X$32095 546 608 547 644 645 cell_1rw
* cell instance $32096 m0 *1 169.2,131.04
X$32096 546 610 547 644 645 cell_1rw
* cell instance $32097 r0 *1 169.2,131.04
X$32097 546 611 547 644 645 cell_1rw
* cell instance $32098 m0 *1 169.2,133.77
X$32098 546 612 547 644 645 cell_1rw
* cell instance $32099 r0 *1 169.2,133.77
X$32099 546 613 547 644 645 cell_1rw
* cell instance $32100 m0 *1 169.2,136.5
X$32100 546 615 547 644 645 cell_1rw
* cell instance $32101 m0 *1 169.2,139.23
X$32101 546 617 547 644 645 cell_1rw
* cell instance $32102 r0 *1 169.2,136.5
X$32102 546 614 547 644 645 cell_1rw
* cell instance $32103 r0 *1 169.2,139.23
X$32103 546 616 547 644 645 cell_1rw
* cell instance $32104 m0 *1 169.2,141.96
X$32104 546 618 547 644 645 cell_1rw
* cell instance $32105 r0 *1 169.2,141.96
X$32105 546 619 547 644 645 cell_1rw
* cell instance $32106 m0 *1 169.2,144.69
X$32106 546 620 547 644 645 cell_1rw
* cell instance $32107 r0 *1 169.2,144.69
X$32107 546 621 547 644 645 cell_1rw
* cell instance $32108 m0 *1 169.2,147.42
X$32108 546 622 547 644 645 cell_1rw
* cell instance $32109 r0 *1 169.2,147.42
X$32109 546 623 547 644 645 cell_1rw
* cell instance $32110 m0 *1 169.2,150.15
X$32110 546 624 547 644 645 cell_1rw
* cell instance $32111 r0 *1 169.2,150.15
X$32111 546 625 547 644 645 cell_1rw
* cell instance $32112 m0 *1 169.2,152.88
X$32112 546 626 547 644 645 cell_1rw
* cell instance $32113 m0 *1 169.2,155.61
X$32113 546 628 547 644 645 cell_1rw
* cell instance $32114 r0 *1 169.2,152.88
X$32114 546 627 547 644 645 cell_1rw
* cell instance $32115 r0 *1 169.2,155.61
X$32115 546 629 547 644 645 cell_1rw
* cell instance $32116 m0 *1 169.2,158.34
X$32116 546 630 547 644 645 cell_1rw
* cell instance $32117 r0 *1 169.2,158.34
X$32117 546 631 547 644 645 cell_1rw
* cell instance $32118 m0 *1 169.2,161.07
X$32118 546 632 547 644 645 cell_1rw
* cell instance $32119 r0 *1 169.2,161.07
X$32119 546 633 547 644 645 cell_1rw
* cell instance $32120 m0 *1 169.2,163.8
X$32120 546 634 547 644 645 cell_1rw
* cell instance $32121 r0 *1 169.2,163.8
X$32121 546 635 547 644 645 cell_1rw
* cell instance $32122 m0 *1 169.2,166.53
X$32122 546 637 547 644 645 cell_1rw
* cell instance $32123 r0 *1 169.2,166.53
X$32123 546 636 547 644 645 cell_1rw
* cell instance $32124 m0 *1 169.2,169.26
X$32124 546 639 547 644 645 cell_1rw
* cell instance $32125 r0 *1 169.2,169.26
X$32125 546 638 547 644 645 cell_1rw
* cell instance $32126 m0 *1 169.2,171.99
X$32126 546 640 547 644 645 cell_1rw
* cell instance $32127 r0 *1 169.2,171.99
X$32127 546 641 547 644 645 cell_1rw
* cell instance $32128 m0 *1 169.2,174.72
X$32128 546 642 547 644 645 cell_1rw
* cell instance $32129 r0 *1 169.2,174.72
X$32129 546 643 547 644 645 cell_1rw
* cell instance $32130 m0 *1 169.905,90.09
X$32130 548 581 549 644 645 cell_1rw
* cell instance $32131 r0 *1 169.905,90.09
X$32131 548 580 549 644 645 cell_1rw
* cell instance $32132 m0 *1 169.905,92.82
X$32132 548 583 549 644 645 cell_1rw
* cell instance $32133 r0 *1 169.905,92.82
X$32133 548 582 549 644 645 cell_1rw
* cell instance $32134 m0 *1 169.905,95.55
X$32134 548 584 549 644 645 cell_1rw
* cell instance $32135 r0 *1 169.905,95.55
X$32135 548 585 549 644 645 cell_1rw
* cell instance $32136 m0 *1 169.905,98.28
X$32136 548 586 549 644 645 cell_1rw
* cell instance $32137 r0 *1 169.905,98.28
X$32137 548 587 549 644 645 cell_1rw
* cell instance $32138 m0 *1 169.905,101.01
X$32138 548 588 549 644 645 cell_1rw
* cell instance $32139 r0 *1 169.905,101.01
X$32139 548 589 549 644 645 cell_1rw
* cell instance $32140 m0 *1 169.905,103.74
X$32140 548 590 549 644 645 cell_1rw
* cell instance $32141 r0 *1 169.905,103.74
X$32141 548 591 549 644 645 cell_1rw
* cell instance $32142 m0 *1 169.905,106.47
X$32142 548 593 549 644 645 cell_1rw
* cell instance $32143 m0 *1 169.905,109.2
X$32143 548 594 549 644 645 cell_1rw
* cell instance $32144 r0 *1 169.905,106.47
X$32144 548 592 549 644 645 cell_1rw
* cell instance $32145 r0 *1 169.905,109.2
X$32145 548 595 549 644 645 cell_1rw
* cell instance $32146 m0 *1 169.905,111.93
X$32146 548 597 549 644 645 cell_1rw
* cell instance $32147 r0 *1 169.905,111.93
X$32147 548 596 549 644 645 cell_1rw
* cell instance $32148 m0 *1 169.905,114.66
X$32148 548 598 549 644 645 cell_1rw
* cell instance $32149 r0 *1 169.905,114.66
X$32149 548 599 549 644 645 cell_1rw
* cell instance $32150 m0 *1 169.905,117.39
X$32150 548 600 549 644 645 cell_1rw
* cell instance $32151 r0 *1 169.905,117.39
X$32151 548 601 549 644 645 cell_1rw
* cell instance $32152 m0 *1 169.905,120.12
X$32152 548 602 549 644 645 cell_1rw
* cell instance $32153 r0 *1 169.905,120.12
X$32153 548 603 549 644 645 cell_1rw
* cell instance $32154 m0 *1 169.905,122.85
X$32154 548 604 549 644 645 cell_1rw
* cell instance $32155 r0 *1 169.905,122.85
X$32155 548 605 549 644 645 cell_1rw
* cell instance $32156 m0 *1 169.905,125.58
X$32156 548 606 549 644 645 cell_1rw
* cell instance $32157 r0 *1 169.905,125.58
X$32157 548 607 549 644 645 cell_1rw
* cell instance $32158 m0 *1 169.905,128.31
X$32158 548 609 549 644 645 cell_1rw
* cell instance $32159 r0 *1 169.905,128.31
X$32159 548 608 549 644 645 cell_1rw
* cell instance $32160 m0 *1 169.905,131.04
X$32160 548 610 549 644 645 cell_1rw
* cell instance $32161 r0 *1 169.905,131.04
X$32161 548 611 549 644 645 cell_1rw
* cell instance $32162 m0 *1 169.905,133.77
X$32162 548 612 549 644 645 cell_1rw
* cell instance $32163 r0 *1 169.905,133.77
X$32163 548 613 549 644 645 cell_1rw
* cell instance $32164 m0 *1 169.905,136.5
X$32164 548 615 549 644 645 cell_1rw
* cell instance $32165 r0 *1 169.905,136.5
X$32165 548 614 549 644 645 cell_1rw
* cell instance $32166 m0 *1 169.905,139.23
X$32166 548 617 549 644 645 cell_1rw
* cell instance $32167 r0 *1 169.905,139.23
X$32167 548 616 549 644 645 cell_1rw
* cell instance $32168 m0 *1 169.905,141.96
X$32168 548 618 549 644 645 cell_1rw
* cell instance $32169 r0 *1 169.905,141.96
X$32169 548 619 549 644 645 cell_1rw
* cell instance $32170 m0 *1 169.905,144.69
X$32170 548 620 549 644 645 cell_1rw
* cell instance $32171 r0 *1 169.905,144.69
X$32171 548 621 549 644 645 cell_1rw
* cell instance $32172 m0 *1 169.905,147.42
X$32172 548 622 549 644 645 cell_1rw
* cell instance $32173 r0 *1 169.905,147.42
X$32173 548 623 549 644 645 cell_1rw
* cell instance $32174 m0 *1 169.905,150.15
X$32174 548 624 549 644 645 cell_1rw
* cell instance $32175 r0 *1 169.905,150.15
X$32175 548 625 549 644 645 cell_1rw
* cell instance $32176 m0 *1 169.905,152.88
X$32176 548 626 549 644 645 cell_1rw
* cell instance $32177 r0 *1 169.905,152.88
X$32177 548 627 549 644 645 cell_1rw
* cell instance $32178 m0 *1 169.905,155.61
X$32178 548 628 549 644 645 cell_1rw
* cell instance $32179 r0 *1 169.905,155.61
X$32179 548 629 549 644 645 cell_1rw
* cell instance $32180 m0 *1 169.905,158.34
X$32180 548 630 549 644 645 cell_1rw
* cell instance $32181 r0 *1 169.905,158.34
X$32181 548 631 549 644 645 cell_1rw
* cell instance $32182 m0 *1 169.905,161.07
X$32182 548 632 549 644 645 cell_1rw
* cell instance $32183 r0 *1 169.905,161.07
X$32183 548 633 549 644 645 cell_1rw
* cell instance $32184 m0 *1 169.905,163.8
X$32184 548 634 549 644 645 cell_1rw
* cell instance $32185 r0 *1 169.905,163.8
X$32185 548 635 549 644 645 cell_1rw
* cell instance $32186 m0 *1 169.905,166.53
X$32186 548 637 549 644 645 cell_1rw
* cell instance $32187 r0 *1 169.905,166.53
X$32187 548 636 549 644 645 cell_1rw
* cell instance $32188 m0 *1 169.905,169.26
X$32188 548 639 549 644 645 cell_1rw
* cell instance $32189 r0 *1 169.905,169.26
X$32189 548 638 549 644 645 cell_1rw
* cell instance $32190 m0 *1 169.905,171.99
X$32190 548 640 549 644 645 cell_1rw
* cell instance $32191 r0 *1 169.905,171.99
X$32191 548 641 549 644 645 cell_1rw
* cell instance $32192 m0 *1 169.905,174.72
X$32192 548 642 549 644 645 cell_1rw
* cell instance $32193 r0 *1 169.905,174.72
X$32193 548 643 549 644 645 cell_1rw
* cell instance $32194 m0 *1 170.61,90.09
X$32194 550 581 551 644 645 cell_1rw
* cell instance $32195 r0 *1 170.61,90.09
X$32195 550 580 551 644 645 cell_1rw
* cell instance $32196 m0 *1 170.61,92.82
X$32196 550 583 551 644 645 cell_1rw
* cell instance $32197 r0 *1 170.61,92.82
X$32197 550 582 551 644 645 cell_1rw
* cell instance $32198 m0 *1 170.61,95.55
X$32198 550 584 551 644 645 cell_1rw
* cell instance $32199 r0 *1 170.61,95.55
X$32199 550 585 551 644 645 cell_1rw
* cell instance $32200 m0 *1 170.61,98.28
X$32200 550 586 551 644 645 cell_1rw
* cell instance $32201 r0 *1 170.61,98.28
X$32201 550 587 551 644 645 cell_1rw
* cell instance $32202 m0 *1 170.61,101.01
X$32202 550 588 551 644 645 cell_1rw
* cell instance $32203 r0 *1 170.61,101.01
X$32203 550 589 551 644 645 cell_1rw
* cell instance $32204 m0 *1 170.61,103.74
X$32204 550 590 551 644 645 cell_1rw
* cell instance $32205 r0 *1 170.61,103.74
X$32205 550 591 551 644 645 cell_1rw
* cell instance $32206 m0 *1 170.61,106.47
X$32206 550 593 551 644 645 cell_1rw
* cell instance $32207 r0 *1 170.61,106.47
X$32207 550 592 551 644 645 cell_1rw
* cell instance $32208 m0 *1 170.61,109.2
X$32208 550 594 551 644 645 cell_1rw
* cell instance $32209 r0 *1 170.61,109.2
X$32209 550 595 551 644 645 cell_1rw
* cell instance $32210 m0 *1 170.61,111.93
X$32210 550 597 551 644 645 cell_1rw
* cell instance $32211 r0 *1 170.61,111.93
X$32211 550 596 551 644 645 cell_1rw
* cell instance $32212 m0 *1 170.61,114.66
X$32212 550 598 551 644 645 cell_1rw
* cell instance $32213 r0 *1 170.61,114.66
X$32213 550 599 551 644 645 cell_1rw
* cell instance $32214 m0 *1 170.61,117.39
X$32214 550 600 551 644 645 cell_1rw
* cell instance $32215 r0 *1 170.61,117.39
X$32215 550 601 551 644 645 cell_1rw
* cell instance $32216 m0 *1 170.61,120.12
X$32216 550 602 551 644 645 cell_1rw
* cell instance $32217 r0 *1 170.61,120.12
X$32217 550 603 551 644 645 cell_1rw
* cell instance $32218 m0 *1 170.61,122.85
X$32218 550 604 551 644 645 cell_1rw
* cell instance $32219 r0 *1 170.61,122.85
X$32219 550 605 551 644 645 cell_1rw
* cell instance $32220 m0 *1 170.61,125.58
X$32220 550 606 551 644 645 cell_1rw
* cell instance $32221 r0 *1 170.61,125.58
X$32221 550 607 551 644 645 cell_1rw
* cell instance $32222 m0 *1 170.61,128.31
X$32222 550 609 551 644 645 cell_1rw
* cell instance $32223 r0 *1 170.61,128.31
X$32223 550 608 551 644 645 cell_1rw
* cell instance $32224 m0 *1 170.61,131.04
X$32224 550 610 551 644 645 cell_1rw
* cell instance $32225 r0 *1 170.61,131.04
X$32225 550 611 551 644 645 cell_1rw
* cell instance $32226 m0 *1 170.61,133.77
X$32226 550 612 551 644 645 cell_1rw
* cell instance $32227 r0 *1 170.61,133.77
X$32227 550 613 551 644 645 cell_1rw
* cell instance $32228 m0 *1 170.61,136.5
X$32228 550 615 551 644 645 cell_1rw
* cell instance $32229 r0 *1 170.61,136.5
X$32229 550 614 551 644 645 cell_1rw
* cell instance $32230 m0 *1 170.61,139.23
X$32230 550 617 551 644 645 cell_1rw
* cell instance $32231 r0 *1 170.61,139.23
X$32231 550 616 551 644 645 cell_1rw
* cell instance $32232 m0 *1 170.61,141.96
X$32232 550 618 551 644 645 cell_1rw
* cell instance $32233 m0 *1 170.61,144.69
X$32233 550 620 551 644 645 cell_1rw
* cell instance $32234 r0 *1 170.61,141.96
X$32234 550 619 551 644 645 cell_1rw
* cell instance $32235 r0 *1 170.61,144.69
X$32235 550 621 551 644 645 cell_1rw
* cell instance $32236 m0 *1 170.61,147.42
X$32236 550 622 551 644 645 cell_1rw
* cell instance $32237 m0 *1 170.61,150.15
X$32237 550 624 551 644 645 cell_1rw
* cell instance $32238 r0 *1 170.61,147.42
X$32238 550 623 551 644 645 cell_1rw
* cell instance $32239 r0 *1 170.61,150.15
X$32239 550 625 551 644 645 cell_1rw
* cell instance $32240 m0 *1 170.61,152.88
X$32240 550 626 551 644 645 cell_1rw
* cell instance $32241 m0 *1 170.61,155.61
X$32241 550 628 551 644 645 cell_1rw
* cell instance $32242 r0 *1 170.61,152.88
X$32242 550 627 551 644 645 cell_1rw
* cell instance $32243 r0 *1 170.61,155.61
X$32243 550 629 551 644 645 cell_1rw
* cell instance $32244 m0 *1 170.61,158.34
X$32244 550 630 551 644 645 cell_1rw
* cell instance $32245 r0 *1 170.61,158.34
X$32245 550 631 551 644 645 cell_1rw
* cell instance $32246 m0 *1 170.61,161.07
X$32246 550 632 551 644 645 cell_1rw
* cell instance $32247 r0 *1 170.61,161.07
X$32247 550 633 551 644 645 cell_1rw
* cell instance $32248 m0 *1 170.61,163.8
X$32248 550 634 551 644 645 cell_1rw
* cell instance $32249 r0 *1 170.61,163.8
X$32249 550 635 551 644 645 cell_1rw
* cell instance $32250 m0 *1 170.61,166.53
X$32250 550 637 551 644 645 cell_1rw
* cell instance $32251 r0 *1 170.61,166.53
X$32251 550 636 551 644 645 cell_1rw
* cell instance $32252 m0 *1 170.61,169.26
X$32252 550 639 551 644 645 cell_1rw
* cell instance $32253 r0 *1 170.61,169.26
X$32253 550 638 551 644 645 cell_1rw
* cell instance $32254 m0 *1 170.61,171.99
X$32254 550 640 551 644 645 cell_1rw
* cell instance $32255 m0 *1 170.61,174.72
X$32255 550 642 551 644 645 cell_1rw
* cell instance $32256 r0 *1 170.61,171.99
X$32256 550 641 551 644 645 cell_1rw
* cell instance $32257 r0 *1 170.61,174.72
X$32257 550 643 551 644 645 cell_1rw
* cell instance $32258 m0 *1 171.315,90.09
X$32258 552 581 553 644 645 cell_1rw
* cell instance $32259 r0 *1 171.315,90.09
X$32259 552 580 553 644 645 cell_1rw
* cell instance $32260 m0 *1 171.315,92.82
X$32260 552 583 553 644 645 cell_1rw
* cell instance $32261 r0 *1 171.315,92.82
X$32261 552 582 553 644 645 cell_1rw
* cell instance $32262 m0 *1 171.315,95.55
X$32262 552 584 553 644 645 cell_1rw
* cell instance $32263 r0 *1 171.315,95.55
X$32263 552 585 553 644 645 cell_1rw
* cell instance $32264 m0 *1 171.315,98.28
X$32264 552 586 553 644 645 cell_1rw
* cell instance $32265 r0 *1 171.315,98.28
X$32265 552 587 553 644 645 cell_1rw
* cell instance $32266 m0 *1 171.315,101.01
X$32266 552 588 553 644 645 cell_1rw
* cell instance $32267 m0 *1 171.315,103.74
X$32267 552 590 553 644 645 cell_1rw
* cell instance $32268 r0 *1 171.315,101.01
X$32268 552 589 553 644 645 cell_1rw
* cell instance $32269 r0 *1 171.315,103.74
X$32269 552 591 553 644 645 cell_1rw
* cell instance $32270 m0 *1 171.315,106.47
X$32270 552 593 553 644 645 cell_1rw
* cell instance $32271 r0 *1 171.315,106.47
X$32271 552 592 553 644 645 cell_1rw
* cell instance $32272 m0 *1 171.315,109.2
X$32272 552 594 553 644 645 cell_1rw
* cell instance $32273 r0 *1 171.315,109.2
X$32273 552 595 553 644 645 cell_1rw
* cell instance $32274 m0 *1 171.315,111.93
X$32274 552 597 553 644 645 cell_1rw
* cell instance $32275 r0 *1 171.315,111.93
X$32275 552 596 553 644 645 cell_1rw
* cell instance $32276 m0 *1 171.315,114.66
X$32276 552 598 553 644 645 cell_1rw
* cell instance $32277 r0 *1 171.315,114.66
X$32277 552 599 553 644 645 cell_1rw
* cell instance $32278 m0 *1 171.315,117.39
X$32278 552 600 553 644 645 cell_1rw
* cell instance $32279 r0 *1 171.315,117.39
X$32279 552 601 553 644 645 cell_1rw
* cell instance $32280 m0 *1 171.315,120.12
X$32280 552 602 553 644 645 cell_1rw
* cell instance $32281 r0 *1 171.315,120.12
X$32281 552 603 553 644 645 cell_1rw
* cell instance $32282 m0 *1 171.315,122.85
X$32282 552 604 553 644 645 cell_1rw
* cell instance $32283 r0 *1 171.315,122.85
X$32283 552 605 553 644 645 cell_1rw
* cell instance $32284 m0 *1 171.315,125.58
X$32284 552 606 553 644 645 cell_1rw
* cell instance $32285 r0 *1 171.315,125.58
X$32285 552 607 553 644 645 cell_1rw
* cell instance $32286 m0 *1 171.315,128.31
X$32286 552 609 553 644 645 cell_1rw
* cell instance $32287 r0 *1 171.315,128.31
X$32287 552 608 553 644 645 cell_1rw
* cell instance $32288 m0 *1 171.315,131.04
X$32288 552 610 553 644 645 cell_1rw
* cell instance $32289 r0 *1 171.315,131.04
X$32289 552 611 553 644 645 cell_1rw
* cell instance $32290 m0 *1 171.315,133.77
X$32290 552 612 553 644 645 cell_1rw
* cell instance $32291 r0 *1 171.315,133.77
X$32291 552 613 553 644 645 cell_1rw
* cell instance $32292 m0 *1 171.315,136.5
X$32292 552 615 553 644 645 cell_1rw
* cell instance $32293 r0 *1 171.315,136.5
X$32293 552 614 553 644 645 cell_1rw
* cell instance $32294 m0 *1 171.315,139.23
X$32294 552 617 553 644 645 cell_1rw
* cell instance $32295 r0 *1 171.315,139.23
X$32295 552 616 553 644 645 cell_1rw
* cell instance $32296 m0 *1 171.315,141.96
X$32296 552 618 553 644 645 cell_1rw
* cell instance $32297 m0 *1 171.315,144.69
X$32297 552 620 553 644 645 cell_1rw
* cell instance $32298 r0 *1 171.315,141.96
X$32298 552 619 553 644 645 cell_1rw
* cell instance $32299 r0 *1 171.315,144.69
X$32299 552 621 553 644 645 cell_1rw
* cell instance $32300 m0 *1 171.315,147.42
X$32300 552 622 553 644 645 cell_1rw
* cell instance $32301 r0 *1 171.315,147.42
X$32301 552 623 553 644 645 cell_1rw
* cell instance $32302 m0 *1 171.315,150.15
X$32302 552 624 553 644 645 cell_1rw
* cell instance $32303 m0 *1 171.315,152.88
X$32303 552 626 553 644 645 cell_1rw
* cell instance $32304 r0 *1 171.315,150.15
X$32304 552 625 553 644 645 cell_1rw
* cell instance $32305 m0 *1 171.315,155.61
X$32305 552 628 553 644 645 cell_1rw
* cell instance $32306 r0 *1 171.315,152.88
X$32306 552 627 553 644 645 cell_1rw
* cell instance $32307 r0 *1 171.315,155.61
X$32307 552 629 553 644 645 cell_1rw
* cell instance $32308 m0 *1 171.315,158.34
X$32308 552 630 553 644 645 cell_1rw
* cell instance $32309 r0 *1 171.315,158.34
X$32309 552 631 553 644 645 cell_1rw
* cell instance $32310 m0 *1 171.315,161.07
X$32310 552 632 553 644 645 cell_1rw
* cell instance $32311 r0 *1 171.315,161.07
X$32311 552 633 553 644 645 cell_1rw
* cell instance $32312 m0 *1 171.315,163.8
X$32312 552 634 553 644 645 cell_1rw
* cell instance $32313 r0 *1 171.315,163.8
X$32313 552 635 553 644 645 cell_1rw
* cell instance $32314 m0 *1 171.315,166.53
X$32314 552 637 553 644 645 cell_1rw
* cell instance $32315 r0 *1 171.315,166.53
X$32315 552 636 553 644 645 cell_1rw
* cell instance $32316 m0 *1 171.315,169.26
X$32316 552 639 553 644 645 cell_1rw
* cell instance $32317 r0 *1 171.315,169.26
X$32317 552 638 553 644 645 cell_1rw
* cell instance $32318 m0 *1 171.315,171.99
X$32318 552 640 553 644 645 cell_1rw
* cell instance $32319 m0 *1 171.315,174.72
X$32319 552 642 553 644 645 cell_1rw
* cell instance $32320 r0 *1 171.315,171.99
X$32320 552 641 553 644 645 cell_1rw
* cell instance $32321 r0 *1 171.315,174.72
X$32321 552 643 553 644 645 cell_1rw
* cell instance $32322 m0 *1 172.02,90.09
X$32322 554 581 555 644 645 cell_1rw
* cell instance $32323 r0 *1 172.02,90.09
X$32323 554 580 555 644 645 cell_1rw
* cell instance $32324 m0 *1 172.02,92.82
X$32324 554 583 555 644 645 cell_1rw
* cell instance $32325 r0 *1 172.02,92.82
X$32325 554 582 555 644 645 cell_1rw
* cell instance $32326 m0 *1 172.02,95.55
X$32326 554 584 555 644 645 cell_1rw
* cell instance $32327 r0 *1 172.02,95.55
X$32327 554 585 555 644 645 cell_1rw
* cell instance $32328 m0 *1 172.02,98.28
X$32328 554 586 555 644 645 cell_1rw
* cell instance $32329 r0 *1 172.02,98.28
X$32329 554 587 555 644 645 cell_1rw
* cell instance $32330 m0 *1 172.02,101.01
X$32330 554 588 555 644 645 cell_1rw
* cell instance $32331 r0 *1 172.02,101.01
X$32331 554 589 555 644 645 cell_1rw
* cell instance $32332 m0 *1 172.02,103.74
X$32332 554 590 555 644 645 cell_1rw
* cell instance $32333 r0 *1 172.02,103.74
X$32333 554 591 555 644 645 cell_1rw
* cell instance $32334 m0 *1 172.02,106.47
X$32334 554 593 555 644 645 cell_1rw
* cell instance $32335 r0 *1 172.02,106.47
X$32335 554 592 555 644 645 cell_1rw
* cell instance $32336 m0 *1 172.02,109.2
X$32336 554 594 555 644 645 cell_1rw
* cell instance $32337 r0 *1 172.02,109.2
X$32337 554 595 555 644 645 cell_1rw
* cell instance $32338 m0 *1 172.02,111.93
X$32338 554 597 555 644 645 cell_1rw
* cell instance $32339 r0 *1 172.02,111.93
X$32339 554 596 555 644 645 cell_1rw
* cell instance $32340 m0 *1 172.02,114.66
X$32340 554 598 555 644 645 cell_1rw
* cell instance $32341 r0 *1 172.02,114.66
X$32341 554 599 555 644 645 cell_1rw
* cell instance $32342 m0 *1 172.02,117.39
X$32342 554 600 555 644 645 cell_1rw
* cell instance $32343 r0 *1 172.02,117.39
X$32343 554 601 555 644 645 cell_1rw
* cell instance $32344 m0 *1 172.02,120.12
X$32344 554 602 555 644 645 cell_1rw
* cell instance $32345 r0 *1 172.02,120.12
X$32345 554 603 555 644 645 cell_1rw
* cell instance $32346 m0 *1 172.02,122.85
X$32346 554 604 555 644 645 cell_1rw
* cell instance $32347 r0 *1 172.02,122.85
X$32347 554 605 555 644 645 cell_1rw
* cell instance $32348 m0 *1 172.02,125.58
X$32348 554 606 555 644 645 cell_1rw
* cell instance $32349 r0 *1 172.02,125.58
X$32349 554 607 555 644 645 cell_1rw
* cell instance $32350 m0 *1 172.02,128.31
X$32350 554 609 555 644 645 cell_1rw
* cell instance $32351 r0 *1 172.02,128.31
X$32351 554 608 555 644 645 cell_1rw
* cell instance $32352 m0 *1 172.02,131.04
X$32352 554 610 555 644 645 cell_1rw
* cell instance $32353 r0 *1 172.02,131.04
X$32353 554 611 555 644 645 cell_1rw
* cell instance $32354 m0 *1 172.02,133.77
X$32354 554 612 555 644 645 cell_1rw
* cell instance $32355 r0 *1 172.02,133.77
X$32355 554 613 555 644 645 cell_1rw
* cell instance $32356 m0 *1 172.02,136.5
X$32356 554 615 555 644 645 cell_1rw
* cell instance $32357 r0 *1 172.02,136.5
X$32357 554 614 555 644 645 cell_1rw
* cell instance $32358 m0 *1 172.02,139.23
X$32358 554 617 555 644 645 cell_1rw
* cell instance $32359 r0 *1 172.02,139.23
X$32359 554 616 555 644 645 cell_1rw
* cell instance $32360 m0 *1 172.02,141.96
X$32360 554 618 555 644 645 cell_1rw
* cell instance $32361 r0 *1 172.02,141.96
X$32361 554 619 555 644 645 cell_1rw
* cell instance $32362 m0 *1 172.02,144.69
X$32362 554 620 555 644 645 cell_1rw
* cell instance $32363 r0 *1 172.02,144.69
X$32363 554 621 555 644 645 cell_1rw
* cell instance $32364 m0 *1 172.02,147.42
X$32364 554 622 555 644 645 cell_1rw
* cell instance $32365 r0 *1 172.02,147.42
X$32365 554 623 555 644 645 cell_1rw
* cell instance $32366 m0 *1 172.02,150.15
X$32366 554 624 555 644 645 cell_1rw
* cell instance $32367 r0 *1 172.02,150.15
X$32367 554 625 555 644 645 cell_1rw
* cell instance $32368 m0 *1 172.02,152.88
X$32368 554 626 555 644 645 cell_1rw
* cell instance $32369 m0 *1 172.02,155.61
X$32369 554 628 555 644 645 cell_1rw
* cell instance $32370 r0 *1 172.02,152.88
X$32370 554 627 555 644 645 cell_1rw
* cell instance $32371 r0 *1 172.02,155.61
X$32371 554 629 555 644 645 cell_1rw
* cell instance $32372 m0 *1 172.02,158.34
X$32372 554 630 555 644 645 cell_1rw
* cell instance $32373 r0 *1 172.02,158.34
X$32373 554 631 555 644 645 cell_1rw
* cell instance $32374 m0 *1 172.02,161.07
X$32374 554 632 555 644 645 cell_1rw
* cell instance $32375 r0 *1 172.02,161.07
X$32375 554 633 555 644 645 cell_1rw
* cell instance $32376 m0 *1 172.02,163.8
X$32376 554 634 555 644 645 cell_1rw
* cell instance $32377 r0 *1 172.02,163.8
X$32377 554 635 555 644 645 cell_1rw
* cell instance $32378 m0 *1 172.02,166.53
X$32378 554 637 555 644 645 cell_1rw
* cell instance $32379 r0 *1 172.02,166.53
X$32379 554 636 555 644 645 cell_1rw
* cell instance $32380 m0 *1 172.02,169.26
X$32380 554 639 555 644 645 cell_1rw
* cell instance $32381 r0 *1 172.02,169.26
X$32381 554 638 555 644 645 cell_1rw
* cell instance $32382 m0 *1 172.02,171.99
X$32382 554 640 555 644 645 cell_1rw
* cell instance $32383 m0 *1 172.02,174.72
X$32383 554 642 555 644 645 cell_1rw
* cell instance $32384 r0 *1 172.02,171.99
X$32384 554 641 555 644 645 cell_1rw
* cell instance $32385 r0 *1 172.02,174.72
X$32385 554 643 555 644 645 cell_1rw
* cell instance $32386 m0 *1 172.725,90.09
X$32386 556 581 557 644 645 cell_1rw
* cell instance $32387 r0 *1 172.725,90.09
X$32387 556 580 557 644 645 cell_1rw
* cell instance $32388 m0 *1 172.725,92.82
X$32388 556 583 557 644 645 cell_1rw
* cell instance $32389 r0 *1 172.725,92.82
X$32389 556 582 557 644 645 cell_1rw
* cell instance $32390 m0 *1 172.725,95.55
X$32390 556 584 557 644 645 cell_1rw
* cell instance $32391 r0 *1 172.725,95.55
X$32391 556 585 557 644 645 cell_1rw
* cell instance $32392 m0 *1 172.725,98.28
X$32392 556 586 557 644 645 cell_1rw
* cell instance $32393 m0 *1 172.725,101.01
X$32393 556 588 557 644 645 cell_1rw
* cell instance $32394 r0 *1 172.725,98.28
X$32394 556 587 557 644 645 cell_1rw
* cell instance $32395 r0 *1 172.725,101.01
X$32395 556 589 557 644 645 cell_1rw
* cell instance $32396 m0 *1 172.725,103.74
X$32396 556 590 557 644 645 cell_1rw
* cell instance $32397 m0 *1 172.725,106.47
X$32397 556 593 557 644 645 cell_1rw
* cell instance $32398 r0 *1 172.725,103.74
X$32398 556 591 557 644 645 cell_1rw
* cell instance $32399 r0 *1 172.725,106.47
X$32399 556 592 557 644 645 cell_1rw
* cell instance $32400 m0 *1 172.725,109.2
X$32400 556 594 557 644 645 cell_1rw
* cell instance $32401 r0 *1 172.725,109.2
X$32401 556 595 557 644 645 cell_1rw
* cell instance $32402 m0 *1 172.725,111.93
X$32402 556 597 557 644 645 cell_1rw
* cell instance $32403 m0 *1 172.725,114.66
X$32403 556 598 557 644 645 cell_1rw
* cell instance $32404 r0 *1 172.725,111.93
X$32404 556 596 557 644 645 cell_1rw
* cell instance $32405 r0 *1 172.725,114.66
X$32405 556 599 557 644 645 cell_1rw
* cell instance $32406 m0 *1 172.725,117.39
X$32406 556 600 557 644 645 cell_1rw
* cell instance $32407 r0 *1 172.725,117.39
X$32407 556 601 557 644 645 cell_1rw
* cell instance $32408 m0 *1 172.725,120.12
X$32408 556 602 557 644 645 cell_1rw
* cell instance $32409 r0 *1 172.725,120.12
X$32409 556 603 557 644 645 cell_1rw
* cell instance $32410 m0 *1 172.725,122.85
X$32410 556 604 557 644 645 cell_1rw
* cell instance $32411 r0 *1 172.725,122.85
X$32411 556 605 557 644 645 cell_1rw
* cell instance $32412 m0 *1 172.725,125.58
X$32412 556 606 557 644 645 cell_1rw
* cell instance $32413 m0 *1 172.725,128.31
X$32413 556 609 557 644 645 cell_1rw
* cell instance $32414 r0 *1 172.725,125.58
X$32414 556 607 557 644 645 cell_1rw
* cell instance $32415 r0 *1 172.725,128.31
X$32415 556 608 557 644 645 cell_1rw
* cell instance $32416 m0 *1 172.725,131.04
X$32416 556 610 557 644 645 cell_1rw
* cell instance $32417 r0 *1 172.725,131.04
X$32417 556 611 557 644 645 cell_1rw
* cell instance $32418 m0 *1 172.725,133.77
X$32418 556 612 557 644 645 cell_1rw
* cell instance $32419 m0 *1 172.725,136.5
X$32419 556 615 557 644 645 cell_1rw
* cell instance $32420 r0 *1 172.725,133.77
X$32420 556 613 557 644 645 cell_1rw
* cell instance $32421 r0 *1 172.725,136.5
X$32421 556 614 557 644 645 cell_1rw
* cell instance $32422 m0 *1 172.725,139.23
X$32422 556 617 557 644 645 cell_1rw
* cell instance $32423 m0 *1 172.725,141.96
X$32423 556 618 557 644 645 cell_1rw
* cell instance $32424 r0 *1 172.725,139.23
X$32424 556 616 557 644 645 cell_1rw
* cell instance $32425 r0 *1 172.725,141.96
X$32425 556 619 557 644 645 cell_1rw
* cell instance $32426 m0 *1 172.725,144.69
X$32426 556 620 557 644 645 cell_1rw
* cell instance $32427 r0 *1 172.725,144.69
X$32427 556 621 557 644 645 cell_1rw
* cell instance $32428 m0 *1 172.725,147.42
X$32428 556 622 557 644 645 cell_1rw
* cell instance $32429 r0 *1 172.725,147.42
X$32429 556 623 557 644 645 cell_1rw
* cell instance $32430 m0 *1 172.725,150.15
X$32430 556 624 557 644 645 cell_1rw
* cell instance $32431 r0 *1 172.725,150.15
X$32431 556 625 557 644 645 cell_1rw
* cell instance $32432 m0 *1 172.725,152.88
X$32432 556 626 557 644 645 cell_1rw
* cell instance $32433 r0 *1 172.725,152.88
X$32433 556 627 557 644 645 cell_1rw
* cell instance $32434 m0 *1 172.725,155.61
X$32434 556 628 557 644 645 cell_1rw
* cell instance $32435 r0 *1 172.725,155.61
X$32435 556 629 557 644 645 cell_1rw
* cell instance $32436 m0 *1 172.725,158.34
X$32436 556 630 557 644 645 cell_1rw
* cell instance $32437 r0 *1 172.725,158.34
X$32437 556 631 557 644 645 cell_1rw
* cell instance $32438 m0 *1 172.725,161.07
X$32438 556 632 557 644 645 cell_1rw
* cell instance $32439 r0 *1 172.725,161.07
X$32439 556 633 557 644 645 cell_1rw
* cell instance $32440 m0 *1 172.725,163.8
X$32440 556 634 557 644 645 cell_1rw
* cell instance $32441 r0 *1 172.725,163.8
X$32441 556 635 557 644 645 cell_1rw
* cell instance $32442 m0 *1 172.725,166.53
X$32442 556 637 557 644 645 cell_1rw
* cell instance $32443 m0 *1 172.725,169.26
X$32443 556 639 557 644 645 cell_1rw
* cell instance $32444 r0 *1 172.725,166.53
X$32444 556 636 557 644 645 cell_1rw
* cell instance $32445 r0 *1 172.725,169.26
X$32445 556 638 557 644 645 cell_1rw
* cell instance $32446 m0 *1 172.725,171.99
X$32446 556 640 557 644 645 cell_1rw
* cell instance $32447 r0 *1 172.725,171.99
X$32447 556 641 557 644 645 cell_1rw
* cell instance $32448 m0 *1 172.725,174.72
X$32448 556 642 557 644 645 cell_1rw
* cell instance $32449 r0 *1 172.725,174.72
X$32449 556 643 557 644 645 cell_1rw
* cell instance $32450 m0 *1 173.43,90.09
X$32450 558 581 559 644 645 cell_1rw
* cell instance $32451 r0 *1 173.43,90.09
X$32451 558 580 559 644 645 cell_1rw
* cell instance $32452 m0 *1 173.43,92.82
X$32452 558 583 559 644 645 cell_1rw
* cell instance $32453 r0 *1 173.43,92.82
X$32453 558 582 559 644 645 cell_1rw
* cell instance $32454 m0 *1 173.43,95.55
X$32454 558 584 559 644 645 cell_1rw
* cell instance $32455 r0 *1 173.43,95.55
X$32455 558 585 559 644 645 cell_1rw
* cell instance $32456 m0 *1 173.43,98.28
X$32456 558 586 559 644 645 cell_1rw
* cell instance $32457 r0 *1 173.43,98.28
X$32457 558 587 559 644 645 cell_1rw
* cell instance $32458 m0 *1 173.43,101.01
X$32458 558 588 559 644 645 cell_1rw
* cell instance $32459 r0 *1 173.43,101.01
X$32459 558 589 559 644 645 cell_1rw
* cell instance $32460 m0 *1 173.43,103.74
X$32460 558 590 559 644 645 cell_1rw
* cell instance $32461 m0 *1 173.43,106.47
X$32461 558 593 559 644 645 cell_1rw
* cell instance $32462 r0 *1 173.43,103.74
X$32462 558 591 559 644 645 cell_1rw
* cell instance $32463 r0 *1 173.43,106.47
X$32463 558 592 559 644 645 cell_1rw
* cell instance $32464 m0 *1 173.43,109.2
X$32464 558 594 559 644 645 cell_1rw
* cell instance $32465 m0 *1 173.43,111.93
X$32465 558 597 559 644 645 cell_1rw
* cell instance $32466 r0 *1 173.43,109.2
X$32466 558 595 559 644 645 cell_1rw
* cell instance $32467 r0 *1 173.43,111.93
X$32467 558 596 559 644 645 cell_1rw
* cell instance $32468 m0 *1 173.43,114.66
X$32468 558 598 559 644 645 cell_1rw
* cell instance $32469 m0 *1 173.43,117.39
X$32469 558 600 559 644 645 cell_1rw
* cell instance $32470 r0 *1 173.43,114.66
X$32470 558 599 559 644 645 cell_1rw
* cell instance $32471 r0 *1 173.43,117.39
X$32471 558 601 559 644 645 cell_1rw
* cell instance $32472 m0 *1 173.43,120.12
X$32472 558 602 559 644 645 cell_1rw
* cell instance $32473 r0 *1 173.43,120.12
X$32473 558 603 559 644 645 cell_1rw
* cell instance $32474 m0 *1 173.43,122.85
X$32474 558 604 559 644 645 cell_1rw
* cell instance $32475 r0 *1 173.43,122.85
X$32475 558 605 559 644 645 cell_1rw
* cell instance $32476 m0 *1 173.43,125.58
X$32476 558 606 559 644 645 cell_1rw
* cell instance $32477 r0 *1 173.43,125.58
X$32477 558 607 559 644 645 cell_1rw
* cell instance $32478 m0 *1 173.43,128.31
X$32478 558 609 559 644 645 cell_1rw
* cell instance $32479 r0 *1 173.43,128.31
X$32479 558 608 559 644 645 cell_1rw
* cell instance $32480 m0 *1 173.43,131.04
X$32480 558 610 559 644 645 cell_1rw
* cell instance $32481 r0 *1 173.43,131.04
X$32481 558 611 559 644 645 cell_1rw
* cell instance $32482 m0 *1 173.43,133.77
X$32482 558 612 559 644 645 cell_1rw
* cell instance $32483 r0 *1 173.43,133.77
X$32483 558 613 559 644 645 cell_1rw
* cell instance $32484 m0 *1 173.43,136.5
X$32484 558 615 559 644 645 cell_1rw
* cell instance $32485 r0 *1 173.43,136.5
X$32485 558 614 559 644 645 cell_1rw
* cell instance $32486 m0 *1 173.43,139.23
X$32486 558 617 559 644 645 cell_1rw
* cell instance $32487 r0 *1 173.43,139.23
X$32487 558 616 559 644 645 cell_1rw
* cell instance $32488 m0 *1 173.43,141.96
X$32488 558 618 559 644 645 cell_1rw
* cell instance $32489 r0 *1 173.43,141.96
X$32489 558 619 559 644 645 cell_1rw
* cell instance $32490 m0 *1 173.43,144.69
X$32490 558 620 559 644 645 cell_1rw
* cell instance $32491 r0 *1 173.43,144.69
X$32491 558 621 559 644 645 cell_1rw
* cell instance $32492 m0 *1 173.43,147.42
X$32492 558 622 559 644 645 cell_1rw
* cell instance $32493 r0 *1 173.43,147.42
X$32493 558 623 559 644 645 cell_1rw
* cell instance $32494 m0 *1 173.43,150.15
X$32494 558 624 559 644 645 cell_1rw
* cell instance $32495 r0 *1 173.43,150.15
X$32495 558 625 559 644 645 cell_1rw
* cell instance $32496 m0 *1 173.43,152.88
X$32496 558 626 559 644 645 cell_1rw
* cell instance $32497 r0 *1 173.43,152.88
X$32497 558 627 559 644 645 cell_1rw
* cell instance $32498 m0 *1 173.43,155.61
X$32498 558 628 559 644 645 cell_1rw
* cell instance $32499 r0 *1 173.43,155.61
X$32499 558 629 559 644 645 cell_1rw
* cell instance $32500 m0 *1 173.43,158.34
X$32500 558 630 559 644 645 cell_1rw
* cell instance $32501 r0 *1 173.43,158.34
X$32501 558 631 559 644 645 cell_1rw
* cell instance $32502 m0 *1 173.43,161.07
X$32502 558 632 559 644 645 cell_1rw
* cell instance $32503 r0 *1 173.43,161.07
X$32503 558 633 559 644 645 cell_1rw
* cell instance $32504 m0 *1 173.43,163.8
X$32504 558 634 559 644 645 cell_1rw
* cell instance $32505 m0 *1 173.43,166.53
X$32505 558 637 559 644 645 cell_1rw
* cell instance $32506 r0 *1 173.43,163.8
X$32506 558 635 559 644 645 cell_1rw
* cell instance $32507 m0 *1 173.43,169.26
X$32507 558 639 559 644 645 cell_1rw
* cell instance $32508 r0 *1 173.43,166.53
X$32508 558 636 559 644 645 cell_1rw
* cell instance $32509 m0 *1 173.43,171.99
X$32509 558 640 559 644 645 cell_1rw
* cell instance $32510 r0 *1 173.43,169.26
X$32510 558 638 559 644 645 cell_1rw
* cell instance $32511 m0 *1 173.43,174.72
X$32511 558 642 559 644 645 cell_1rw
* cell instance $32512 r0 *1 173.43,171.99
X$32512 558 641 559 644 645 cell_1rw
* cell instance $32513 r0 *1 173.43,174.72
X$32513 558 643 559 644 645 cell_1rw
* cell instance $32514 m0 *1 174.135,90.09
X$32514 560 581 561 644 645 cell_1rw
* cell instance $32515 r0 *1 174.135,90.09
X$32515 560 580 561 644 645 cell_1rw
* cell instance $32516 m0 *1 174.135,92.82
X$32516 560 583 561 644 645 cell_1rw
* cell instance $32517 r0 *1 174.135,92.82
X$32517 560 582 561 644 645 cell_1rw
* cell instance $32518 m0 *1 174.135,95.55
X$32518 560 584 561 644 645 cell_1rw
* cell instance $32519 r0 *1 174.135,95.55
X$32519 560 585 561 644 645 cell_1rw
* cell instance $32520 m0 *1 174.135,98.28
X$32520 560 586 561 644 645 cell_1rw
* cell instance $32521 r0 *1 174.135,98.28
X$32521 560 587 561 644 645 cell_1rw
* cell instance $32522 m0 *1 174.135,101.01
X$32522 560 588 561 644 645 cell_1rw
* cell instance $32523 r0 *1 174.135,101.01
X$32523 560 589 561 644 645 cell_1rw
* cell instance $32524 m0 *1 174.135,103.74
X$32524 560 590 561 644 645 cell_1rw
* cell instance $32525 r0 *1 174.135,103.74
X$32525 560 591 561 644 645 cell_1rw
* cell instance $32526 m0 *1 174.135,106.47
X$32526 560 593 561 644 645 cell_1rw
* cell instance $32527 m0 *1 174.135,109.2
X$32527 560 594 561 644 645 cell_1rw
* cell instance $32528 r0 *1 174.135,106.47
X$32528 560 592 561 644 645 cell_1rw
* cell instance $32529 r0 *1 174.135,109.2
X$32529 560 595 561 644 645 cell_1rw
* cell instance $32530 m0 *1 174.135,111.93
X$32530 560 597 561 644 645 cell_1rw
* cell instance $32531 r0 *1 174.135,111.93
X$32531 560 596 561 644 645 cell_1rw
* cell instance $32532 m0 *1 174.135,114.66
X$32532 560 598 561 644 645 cell_1rw
* cell instance $32533 m0 *1 174.135,117.39
X$32533 560 600 561 644 645 cell_1rw
* cell instance $32534 r0 *1 174.135,114.66
X$32534 560 599 561 644 645 cell_1rw
* cell instance $32535 r0 *1 174.135,117.39
X$32535 560 601 561 644 645 cell_1rw
* cell instance $32536 m0 *1 174.135,120.12
X$32536 560 602 561 644 645 cell_1rw
* cell instance $32537 r0 *1 174.135,120.12
X$32537 560 603 561 644 645 cell_1rw
* cell instance $32538 m0 *1 174.135,122.85
X$32538 560 604 561 644 645 cell_1rw
* cell instance $32539 r0 *1 174.135,122.85
X$32539 560 605 561 644 645 cell_1rw
* cell instance $32540 m0 *1 174.135,125.58
X$32540 560 606 561 644 645 cell_1rw
* cell instance $32541 r0 *1 174.135,125.58
X$32541 560 607 561 644 645 cell_1rw
* cell instance $32542 m0 *1 174.135,128.31
X$32542 560 609 561 644 645 cell_1rw
* cell instance $32543 r0 *1 174.135,128.31
X$32543 560 608 561 644 645 cell_1rw
* cell instance $32544 m0 *1 174.135,131.04
X$32544 560 610 561 644 645 cell_1rw
* cell instance $32545 r0 *1 174.135,131.04
X$32545 560 611 561 644 645 cell_1rw
* cell instance $32546 m0 *1 174.135,133.77
X$32546 560 612 561 644 645 cell_1rw
* cell instance $32547 r0 *1 174.135,133.77
X$32547 560 613 561 644 645 cell_1rw
* cell instance $32548 m0 *1 174.135,136.5
X$32548 560 615 561 644 645 cell_1rw
* cell instance $32549 r0 *1 174.135,136.5
X$32549 560 614 561 644 645 cell_1rw
* cell instance $32550 m0 *1 174.135,139.23
X$32550 560 617 561 644 645 cell_1rw
* cell instance $32551 r0 *1 174.135,139.23
X$32551 560 616 561 644 645 cell_1rw
* cell instance $32552 m0 *1 174.135,141.96
X$32552 560 618 561 644 645 cell_1rw
* cell instance $32553 m0 *1 174.135,144.69
X$32553 560 620 561 644 645 cell_1rw
* cell instance $32554 r0 *1 174.135,141.96
X$32554 560 619 561 644 645 cell_1rw
* cell instance $32555 r0 *1 174.135,144.69
X$32555 560 621 561 644 645 cell_1rw
* cell instance $32556 m0 *1 174.135,147.42
X$32556 560 622 561 644 645 cell_1rw
* cell instance $32557 r0 *1 174.135,147.42
X$32557 560 623 561 644 645 cell_1rw
* cell instance $32558 m0 *1 174.135,150.15
X$32558 560 624 561 644 645 cell_1rw
* cell instance $32559 m0 *1 174.135,152.88
X$32559 560 626 561 644 645 cell_1rw
* cell instance $32560 r0 *1 174.135,150.15
X$32560 560 625 561 644 645 cell_1rw
* cell instance $32561 m0 *1 174.135,155.61
X$32561 560 628 561 644 645 cell_1rw
* cell instance $32562 r0 *1 174.135,152.88
X$32562 560 627 561 644 645 cell_1rw
* cell instance $32563 m0 *1 174.135,158.34
X$32563 560 630 561 644 645 cell_1rw
* cell instance $32564 r0 *1 174.135,155.61
X$32564 560 629 561 644 645 cell_1rw
* cell instance $32565 m0 *1 174.135,161.07
X$32565 560 632 561 644 645 cell_1rw
* cell instance $32566 r0 *1 174.135,158.34
X$32566 560 631 561 644 645 cell_1rw
* cell instance $32567 r0 *1 174.135,161.07
X$32567 560 633 561 644 645 cell_1rw
* cell instance $32568 m0 *1 174.135,163.8
X$32568 560 634 561 644 645 cell_1rw
* cell instance $32569 m0 *1 174.135,166.53
X$32569 560 637 561 644 645 cell_1rw
* cell instance $32570 r0 *1 174.135,163.8
X$32570 560 635 561 644 645 cell_1rw
* cell instance $32571 r0 *1 174.135,166.53
X$32571 560 636 561 644 645 cell_1rw
* cell instance $32572 m0 *1 174.135,169.26
X$32572 560 639 561 644 645 cell_1rw
* cell instance $32573 r0 *1 174.135,169.26
X$32573 560 638 561 644 645 cell_1rw
* cell instance $32574 m0 *1 174.135,171.99
X$32574 560 640 561 644 645 cell_1rw
* cell instance $32575 r0 *1 174.135,171.99
X$32575 560 641 561 644 645 cell_1rw
* cell instance $32576 m0 *1 174.135,174.72
X$32576 560 642 561 644 645 cell_1rw
* cell instance $32577 r0 *1 174.135,174.72
X$32577 560 643 561 644 645 cell_1rw
* cell instance $32578 m0 *1 174.84,90.09
X$32578 562 581 563 644 645 cell_1rw
* cell instance $32579 r0 *1 174.84,90.09
X$32579 562 580 563 644 645 cell_1rw
* cell instance $32580 m0 *1 174.84,92.82
X$32580 562 583 563 644 645 cell_1rw
* cell instance $32581 m0 *1 174.84,95.55
X$32581 562 584 563 644 645 cell_1rw
* cell instance $32582 r0 *1 174.84,92.82
X$32582 562 582 563 644 645 cell_1rw
* cell instance $32583 r0 *1 174.84,95.55
X$32583 562 585 563 644 645 cell_1rw
* cell instance $32584 m0 *1 174.84,98.28
X$32584 562 586 563 644 645 cell_1rw
* cell instance $32585 m0 *1 174.84,101.01
X$32585 562 588 563 644 645 cell_1rw
* cell instance $32586 r0 *1 174.84,98.28
X$32586 562 587 563 644 645 cell_1rw
* cell instance $32587 r0 *1 174.84,101.01
X$32587 562 589 563 644 645 cell_1rw
* cell instance $32588 m0 *1 174.84,103.74
X$32588 562 590 563 644 645 cell_1rw
* cell instance $32589 m0 *1 174.84,106.47
X$32589 562 593 563 644 645 cell_1rw
* cell instance $32590 r0 *1 174.84,103.74
X$32590 562 591 563 644 645 cell_1rw
* cell instance $32591 r0 *1 174.84,106.47
X$32591 562 592 563 644 645 cell_1rw
* cell instance $32592 m0 *1 174.84,109.2
X$32592 562 594 563 644 645 cell_1rw
* cell instance $32593 m0 *1 174.84,111.93
X$32593 562 597 563 644 645 cell_1rw
* cell instance $32594 r0 *1 174.84,109.2
X$32594 562 595 563 644 645 cell_1rw
* cell instance $32595 r0 *1 174.84,111.93
X$32595 562 596 563 644 645 cell_1rw
* cell instance $32596 m0 *1 174.84,114.66
X$32596 562 598 563 644 645 cell_1rw
* cell instance $32597 r0 *1 174.84,114.66
X$32597 562 599 563 644 645 cell_1rw
* cell instance $32598 m0 *1 174.84,117.39
X$32598 562 600 563 644 645 cell_1rw
* cell instance $32599 r0 *1 174.84,117.39
X$32599 562 601 563 644 645 cell_1rw
* cell instance $32600 m0 *1 174.84,120.12
X$32600 562 602 563 644 645 cell_1rw
* cell instance $32601 m0 *1 174.84,122.85
X$32601 562 604 563 644 645 cell_1rw
* cell instance $32602 r0 *1 174.84,120.12
X$32602 562 603 563 644 645 cell_1rw
* cell instance $32603 r0 *1 174.84,122.85
X$32603 562 605 563 644 645 cell_1rw
* cell instance $32604 m0 *1 174.84,125.58
X$32604 562 606 563 644 645 cell_1rw
* cell instance $32605 r0 *1 174.84,125.58
X$32605 562 607 563 644 645 cell_1rw
* cell instance $32606 m0 *1 174.84,128.31
X$32606 562 609 563 644 645 cell_1rw
* cell instance $32607 r0 *1 174.84,128.31
X$32607 562 608 563 644 645 cell_1rw
* cell instance $32608 m0 *1 174.84,131.04
X$32608 562 610 563 644 645 cell_1rw
* cell instance $32609 r0 *1 174.84,131.04
X$32609 562 611 563 644 645 cell_1rw
* cell instance $32610 m0 *1 174.84,133.77
X$32610 562 612 563 644 645 cell_1rw
* cell instance $32611 m0 *1 174.84,136.5
X$32611 562 615 563 644 645 cell_1rw
* cell instance $32612 r0 *1 174.84,133.77
X$32612 562 613 563 644 645 cell_1rw
* cell instance $32613 m0 *1 174.84,139.23
X$32613 562 617 563 644 645 cell_1rw
* cell instance $32614 r0 *1 174.84,136.5
X$32614 562 614 563 644 645 cell_1rw
* cell instance $32615 r0 *1 174.84,139.23
X$32615 562 616 563 644 645 cell_1rw
* cell instance $32616 m0 *1 174.84,141.96
X$32616 562 618 563 644 645 cell_1rw
* cell instance $32617 r0 *1 174.84,141.96
X$32617 562 619 563 644 645 cell_1rw
* cell instance $32618 m0 *1 174.84,144.69
X$32618 562 620 563 644 645 cell_1rw
* cell instance $32619 r0 *1 174.84,144.69
X$32619 562 621 563 644 645 cell_1rw
* cell instance $32620 m0 *1 174.84,147.42
X$32620 562 622 563 644 645 cell_1rw
* cell instance $32621 r0 *1 174.84,147.42
X$32621 562 623 563 644 645 cell_1rw
* cell instance $32622 m0 *1 174.84,150.15
X$32622 562 624 563 644 645 cell_1rw
* cell instance $32623 r0 *1 174.84,150.15
X$32623 562 625 563 644 645 cell_1rw
* cell instance $32624 m0 *1 174.84,152.88
X$32624 562 626 563 644 645 cell_1rw
* cell instance $32625 r0 *1 174.84,152.88
X$32625 562 627 563 644 645 cell_1rw
* cell instance $32626 m0 *1 174.84,155.61
X$32626 562 628 563 644 645 cell_1rw
* cell instance $32627 r0 *1 174.84,155.61
X$32627 562 629 563 644 645 cell_1rw
* cell instance $32628 m0 *1 174.84,158.34
X$32628 562 630 563 644 645 cell_1rw
* cell instance $32629 r0 *1 174.84,158.34
X$32629 562 631 563 644 645 cell_1rw
* cell instance $32630 m0 *1 174.84,161.07
X$32630 562 632 563 644 645 cell_1rw
* cell instance $32631 m0 *1 174.84,163.8
X$32631 562 634 563 644 645 cell_1rw
* cell instance $32632 r0 *1 174.84,161.07
X$32632 562 633 563 644 645 cell_1rw
* cell instance $32633 r0 *1 174.84,163.8
X$32633 562 635 563 644 645 cell_1rw
* cell instance $32634 m0 *1 174.84,166.53
X$32634 562 637 563 644 645 cell_1rw
* cell instance $32635 r0 *1 174.84,166.53
X$32635 562 636 563 644 645 cell_1rw
* cell instance $32636 m0 *1 174.84,169.26
X$32636 562 639 563 644 645 cell_1rw
* cell instance $32637 r0 *1 174.84,169.26
X$32637 562 638 563 644 645 cell_1rw
* cell instance $32638 m0 *1 174.84,171.99
X$32638 562 640 563 644 645 cell_1rw
* cell instance $32639 m0 *1 174.84,174.72
X$32639 562 642 563 644 645 cell_1rw
* cell instance $32640 r0 *1 174.84,171.99
X$32640 562 641 563 644 645 cell_1rw
* cell instance $32641 r0 *1 174.84,174.72
X$32641 562 643 563 644 645 cell_1rw
* cell instance $32642 m0 *1 175.545,90.09
X$32642 564 581 565 644 645 cell_1rw
* cell instance $32643 r0 *1 175.545,90.09
X$32643 564 580 565 644 645 cell_1rw
* cell instance $32644 m0 *1 175.545,92.82
X$32644 564 583 565 644 645 cell_1rw
* cell instance $32645 r0 *1 175.545,92.82
X$32645 564 582 565 644 645 cell_1rw
* cell instance $32646 m0 *1 175.545,95.55
X$32646 564 584 565 644 645 cell_1rw
* cell instance $32647 m0 *1 175.545,98.28
X$32647 564 586 565 644 645 cell_1rw
* cell instance $32648 r0 *1 175.545,95.55
X$32648 564 585 565 644 645 cell_1rw
* cell instance $32649 m0 *1 175.545,101.01
X$32649 564 588 565 644 645 cell_1rw
* cell instance $32650 r0 *1 175.545,98.28
X$32650 564 587 565 644 645 cell_1rw
* cell instance $32651 r0 *1 175.545,101.01
X$32651 564 589 565 644 645 cell_1rw
* cell instance $32652 m0 *1 175.545,103.74
X$32652 564 590 565 644 645 cell_1rw
* cell instance $32653 r0 *1 175.545,103.74
X$32653 564 591 565 644 645 cell_1rw
* cell instance $32654 m0 *1 175.545,106.47
X$32654 564 593 565 644 645 cell_1rw
* cell instance $32655 m0 *1 175.545,109.2
X$32655 564 594 565 644 645 cell_1rw
* cell instance $32656 r0 *1 175.545,106.47
X$32656 564 592 565 644 645 cell_1rw
* cell instance $32657 r0 *1 175.545,109.2
X$32657 564 595 565 644 645 cell_1rw
* cell instance $32658 m0 *1 175.545,111.93
X$32658 564 597 565 644 645 cell_1rw
* cell instance $32659 r0 *1 175.545,111.93
X$32659 564 596 565 644 645 cell_1rw
* cell instance $32660 m0 *1 175.545,114.66
X$32660 564 598 565 644 645 cell_1rw
* cell instance $32661 r0 *1 175.545,114.66
X$32661 564 599 565 644 645 cell_1rw
* cell instance $32662 m0 *1 175.545,117.39
X$32662 564 600 565 644 645 cell_1rw
* cell instance $32663 r0 *1 175.545,117.39
X$32663 564 601 565 644 645 cell_1rw
* cell instance $32664 m0 *1 175.545,120.12
X$32664 564 602 565 644 645 cell_1rw
* cell instance $32665 r0 *1 175.545,120.12
X$32665 564 603 565 644 645 cell_1rw
* cell instance $32666 m0 *1 175.545,122.85
X$32666 564 604 565 644 645 cell_1rw
* cell instance $32667 r0 *1 175.545,122.85
X$32667 564 605 565 644 645 cell_1rw
* cell instance $32668 m0 *1 175.545,125.58
X$32668 564 606 565 644 645 cell_1rw
* cell instance $32669 r0 *1 175.545,125.58
X$32669 564 607 565 644 645 cell_1rw
* cell instance $32670 m0 *1 175.545,128.31
X$32670 564 609 565 644 645 cell_1rw
* cell instance $32671 r0 *1 175.545,128.31
X$32671 564 608 565 644 645 cell_1rw
* cell instance $32672 m0 *1 175.545,131.04
X$32672 564 610 565 644 645 cell_1rw
* cell instance $32673 m0 *1 175.545,133.77
X$32673 564 612 565 644 645 cell_1rw
* cell instance $32674 r0 *1 175.545,131.04
X$32674 564 611 565 644 645 cell_1rw
* cell instance $32675 r0 *1 175.545,133.77
X$32675 564 613 565 644 645 cell_1rw
* cell instance $32676 m0 *1 175.545,136.5
X$32676 564 615 565 644 645 cell_1rw
* cell instance $32677 r0 *1 175.545,136.5
X$32677 564 614 565 644 645 cell_1rw
* cell instance $32678 m0 *1 175.545,139.23
X$32678 564 617 565 644 645 cell_1rw
* cell instance $32679 r0 *1 175.545,139.23
X$32679 564 616 565 644 645 cell_1rw
* cell instance $32680 m0 *1 175.545,141.96
X$32680 564 618 565 644 645 cell_1rw
* cell instance $32681 r0 *1 175.545,141.96
X$32681 564 619 565 644 645 cell_1rw
* cell instance $32682 m0 *1 175.545,144.69
X$32682 564 620 565 644 645 cell_1rw
* cell instance $32683 m0 *1 175.545,147.42
X$32683 564 622 565 644 645 cell_1rw
* cell instance $32684 r0 *1 175.545,144.69
X$32684 564 621 565 644 645 cell_1rw
* cell instance $32685 r0 *1 175.545,147.42
X$32685 564 623 565 644 645 cell_1rw
* cell instance $32686 m0 *1 175.545,150.15
X$32686 564 624 565 644 645 cell_1rw
* cell instance $32687 m0 *1 175.545,152.88
X$32687 564 626 565 644 645 cell_1rw
* cell instance $32688 r0 *1 175.545,150.15
X$32688 564 625 565 644 645 cell_1rw
* cell instance $32689 r0 *1 175.545,152.88
X$32689 564 627 565 644 645 cell_1rw
* cell instance $32690 m0 *1 175.545,155.61
X$32690 564 628 565 644 645 cell_1rw
* cell instance $32691 r0 *1 175.545,155.61
X$32691 564 629 565 644 645 cell_1rw
* cell instance $32692 m0 *1 175.545,158.34
X$32692 564 630 565 644 645 cell_1rw
* cell instance $32693 m0 *1 175.545,161.07
X$32693 564 632 565 644 645 cell_1rw
* cell instance $32694 r0 *1 175.545,158.34
X$32694 564 631 565 644 645 cell_1rw
* cell instance $32695 r0 *1 175.545,161.07
X$32695 564 633 565 644 645 cell_1rw
* cell instance $32696 m0 *1 175.545,163.8
X$32696 564 634 565 644 645 cell_1rw
* cell instance $32697 r0 *1 175.545,163.8
X$32697 564 635 565 644 645 cell_1rw
* cell instance $32698 m0 *1 175.545,166.53
X$32698 564 637 565 644 645 cell_1rw
* cell instance $32699 r0 *1 175.545,166.53
X$32699 564 636 565 644 645 cell_1rw
* cell instance $32700 m0 *1 175.545,169.26
X$32700 564 639 565 644 645 cell_1rw
* cell instance $32701 r0 *1 175.545,169.26
X$32701 564 638 565 644 645 cell_1rw
* cell instance $32702 m0 *1 175.545,171.99
X$32702 564 640 565 644 645 cell_1rw
* cell instance $32703 r0 *1 175.545,171.99
X$32703 564 641 565 644 645 cell_1rw
* cell instance $32704 m0 *1 175.545,174.72
X$32704 564 642 565 644 645 cell_1rw
* cell instance $32705 r0 *1 175.545,174.72
X$32705 564 643 565 644 645 cell_1rw
* cell instance $32706 m0 *1 176.25,90.09
X$32706 566 581 567 644 645 cell_1rw
* cell instance $32707 r0 *1 176.25,90.09
X$32707 566 580 567 644 645 cell_1rw
* cell instance $32708 m0 *1 176.25,92.82
X$32708 566 583 567 644 645 cell_1rw
* cell instance $32709 r0 *1 176.25,92.82
X$32709 566 582 567 644 645 cell_1rw
* cell instance $32710 m0 *1 176.25,95.55
X$32710 566 584 567 644 645 cell_1rw
* cell instance $32711 r0 *1 176.25,95.55
X$32711 566 585 567 644 645 cell_1rw
* cell instance $32712 m0 *1 176.25,98.28
X$32712 566 586 567 644 645 cell_1rw
* cell instance $32713 r0 *1 176.25,98.28
X$32713 566 587 567 644 645 cell_1rw
* cell instance $32714 m0 *1 176.25,101.01
X$32714 566 588 567 644 645 cell_1rw
* cell instance $32715 r0 *1 176.25,101.01
X$32715 566 589 567 644 645 cell_1rw
* cell instance $32716 m0 *1 176.25,103.74
X$32716 566 590 567 644 645 cell_1rw
* cell instance $32717 m0 *1 176.25,106.47
X$32717 566 593 567 644 645 cell_1rw
* cell instance $32718 r0 *1 176.25,103.74
X$32718 566 591 567 644 645 cell_1rw
* cell instance $32719 r0 *1 176.25,106.47
X$32719 566 592 567 644 645 cell_1rw
* cell instance $32720 m0 *1 176.25,109.2
X$32720 566 594 567 644 645 cell_1rw
* cell instance $32721 r0 *1 176.25,109.2
X$32721 566 595 567 644 645 cell_1rw
* cell instance $32722 m0 *1 176.25,111.93
X$32722 566 597 567 644 645 cell_1rw
* cell instance $32723 r0 *1 176.25,111.93
X$32723 566 596 567 644 645 cell_1rw
* cell instance $32724 m0 *1 176.25,114.66
X$32724 566 598 567 644 645 cell_1rw
* cell instance $32725 r0 *1 176.25,114.66
X$32725 566 599 567 644 645 cell_1rw
* cell instance $32726 m0 *1 176.25,117.39
X$32726 566 600 567 644 645 cell_1rw
* cell instance $32727 r0 *1 176.25,117.39
X$32727 566 601 567 644 645 cell_1rw
* cell instance $32728 m0 *1 176.25,120.12
X$32728 566 602 567 644 645 cell_1rw
* cell instance $32729 r0 *1 176.25,120.12
X$32729 566 603 567 644 645 cell_1rw
* cell instance $32730 m0 *1 176.25,122.85
X$32730 566 604 567 644 645 cell_1rw
* cell instance $32731 r0 *1 176.25,122.85
X$32731 566 605 567 644 645 cell_1rw
* cell instance $32732 m0 *1 176.25,125.58
X$32732 566 606 567 644 645 cell_1rw
* cell instance $32733 r0 *1 176.25,125.58
X$32733 566 607 567 644 645 cell_1rw
* cell instance $32734 m0 *1 176.25,128.31
X$32734 566 609 567 644 645 cell_1rw
* cell instance $32735 m0 *1 176.25,131.04
X$32735 566 610 567 644 645 cell_1rw
* cell instance $32736 r0 *1 176.25,128.31
X$32736 566 608 567 644 645 cell_1rw
* cell instance $32737 r0 *1 176.25,131.04
X$32737 566 611 567 644 645 cell_1rw
* cell instance $32738 m0 *1 176.25,133.77
X$32738 566 612 567 644 645 cell_1rw
* cell instance $32739 r0 *1 176.25,133.77
X$32739 566 613 567 644 645 cell_1rw
* cell instance $32740 m0 *1 176.25,136.5
X$32740 566 615 567 644 645 cell_1rw
* cell instance $32741 r0 *1 176.25,136.5
X$32741 566 614 567 644 645 cell_1rw
* cell instance $32742 m0 *1 176.25,139.23
X$32742 566 617 567 644 645 cell_1rw
* cell instance $32743 r0 *1 176.25,139.23
X$32743 566 616 567 644 645 cell_1rw
* cell instance $32744 m0 *1 176.25,141.96
X$32744 566 618 567 644 645 cell_1rw
* cell instance $32745 r0 *1 176.25,141.96
X$32745 566 619 567 644 645 cell_1rw
* cell instance $32746 m0 *1 176.25,144.69
X$32746 566 620 567 644 645 cell_1rw
* cell instance $32747 m0 *1 176.25,147.42
X$32747 566 622 567 644 645 cell_1rw
* cell instance $32748 r0 *1 176.25,144.69
X$32748 566 621 567 644 645 cell_1rw
* cell instance $32749 r0 *1 176.25,147.42
X$32749 566 623 567 644 645 cell_1rw
* cell instance $32750 m0 *1 176.25,150.15
X$32750 566 624 567 644 645 cell_1rw
* cell instance $32751 r0 *1 176.25,150.15
X$32751 566 625 567 644 645 cell_1rw
* cell instance $32752 m0 *1 176.25,152.88
X$32752 566 626 567 644 645 cell_1rw
* cell instance $32753 r0 *1 176.25,152.88
X$32753 566 627 567 644 645 cell_1rw
* cell instance $32754 m0 *1 176.25,155.61
X$32754 566 628 567 644 645 cell_1rw
* cell instance $32755 r0 *1 176.25,155.61
X$32755 566 629 567 644 645 cell_1rw
* cell instance $32756 m0 *1 176.25,158.34
X$32756 566 630 567 644 645 cell_1rw
* cell instance $32757 m0 *1 176.25,161.07
X$32757 566 632 567 644 645 cell_1rw
* cell instance $32758 r0 *1 176.25,158.34
X$32758 566 631 567 644 645 cell_1rw
* cell instance $32759 r0 *1 176.25,161.07
X$32759 566 633 567 644 645 cell_1rw
* cell instance $32760 m0 *1 176.25,163.8
X$32760 566 634 567 644 645 cell_1rw
* cell instance $32761 r0 *1 176.25,163.8
X$32761 566 635 567 644 645 cell_1rw
* cell instance $32762 m0 *1 176.25,166.53
X$32762 566 637 567 644 645 cell_1rw
* cell instance $32763 r0 *1 176.25,166.53
X$32763 566 636 567 644 645 cell_1rw
* cell instance $32764 m0 *1 176.25,169.26
X$32764 566 639 567 644 645 cell_1rw
* cell instance $32765 r0 *1 176.25,169.26
X$32765 566 638 567 644 645 cell_1rw
* cell instance $32766 m0 *1 176.25,171.99
X$32766 566 640 567 644 645 cell_1rw
* cell instance $32767 m0 *1 176.25,174.72
X$32767 566 642 567 644 645 cell_1rw
* cell instance $32768 r0 *1 176.25,171.99
X$32768 566 641 567 644 645 cell_1rw
* cell instance $32769 r0 *1 176.25,174.72
X$32769 566 643 567 644 645 cell_1rw
* cell instance $32770 m0 *1 176.955,90.09
X$32770 568 581 569 644 645 cell_1rw
* cell instance $32771 r0 *1 176.955,90.09
X$32771 568 580 569 644 645 cell_1rw
* cell instance $32772 m0 *1 176.955,92.82
X$32772 568 583 569 644 645 cell_1rw
* cell instance $32773 m0 *1 176.955,95.55
X$32773 568 584 569 644 645 cell_1rw
* cell instance $32774 r0 *1 176.955,92.82
X$32774 568 582 569 644 645 cell_1rw
* cell instance $32775 r0 *1 176.955,95.55
X$32775 568 585 569 644 645 cell_1rw
* cell instance $32776 m0 *1 176.955,98.28
X$32776 568 586 569 644 645 cell_1rw
* cell instance $32777 r0 *1 176.955,98.28
X$32777 568 587 569 644 645 cell_1rw
* cell instance $32778 m0 *1 176.955,101.01
X$32778 568 588 569 644 645 cell_1rw
* cell instance $32779 r0 *1 176.955,101.01
X$32779 568 589 569 644 645 cell_1rw
* cell instance $32780 m0 *1 176.955,103.74
X$32780 568 590 569 644 645 cell_1rw
* cell instance $32781 r0 *1 176.955,103.74
X$32781 568 591 569 644 645 cell_1rw
* cell instance $32782 m0 *1 176.955,106.47
X$32782 568 593 569 644 645 cell_1rw
* cell instance $32783 m0 *1 176.955,109.2
X$32783 568 594 569 644 645 cell_1rw
* cell instance $32784 r0 *1 176.955,106.47
X$32784 568 592 569 644 645 cell_1rw
* cell instance $32785 r0 *1 176.955,109.2
X$32785 568 595 569 644 645 cell_1rw
* cell instance $32786 m0 *1 176.955,111.93
X$32786 568 597 569 644 645 cell_1rw
* cell instance $32787 r0 *1 176.955,111.93
X$32787 568 596 569 644 645 cell_1rw
* cell instance $32788 m0 *1 176.955,114.66
X$32788 568 598 569 644 645 cell_1rw
* cell instance $32789 r0 *1 176.955,114.66
X$32789 568 599 569 644 645 cell_1rw
* cell instance $32790 m0 *1 176.955,117.39
X$32790 568 600 569 644 645 cell_1rw
* cell instance $32791 r0 *1 176.955,117.39
X$32791 568 601 569 644 645 cell_1rw
* cell instance $32792 m0 *1 176.955,120.12
X$32792 568 602 569 644 645 cell_1rw
* cell instance $32793 m0 *1 176.955,122.85
X$32793 568 604 569 644 645 cell_1rw
* cell instance $32794 r0 *1 176.955,120.12
X$32794 568 603 569 644 645 cell_1rw
* cell instance $32795 r0 *1 176.955,122.85
X$32795 568 605 569 644 645 cell_1rw
* cell instance $32796 m0 *1 176.955,125.58
X$32796 568 606 569 644 645 cell_1rw
* cell instance $32797 r0 *1 176.955,125.58
X$32797 568 607 569 644 645 cell_1rw
* cell instance $32798 m0 *1 176.955,128.31
X$32798 568 609 569 644 645 cell_1rw
* cell instance $32799 r0 *1 176.955,128.31
X$32799 568 608 569 644 645 cell_1rw
* cell instance $32800 m0 *1 176.955,131.04
X$32800 568 610 569 644 645 cell_1rw
* cell instance $32801 m0 *1 176.955,133.77
X$32801 568 612 569 644 645 cell_1rw
* cell instance $32802 r0 *1 176.955,131.04
X$32802 568 611 569 644 645 cell_1rw
* cell instance $32803 r0 *1 176.955,133.77
X$32803 568 613 569 644 645 cell_1rw
* cell instance $32804 m0 *1 176.955,136.5
X$32804 568 615 569 644 645 cell_1rw
* cell instance $32805 r0 *1 176.955,136.5
X$32805 568 614 569 644 645 cell_1rw
* cell instance $32806 m0 *1 176.955,139.23
X$32806 568 617 569 644 645 cell_1rw
* cell instance $32807 m0 *1 176.955,141.96
X$32807 568 618 569 644 645 cell_1rw
* cell instance $32808 r0 *1 176.955,139.23
X$32808 568 616 569 644 645 cell_1rw
* cell instance $32809 r0 *1 176.955,141.96
X$32809 568 619 569 644 645 cell_1rw
* cell instance $32810 m0 *1 176.955,144.69
X$32810 568 620 569 644 645 cell_1rw
* cell instance $32811 r0 *1 176.955,144.69
X$32811 568 621 569 644 645 cell_1rw
* cell instance $32812 m0 *1 176.955,147.42
X$32812 568 622 569 644 645 cell_1rw
* cell instance $32813 r0 *1 176.955,147.42
X$32813 568 623 569 644 645 cell_1rw
* cell instance $32814 m0 *1 176.955,150.15
X$32814 568 624 569 644 645 cell_1rw
* cell instance $32815 r0 *1 176.955,150.15
X$32815 568 625 569 644 645 cell_1rw
* cell instance $32816 m0 *1 176.955,152.88
X$32816 568 626 569 644 645 cell_1rw
* cell instance $32817 r0 *1 176.955,152.88
X$32817 568 627 569 644 645 cell_1rw
* cell instance $32818 m0 *1 176.955,155.61
X$32818 568 628 569 644 645 cell_1rw
* cell instance $32819 r0 *1 176.955,155.61
X$32819 568 629 569 644 645 cell_1rw
* cell instance $32820 m0 *1 176.955,158.34
X$32820 568 630 569 644 645 cell_1rw
* cell instance $32821 r0 *1 176.955,158.34
X$32821 568 631 569 644 645 cell_1rw
* cell instance $32822 m0 *1 176.955,161.07
X$32822 568 632 569 644 645 cell_1rw
* cell instance $32823 r0 *1 176.955,161.07
X$32823 568 633 569 644 645 cell_1rw
* cell instance $32824 m0 *1 176.955,163.8
X$32824 568 634 569 644 645 cell_1rw
* cell instance $32825 r0 *1 176.955,163.8
X$32825 568 635 569 644 645 cell_1rw
* cell instance $32826 m0 *1 176.955,166.53
X$32826 568 637 569 644 645 cell_1rw
* cell instance $32827 r0 *1 176.955,166.53
X$32827 568 636 569 644 645 cell_1rw
* cell instance $32828 m0 *1 176.955,169.26
X$32828 568 639 569 644 645 cell_1rw
* cell instance $32829 r0 *1 176.955,169.26
X$32829 568 638 569 644 645 cell_1rw
* cell instance $32830 m0 *1 176.955,171.99
X$32830 568 640 569 644 645 cell_1rw
* cell instance $32831 r0 *1 176.955,171.99
X$32831 568 641 569 644 645 cell_1rw
* cell instance $32832 m0 *1 176.955,174.72
X$32832 568 642 569 644 645 cell_1rw
* cell instance $32833 r0 *1 176.955,174.72
X$32833 568 643 569 644 645 cell_1rw
* cell instance $32834 m0 *1 177.66,90.09
X$32834 570 581 571 644 645 cell_1rw
* cell instance $32835 m0 *1 177.66,92.82
X$32835 570 583 571 644 645 cell_1rw
* cell instance $32836 r0 *1 177.66,90.09
X$32836 570 580 571 644 645 cell_1rw
* cell instance $32837 m0 *1 177.66,95.55
X$32837 570 584 571 644 645 cell_1rw
* cell instance $32838 r0 *1 177.66,92.82
X$32838 570 582 571 644 645 cell_1rw
* cell instance $32839 r0 *1 177.66,95.55
X$32839 570 585 571 644 645 cell_1rw
* cell instance $32840 m0 *1 177.66,98.28
X$32840 570 586 571 644 645 cell_1rw
* cell instance $32841 r0 *1 177.66,98.28
X$32841 570 587 571 644 645 cell_1rw
* cell instance $32842 m0 *1 177.66,101.01
X$32842 570 588 571 644 645 cell_1rw
* cell instance $32843 r0 *1 177.66,101.01
X$32843 570 589 571 644 645 cell_1rw
* cell instance $32844 m0 *1 177.66,103.74
X$32844 570 590 571 644 645 cell_1rw
* cell instance $32845 r0 *1 177.66,103.74
X$32845 570 591 571 644 645 cell_1rw
* cell instance $32846 m0 *1 177.66,106.47
X$32846 570 593 571 644 645 cell_1rw
* cell instance $32847 m0 *1 177.66,109.2
X$32847 570 594 571 644 645 cell_1rw
* cell instance $32848 r0 *1 177.66,106.47
X$32848 570 592 571 644 645 cell_1rw
* cell instance $32849 r0 *1 177.66,109.2
X$32849 570 595 571 644 645 cell_1rw
* cell instance $32850 m0 *1 177.66,111.93
X$32850 570 597 571 644 645 cell_1rw
* cell instance $32851 r0 *1 177.66,111.93
X$32851 570 596 571 644 645 cell_1rw
* cell instance $32852 m0 *1 177.66,114.66
X$32852 570 598 571 644 645 cell_1rw
* cell instance $32853 r0 *1 177.66,114.66
X$32853 570 599 571 644 645 cell_1rw
* cell instance $32854 m0 *1 177.66,117.39
X$32854 570 600 571 644 645 cell_1rw
* cell instance $32855 m0 *1 177.66,120.12
X$32855 570 602 571 644 645 cell_1rw
* cell instance $32856 r0 *1 177.66,117.39
X$32856 570 601 571 644 645 cell_1rw
* cell instance $32857 r0 *1 177.66,120.12
X$32857 570 603 571 644 645 cell_1rw
* cell instance $32858 m0 *1 177.66,122.85
X$32858 570 604 571 644 645 cell_1rw
* cell instance $32859 r0 *1 177.66,122.85
X$32859 570 605 571 644 645 cell_1rw
* cell instance $32860 m0 *1 177.66,125.58
X$32860 570 606 571 644 645 cell_1rw
* cell instance $32861 r0 *1 177.66,125.58
X$32861 570 607 571 644 645 cell_1rw
* cell instance $32862 m0 *1 177.66,128.31
X$32862 570 609 571 644 645 cell_1rw
* cell instance $32863 r0 *1 177.66,128.31
X$32863 570 608 571 644 645 cell_1rw
* cell instance $32864 m0 *1 177.66,131.04
X$32864 570 610 571 644 645 cell_1rw
* cell instance $32865 r0 *1 177.66,131.04
X$32865 570 611 571 644 645 cell_1rw
* cell instance $32866 m0 *1 177.66,133.77
X$32866 570 612 571 644 645 cell_1rw
* cell instance $32867 r0 *1 177.66,133.77
X$32867 570 613 571 644 645 cell_1rw
* cell instance $32868 m0 *1 177.66,136.5
X$32868 570 615 571 644 645 cell_1rw
* cell instance $32869 r0 *1 177.66,136.5
X$32869 570 614 571 644 645 cell_1rw
* cell instance $32870 m0 *1 177.66,139.23
X$32870 570 617 571 644 645 cell_1rw
* cell instance $32871 r0 *1 177.66,139.23
X$32871 570 616 571 644 645 cell_1rw
* cell instance $32872 m0 *1 177.66,141.96
X$32872 570 618 571 644 645 cell_1rw
* cell instance $32873 r0 *1 177.66,141.96
X$32873 570 619 571 644 645 cell_1rw
* cell instance $32874 m0 *1 177.66,144.69
X$32874 570 620 571 644 645 cell_1rw
* cell instance $32875 r0 *1 177.66,144.69
X$32875 570 621 571 644 645 cell_1rw
* cell instance $32876 m0 *1 177.66,147.42
X$32876 570 622 571 644 645 cell_1rw
* cell instance $32877 r0 *1 177.66,147.42
X$32877 570 623 571 644 645 cell_1rw
* cell instance $32878 m0 *1 177.66,150.15
X$32878 570 624 571 644 645 cell_1rw
* cell instance $32879 r0 *1 177.66,150.15
X$32879 570 625 571 644 645 cell_1rw
* cell instance $32880 m0 *1 177.66,152.88
X$32880 570 626 571 644 645 cell_1rw
* cell instance $32881 r0 *1 177.66,152.88
X$32881 570 627 571 644 645 cell_1rw
* cell instance $32882 m0 *1 177.66,155.61
X$32882 570 628 571 644 645 cell_1rw
* cell instance $32883 r0 *1 177.66,155.61
X$32883 570 629 571 644 645 cell_1rw
* cell instance $32884 m0 *1 177.66,158.34
X$32884 570 630 571 644 645 cell_1rw
* cell instance $32885 r0 *1 177.66,158.34
X$32885 570 631 571 644 645 cell_1rw
* cell instance $32886 m0 *1 177.66,161.07
X$32886 570 632 571 644 645 cell_1rw
* cell instance $32887 m0 *1 177.66,163.8
X$32887 570 634 571 644 645 cell_1rw
* cell instance $32888 r0 *1 177.66,161.07
X$32888 570 633 571 644 645 cell_1rw
* cell instance $32889 r0 *1 177.66,163.8
X$32889 570 635 571 644 645 cell_1rw
* cell instance $32890 m0 *1 177.66,166.53
X$32890 570 637 571 644 645 cell_1rw
* cell instance $32891 r0 *1 177.66,166.53
X$32891 570 636 571 644 645 cell_1rw
* cell instance $32892 m0 *1 177.66,169.26
X$32892 570 639 571 644 645 cell_1rw
* cell instance $32893 r0 *1 177.66,169.26
X$32893 570 638 571 644 645 cell_1rw
* cell instance $32894 m0 *1 177.66,171.99
X$32894 570 640 571 644 645 cell_1rw
* cell instance $32895 r0 *1 177.66,171.99
X$32895 570 641 571 644 645 cell_1rw
* cell instance $32896 m0 *1 177.66,174.72
X$32896 570 642 571 644 645 cell_1rw
* cell instance $32897 r0 *1 177.66,174.72
X$32897 570 643 571 644 645 cell_1rw
* cell instance $32898 m0 *1 178.365,90.09
X$32898 572 581 573 644 645 cell_1rw
* cell instance $32899 m0 *1 178.365,92.82
X$32899 572 583 573 644 645 cell_1rw
* cell instance $32900 r0 *1 178.365,90.09
X$32900 572 580 573 644 645 cell_1rw
* cell instance $32901 r0 *1 178.365,92.82
X$32901 572 582 573 644 645 cell_1rw
* cell instance $32902 m0 *1 178.365,95.55
X$32902 572 584 573 644 645 cell_1rw
* cell instance $32903 m0 *1 178.365,98.28
X$32903 572 586 573 644 645 cell_1rw
* cell instance $32904 r0 *1 178.365,95.55
X$32904 572 585 573 644 645 cell_1rw
* cell instance $32905 r0 *1 178.365,98.28
X$32905 572 587 573 644 645 cell_1rw
* cell instance $32906 m0 *1 178.365,101.01
X$32906 572 588 573 644 645 cell_1rw
* cell instance $32907 m0 *1 178.365,103.74
X$32907 572 590 573 644 645 cell_1rw
* cell instance $32908 r0 *1 178.365,101.01
X$32908 572 589 573 644 645 cell_1rw
* cell instance $32909 r0 *1 178.365,103.74
X$32909 572 591 573 644 645 cell_1rw
* cell instance $32910 m0 *1 178.365,106.47
X$32910 572 593 573 644 645 cell_1rw
* cell instance $32911 r0 *1 178.365,106.47
X$32911 572 592 573 644 645 cell_1rw
* cell instance $32912 m0 *1 178.365,109.2
X$32912 572 594 573 644 645 cell_1rw
* cell instance $32913 r0 *1 178.365,109.2
X$32913 572 595 573 644 645 cell_1rw
* cell instance $32914 m0 *1 178.365,111.93
X$32914 572 597 573 644 645 cell_1rw
* cell instance $32915 r0 *1 178.365,111.93
X$32915 572 596 573 644 645 cell_1rw
* cell instance $32916 m0 *1 178.365,114.66
X$32916 572 598 573 644 645 cell_1rw
* cell instance $32917 r0 *1 178.365,114.66
X$32917 572 599 573 644 645 cell_1rw
* cell instance $32918 m0 *1 178.365,117.39
X$32918 572 600 573 644 645 cell_1rw
* cell instance $32919 r0 *1 178.365,117.39
X$32919 572 601 573 644 645 cell_1rw
* cell instance $32920 m0 *1 178.365,120.12
X$32920 572 602 573 644 645 cell_1rw
* cell instance $32921 r0 *1 178.365,120.12
X$32921 572 603 573 644 645 cell_1rw
* cell instance $32922 m0 *1 178.365,122.85
X$32922 572 604 573 644 645 cell_1rw
* cell instance $32923 r0 *1 178.365,122.85
X$32923 572 605 573 644 645 cell_1rw
* cell instance $32924 m0 *1 178.365,125.58
X$32924 572 606 573 644 645 cell_1rw
* cell instance $32925 r0 *1 178.365,125.58
X$32925 572 607 573 644 645 cell_1rw
* cell instance $32926 m0 *1 178.365,128.31
X$32926 572 609 573 644 645 cell_1rw
* cell instance $32927 r0 *1 178.365,128.31
X$32927 572 608 573 644 645 cell_1rw
* cell instance $32928 m0 *1 178.365,131.04
X$32928 572 610 573 644 645 cell_1rw
* cell instance $32929 m0 *1 178.365,133.77
X$32929 572 612 573 644 645 cell_1rw
* cell instance $32930 r0 *1 178.365,131.04
X$32930 572 611 573 644 645 cell_1rw
* cell instance $32931 r0 *1 178.365,133.77
X$32931 572 613 573 644 645 cell_1rw
* cell instance $32932 m0 *1 178.365,136.5
X$32932 572 615 573 644 645 cell_1rw
* cell instance $32933 m0 *1 178.365,139.23
X$32933 572 617 573 644 645 cell_1rw
* cell instance $32934 r0 *1 178.365,136.5
X$32934 572 614 573 644 645 cell_1rw
* cell instance $32935 r0 *1 178.365,139.23
X$32935 572 616 573 644 645 cell_1rw
* cell instance $32936 m0 *1 178.365,141.96
X$32936 572 618 573 644 645 cell_1rw
* cell instance $32937 r0 *1 178.365,141.96
X$32937 572 619 573 644 645 cell_1rw
* cell instance $32938 m0 *1 178.365,144.69
X$32938 572 620 573 644 645 cell_1rw
* cell instance $32939 r0 *1 178.365,144.69
X$32939 572 621 573 644 645 cell_1rw
* cell instance $32940 m0 *1 178.365,147.42
X$32940 572 622 573 644 645 cell_1rw
* cell instance $32941 r0 *1 178.365,147.42
X$32941 572 623 573 644 645 cell_1rw
* cell instance $32942 m0 *1 178.365,150.15
X$32942 572 624 573 644 645 cell_1rw
* cell instance $32943 r0 *1 178.365,150.15
X$32943 572 625 573 644 645 cell_1rw
* cell instance $32944 m0 *1 178.365,152.88
X$32944 572 626 573 644 645 cell_1rw
* cell instance $32945 r0 *1 178.365,152.88
X$32945 572 627 573 644 645 cell_1rw
* cell instance $32946 m0 *1 178.365,155.61
X$32946 572 628 573 644 645 cell_1rw
* cell instance $32947 m0 *1 178.365,158.34
X$32947 572 630 573 644 645 cell_1rw
* cell instance $32948 r0 *1 178.365,155.61
X$32948 572 629 573 644 645 cell_1rw
* cell instance $32949 m0 *1 178.365,161.07
X$32949 572 632 573 644 645 cell_1rw
* cell instance $32950 r0 *1 178.365,158.34
X$32950 572 631 573 644 645 cell_1rw
* cell instance $32951 m0 *1 178.365,163.8
X$32951 572 634 573 644 645 cell_1rw
* cell instance $32952 r0 *1 178.365,161.07
X$32952 572 633 573 644 645 cell_1rw
* cell instance $32953 r0 *1 178.365,163.8
X$32953 572 635 573 644 645 cell_1rw
* cell instance $32954 m0 *1 178.365,166.53
X$32954 572 637 573 644 645 cell_1rw
* cell instance $32955 r0 *1 178.365,166.53
X$32955 572 636 573 644 645 cell_1rw
* cell instance $32956 m0 *1 178.365,169.26
X$32956 572 639 573 644 645 cell_1rw
* cell instance $32957 r0 *1 178.365,169.26
X$32957 572 638 573 644 645 cell_1rw
* cell instance $32958 m0 *1 178.365,171.99
X$32958 572 640 573 644 645 cell_1rw
* cell instance $32959 m0 *1 178.365,174.72
X$32959 572 642 573 644 645 cell_1rw
* cell instance $32960 r0 *1 178.365,171.99
X$32960 572 641 573 644 645 cell_1rw
* cell instance $32961 r0 *1 178.365,174.72
X$32961 572 643 573 644 645 cell_1rw
* cell instance $32962 m0 *1 179.07,90.09
X$32962 574 581 575 644 645 cell_1rw
* cell instance $32963 r0 *1 179.07,90.09
X$32963 574 580 575 644 645 cell_1rw
* cell instance $32964 m0 *1 179.07,92.82
X$32964 574 583 575 644 645 cell_1rw
* cell instance $32965 r0 *1 179.07,92.82
X$32965 574 582 575 644 645 cell_1rw
* cell instance $32966 m0 *1 179.07,95.55
X$32966 574 584 575 644 645 cell_1rw
* cell instance $32967 m0 *1 179.07,98.28
X$32967 574 586 575 644 645 cell_1rw
* cell instance $32968 r0 *1 179.07,95.55
X$32968 574 585 575 644 645 cell_1rw
* cell instance $32969 r0 *1 179.07,98.28
X$32969 574 587 575 644 645 cell_1rw
* cell instance $32970 m0 *1 179.07,101.01
X$32970 574 588 575 644 645 cell_1rw
* cell instance $32971 r0 *1 179.07,101.01
X$32971 574 589 575 644 645 cell_1rw
* cell instance $32972 m0 *1 179.07,103.74
X$32972 574 590 575 644 645 cell_1rw
* cell instance $32973 r0 *1 179.07,103.74
X$32973 574 591 575 644 645 cell_1rw
* cell instance $32974 m0 *1 179.07,106.47
X$32974 574 593 575 644 645 cell_1rw
* cell instance $32975 m0 *1 179.07,109.2
X$32975 574 594 575 644 645 cell_1rw
* cell instance $32976 r0 *1 179.07,106.47
X$32976 574 592 575 644 645 cell_1rw
* cell instance $32977 r0 *1 179.07,109.2
X$32977 574 595 575 644 645 cell_1rw
* cell instance $32978 m0 *1 179.07,111.93
X$32978 574 597 575 644 645 cell_1rw
* cell instance $32979 m0 *1 179.07,114.66
X$32979 574 598 575 644 645 cell_1rw
* cell instance $32980 r0 *1 179.07,111.93
X$32980 574 596 575 644 645 cell_1rw
* cell instance $32981 r0 *1 179.07,114.66
X$32981 574 599 575 644 645 cell_1rw
* cell instance $32982 m0 *1 179.07,117.39
X$32982 574 600 575 644 645 cell_1rw
* cell instance $32983 r0 *1 179.07,117.39
X$32983 574 601 575 644 645 cell_1rw
* cell instance $32984 m0 *1 179.07,120.12
X$32984 574 602 575 644 645 cell_1rw
* cell instance $32985 r0 *1 179.07,120.12
X$32985 574 603 575 644 645 cell_1rw
* cell instance $32986 m0 *1 179.07,122.85
X$32986 574 604 575 644 645 cell_1rw
* cell instance $32987 r0 *1 179.07,122.85
X$32987 574 605 575 644 645 cell_1rw
* cell instance $32988 m0 *1 179.07,125.58
X$32988 574 606 575 644 645 cell_1rw
* cell instance $32989 r0 *1 179.07,125.58
X$32989 574 607 575 644 645 cell_1rw
* cell instance $32990 m0 *1 179.07,128.31
X$32990 574 609 575 644 645 cell_1rw
* cell instance $32991 r0 *1 179.07,128.31
X$32991 574 608 575 644 645 cell_1rw
* cell instance $32992 m0 *1 179.07,131.04
X$32992 574 610 575 644 645 cell_1rw
* cell instance $32993 r0 *1 179.07,131.04
X$32993 574 611 575 644 645 cell_1rw
* cell instance $32994 m0 *1 179.07,133.77
X$32994 574 612 575 644 645 cell_1rw
* cell instance $32995 r0 *1 179.07,133.77
X$32995 574 613 575 644 645 cell_1rw
* cell instance $32996 m0 *1 179.07,136.5
X$32996 574 615 575 644 645 cell_1rw
* cell instance $32997 r0 *1 179.07,136.5
X$32997 574 614 575 644 645 cell_1rw
* cell instance $32998 m0 *1 179.07,139.23
X$32998 574 617 575 644 645 cell_1rw
* cell instance $32999 r0 *1 179.07,139.23
X$32999 574 616 575 644 645 cell_1rw
* cell instance $33000 m0 *1 179.07,141.96
X$33000 574 618 575 644 645 cell_1rw
* cell instance $33001 r0 *1 179.07,141.96
X$33001 574 619 575 644 645 cell_1rw
* cell instance $33002 m0 *1 179.07,144.69
X$33002 574 620 575 644 645 cell_1rw
* cell instance $33003 r0 *1 179.07,144.69
X$33003 574 621 575 644 645 cell_1rw
* cell instance $33004 m0 *1 179.07,147.42
X$33004 574 622 575 644 645 cell_1rw
* cell instance $33005 m0 *1 179.07,150.15
X$33005 574 624 575 644 645 cell_1rw
* cell instance $33006 r0 *1 179.07,147.42
X$33006 574 623 575 644 645 cell_1rw
* cell instance $33007 r0 *1 179.07,150.15
X$33007 574 625 575 644 645 cell_1rw
* cell instance $33008 m0 *1 179.07,152.88
X$33008 574 626 575 644 645 cell_1rw
* cell instance $33009 r0 *1 179.07,152.88
X$33009 574 627 575 644 645 cell_1rw
* cell instance $33010 m0 *1 179.07,155.61
X$33010 574 628 575 644 645 cell_1rw
* cell instance $33011 r0 *1 179.07,155.61
X$33011 574 629 575 644 645 cell_1rw
* cell instance $33012 m0 *1 179.07,158.34
X$33012 574 630 575 644 645 cell_1rw
* cell instance $33013 r0 *1 179.07,158.34
X$33013 574 631 575 644 645 cell_1rw
* cell instance $33014 m0 *1 179.07,161.07
X$33014 574 632 575 644 645 cell_1rw
* cell instance $33015 r0 *1 179.07,161.07
X$33015 574 633 575 644 645 cell_1rw
* cell instance $33016 m0 *1 179.07,163.8
X$33016 574 634 575 644 645 cell_1rw
* cell instance $33017 r0 *1 179.07,163.8
X$33017 574 635 575 644 645 cell_1rw
* cell instance $33018 m0 *1 179.07,166.53
X$33018 574 637 575 644 645 cell_1rw
* cell instance $33019 r0 *1 179.07,166.53
X$33019 574 636 575 644 645 cell_1rw
* cell instance $33020 m0 *1 179.07,169.26
X$33020 574 639 575 644 645 cell_1rw
* cell instance $33021 r0 *1 179.07,169.26
X$33021 574 638 575 644 645 cell_1rw
* cell instance $33022 m0 *1 179.07,171.99
X$33022 574 640 575 644 645 cell_1rw
* cell instance $33023 r0 *1 179.07,171.99
X$33023 574 641 575 644 645 cell_1rw
* cell instance $33024 m0 *1 179.07,174.72
X$33024 574 642 575 644 645 cell_1rw
* cell instance $33025 r0 *1 179.07,174.72
X$33025 574 643 575 644 645 cell_1rw
* cell instance $33026 m0 *1 179.775,90.09
X$33026 576 581 577 644 645 cell_1rw
* cell instance $33027 r0 *1 179.775,90.09
X$33027 576 580 577 644 645 cell_1rw
* cell instance $33028 m0 *1 179.775,92.82
X$33028 576 583 577 644 645 cell_1rw
* cell instance $33029 r0 *1 179.775,92.82
X$33029 576 582 577 644 645 cell_1rw
* cell instance $33030 m0 *1 179.775,95.55
X$33030 576 584 577 644 645 cell_1rw
* cell instance $33031 r0 *1 179.775,95.55
X$33031 576 585 577 644 645 cell_1rw
* cell instance $33032 m0 *1 179.775,98.28
X$33032 576 586 577 644 645 cell_1rw
* cell instance $33033 r0 *1 179.775,98.28
X$33033 576 587 577 644 645 cell_1rw
* cell instance $33034 m0 *1 179.775,101.01
X$33034 576 588 577 644 645 cell_1rw
* cell instance $33035 r0 *1 179.775,101.01
X$33035 576 589 577 644 645 cell_1rw
* cell instance $33036 m0 *1 179.775,103.74
X$33036 576 590 577 644 645 cell_1rw
* cell instance $33037 r0 *1 179.775,103.74
X$33037 576 591 577 644 645 cell_1rw
* cell instance $33038 m0 *1 179.775,106.47
X$33038 576 593 577 644 645 cell_1rw
* cell instance $33039 r0 *1 179.775,106.47
X$33039 576 592 577 644 645 cell_1rw
* cell instance $33040 m0 *1 179.775,109.2
X$33040 576 594 577 644 645 cell_1rw
* cell instance $33041 r0 *1 179.775,109.2
X$33041 576 595 577 644 645 cell_1rw
* cell instance $33042 m0 *1 179.775,111.93
X$33042 576 597 577 644 645 cell_1rw
* cell instance $33043 r0 *1 179.775,111.93
X$33043 576 596 577 644 645 cell_1rw
* cell instance $33044 m0 *1 179.775,114.66
X$33044 576 598 577 644 645 cell_1rw
* cell instance $33045 r0 *1 179.775,114.66
X$33045 576 599 577 644 645 cell_1rw
* cell instance $33046 m0 *1 179.775,117.39
X$33046 576 600 577 644 645 cell_1rw
* cell instance $33047 r0 *1 179.775,117.39
X$33047 576 601 577 644 645 cell_1rw
* cell instance $33048 m0 *1 179.775,120.12
X$33048 576 602 577 644 645 cell_1rw
* cell instance $33049 r0 *1 179.775,120.12
X$33049 576 603 577 644 645 cell_1rw
* cell instance $33050 m0 *1 179.775,122.85
X$33050 576 604 577 644 645 cell_1rw
* cell instance $33051 r0 *1 179.775,122.85
X$33051 576 605 577 644 645 cell_1rw
* cell instance $33052 m0 *1 179.775,125.58
X$33052 576 606 577 644 645 cell_1rw
* cell instance $33053 m0 *1 179.775,128.31
X$33053 576 609 577 644 645 cell_1rw
* cell instance $33054 r0 *1 179.775,125.58
X$33054 576 607 577 644 645 cell_1rw
* cell instance $33055 r0 *1 179.775,128.31
X$33055 576 608 577 644 645 cell_1rw
* cell instance $33056 m0 *1 179.775,131.04
X$33056 576 610 577 644 645 cell_1rw
* cell instance $33057 r0 *1 179.775,131.04
X$33057 576 611 577 644 645 cell_1rw
* cell instance $33058 m0 *1 179.775,133.77
X$33058 576 612 577 644 645 cell_1rw
* cell instance $33059 r0 *1 179.775,133.77
X$33059 576 613 577 644 645 cell_1rw
* cell instance $33060 m0 *1 179.775,136.5
X$33060 576 615 577 644 645 cell_1rw
* cell instance $33061 r0 *1 179.775,136.5
X$33061 576 614 577 644 645 cell_1rw
* cell instance $33062 m0 *1 179.775,139.23
X$33062 576 617 577 644 645 cell_1rw
* cell instance $33063 m0 *1 179.775,141.96
X$33063 576 618 577 644 645 cell_1rw
* cell instance $33064 r0 *1 179.775,139.23
X$33064 576 616 577 644 645 cell_1rw
* cell instance $33065 r0 *1 179.775,141.96
X$33065 576 619 577 644 645 cell_1rw
* cell instance $33066 m0 *1 179.775,144.69
X$33066 576 620 577 644 645 cell_1rw
* cell instance $33067 r0 *1 179.775,144.69
X$33067 576 621 577 644 645 cell_1rw
* cell instance $33068 m0 *1 179.775,147.42
X$33068 576 622 577 644 645 cell_1rw
* cell instance $33069 m0 *1 179.775,150.15
X$33069 576 624 577 644 645 cell_1rw
* cell instance $33070 r0 *1 179.775,147.42
X$33070 576 623 577 644 645 cell_1rw
* cell instance $33071 r0 *1 179.775,150.15
X$33071 576 625 577 644 645 cell_1rw
* cell instance $33072 m0 *1 179.775,152.88
X$33072 576 626 577 644 645 cell_1rw
* cell instance $33073 r0 *1 179.775,152.88
X$33073 576 627 577 644 645 cell_1rw
* cell instance $33074 m0 *1 179.775,155.61
X$33074 576 628 577 644 645 cell_1rw
* cell instance $33075 r0 *1 179.775,155.61
X$33075 576 629 577 644 645 cell_1rw
* cell instance $33076 m0 *1 179.775,158.34
X$33076 576 630 577 644 645 cell_1rw
* cell instance $33077 r0 *1 179.775,158.34
X$33077 576 631 577 644 645 cell_1rw
* cell instance $33078 m0 *1 179.775,161.07
X$33078 576 632 577 644 645 cell_1rw
* cell instance $33079 m0 *1 179.775,163.8
X$33079 576 634 577 644 645 cell_1rw
* cell instance $33080 r0 *1 179.775,161.07
X$33080 576 633 577 644 645 cell_1rw
* cell instance $33081 r0 *1 179.775,163.8
X$33081 576 635 577 644 645 cell_1rw
* cell instance $33082 m0 *1 179.775,166.53
X$33082 576 637 577 644 645 cell_1rw
* cell instance $33083 r0 *1 179.775,166.53
X$33083 576 636 577 644 645 cell_1rw
* cell instance $33084 m0 *1 179.775,169.26
X$33084 576 639 577 644 645 cell_1rw
* cell instance $33085 r0 *1 179.775,169.26
X$33085 576 638 577 644 645 cell_1rw
* cell instance $33086 m0 *1 179.775,171.99
X$33086 576 640 577 644 645 cell_1rw
* cell instance $33087 r0 *1 179.775,171.99
X$33087 576 641 577 644 645 cell_1rw
* cell instance $33088 m0 *1 179.775,174.72
X$33088 576 642 577 644 645 cell_1rw
* cell instance $33089 r0 *1 179.775,174.72
X$33089 576 643 577 644 645 cell_1rw
* cell instance $33090 m0 *1 180.48,90.09
X$33090 578 581 579 644 645 cell_1rw
* cell instance $33091 r0 *1 180.48,90.09
X$33091 578 580 579 644 645 cell_1rw
* cell instance $33092 m0 *1 180.48,92.82
X$33092 578 583 579 644 645 cell_1rw
* cell instance $33093 r0 *1 180.48,92.82
X$33093 578 582 579 644 645 cell_1rw
* cell instance $33094 m0 *1 180.48,95.55
X$33094 578 584 579 644 645 cell_1rw
* cell instance $33095 r0 *1 180.48,95.55
X$33095 578 585 579 644 645 cell_1rw
* cell instance $33096 m0 *1 180.48,98.28
X$33096 578 586 579 644 645 cell_1rw
* cell instance $33097 r0 *1 180.48,98.28
X$33097 578 587 579 644 645 cell_1rw
* cell instance $33098 m0 *1 180.48,101.01
X$33098 578 588 579 644 645 cell_1rw
* cell instance $33099 m0 *1 180.48,103.74
X$33099 578 590 579 644 645 cell_1rw
* cell instance $33100 r0 *1 180.48,101.01
X$33100 578 589 579 644 645 cell_1rw
* cell instance $33101 r0 *1 180.48,103.74
X$33101 578 591 579 644 645 cell_1rw
* cell instance $33102 m0 *1 180.48,106.47
X$33102 578 593 579 644 645 cell_1rw
* cell instance $33103 r0 *1 180.48,106.47
X$33103 578 592 579 644 645 cell_1rw
* cell instance $33104 m0 *1 180.48,109.2
X$33104 578 594 579 644 645 cell_1rw
* cell instance $33105 r0 *1 180.48,109.2
X$33105 578 595 579 644 645 cell_1rw
* cell instance $33106 m0 *1 180.48,111.93
X$33106 578 597 579 644 645 cell_1rw
* cell instance $33107 r0 *1 180.48,111.93
X$33107 578 596 579 644 645 cell_1rw
* cell instance $33108 m0 *1 180.48,114.66
X$33108 578 598 579 644 645 cell_1rw
* cell instance $33109 m0 *1 180.48,117.39
X$33109 578 600 579 644 645 cell_1rw
* cell instance $33110 r0 *1 180.48,114.66
X$33110 578 599 579 644 645 cell_1rw
* cell instance $33111 r0 *1 180.48,117.39
X$33111 578 601 579 644 645 cell_1rw
* cell instance $33112 m0 *1 180.48,120.12
X$33112 578 602 579 644 645 cell_1rw
* cell instance $33113 r0 *1 180.48,120.12
X$33113 578 603 579 644 645 cell_1rw
* cell instance $33114 m0 *1 180.48,122.85
X$33114 578 604 579 644 645 cell_1rw
* cell instance $33115 r0 *1 180.48,122.85
X$33115 578 605 579 644 645 cell_1rw
* cell instance $33116 m0 *1 180.48,125.58
X$33116 578 606 579 644 645 cell_1rw
* cell instance $33117 r0 *1 180.48,125.58
X$33117 578 607 579 644 645 cell_1rw
* cell instance $33118 m0 *1 180.48,128.31
X$33118 578 609 579 644 645 cell_1rw
* cell instance $33119 r0 *1 180.48,128.31
X$33119 578 608 579 644 645 cell_1rw
* cell instance $33120 m0 *1 180.48,131.04
X$33120 578 610 579 644 645 cell_1rw
* cell instance $33121 r0 *1 180.48,131.04
X$33121 578 611 579 644 645 cell_1rw
* cell instance $33122 m0 *1 180.48,133.77
X$33122 578 612 579 644 645 cell_1rw
* cell instance $33123 r0 *1 180.48,133.77
X$33123 578 613 579 644 645 cell_1rw
* cell instance $33124 m0 *1 180.48,136.5
X$33124 578 615 579 644 645 cell_1rw
* cell instance $33125 r0 *1 180.48,136.5
X$33125 578 614 579 644 645 cell_1rw
* cell instance $33126 m0 *1 180.48,139.23
X$33126 578 617 579 644 645 cell_1rw
* cell instance $33127 r0 *1 180.48,139.23
X$33127 578 616 579 644 645 cell_1rw
* cell instance $33128 m0 *1 180.48,141.96
X$33128 578 618 579 644 645 cell_1rw
* cell instance $33129 m0 *1 180.48,144.69
X$33129 578 620 579 644 645 cell_1rw
* cell instance $33130 r0 *1 180.48,141.96
X$33130 578 619 579 644 645 cell_1rw
* cell instance $33131 r0 *1 180.48,144.69
X$33131 578 621 579 644 645 cell_1rw
* cell instance $33132 m0 *1 180.48,147.42
X$33132 578 622 579 644 645 cell_1rw
* cell instance $33133 r0 *1 180.48,147.42
X$33133 578 623 579 644 645 cell_1rw
* cell instance $33134 m0 *1 180.48,150.15
X$33134 578 624 579 644 645 cell_1rw
* cell instance $33135 r0 *1 180.48,150.15
X$33135 578 625 579 644 645 cell_1rw
* cell instance $33136 m0 *1 180.48,152.88
X$33136 578 626 579 644 645 cell_1rw
* cell instance $33137 r0 *1 180.48,152.88
X$33137 578 627 579 644 645 cell_1rw
* cell instance $33138 m0 *1 180.48,155.61
X$33138 578 628 579 644 645 cell_1rw
* cell instance $33139 r0 *1 180.48,155.61
X$33139 578 629 579 644 645 cell_1rw
* cell instance $33140 m0 *1 180.48,158.34
X$33140 578 630 579 644 645 cell_1rw
* cell instance $33141 m0 *1 180.48,161.07
X$33141 578 632 579 644 645 cell_1rw
* cell instance $33142 r0 *1 180.48,158.34
X$33142 578 631 579 644 645 cell_1rw
* cell instance $33143 m0 *1 180.48,163.8
X$33143 578 634 579 644 645 cell_1rw
* cell instance $33144 r0 *1 180.48,161.07
X$33144 578 633 579 644 645 cell_1rw
* cell instance $33145 r0 *1 180.48,163.8
X$33145 578 635 579 644 645 cell_1rw
* cell instance $33146 m0 *1 180.48,166.53
X$33146 578 637 579 644 645 cell_1rw
* cell instance $33147 r0 *1 180.48,166.53
X$33147 578 636 579 644 645 cell_1rw
* cell instance $33148 m0 *1 180.48,169.26
X$33148 578 639 579 644 645 cell_1rw
* cell instance $33149 r0 *1 180.48,169.26
X$33149 578 638 579 644 645 cell_1rw
* cell instance $33150 m0 *1 180.48,171.99
X$33150 578 640 579 644 645 cell_1rw
* cell instance $33151 r0 *1 180.48,171.99
X$33151 578 641 579 644 645 cell_1rw
* cell instance $33152 m0 *1 180.48,174.72
X$33152 578 642 579 644 645 cell_1rw
* cell instance $33153 r0 *1 180.48,174.72
X$33153 578 643 579 644 645 cell_1rw
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_bitcell_array

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_0
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_0 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0
* pin A
* pin B
* pin C
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0 1 2 3 4 5 6
* net 1 A
* net 2 B
* net 3 C
* net 4 Z
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.2325,2.21 PMOS_VTG
M$1 5 1 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,2.21 PMOS_VTG
M$2 4 2 5 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.022275P PS=0.435U
+ PD=0.435U
* device instance $3 r0 *1 0.6625,2.21 PMOS_VTG
M$3 5 3 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $4 r0 *1 0.2325,0.215 NMOS_VTG
M$4 6 1 8 6 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $5 r0 *1 0.4475,0.215 NMOS_VTG
M$5 8 2 7 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.01485P PS=0.345U PD=0.345U
* device instance $6 r0 *1 0.6625,0.215 NMOS_VTG
M$6 7 3 4 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_0
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_0 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.186 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=5.7575U AS=0.64955625P AD=0.64955625P PS=16.485U
+ PD=16.485U
* device instance $48 r0 *1 0.2325,1.056 PMOS_VTG
M$48 3 1 2 3 PMOS_VTG L=0.05U W=17.2725U AS=1.94866875P AD=1.94866875P
+ PS=28.245U PD=28.245U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_0

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec
* pin Z
* pin A
* pin B
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec 2 3 4 5 6
* net 2 Z
* net 3 A
* net 4 B
* net 5 vdd
* net 6 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 1 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2
* cell instance $2 r0 *1 0.9025,0
X$2 1 2 5 6 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_and2_dec

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec
* pin Z
* pin A
* pin B
* pin C
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec 2 3 4 5 6 7
* net 2 Z
* net 3 A
* net 4 B
* net 5 C
* net 6 vdd
* net 7 gnd
* cell instance $1 r0 *1 0,0
X$1 3 4 5 1 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3
* cell instance $2 r0 *1 1.2475,0
X$2 1 2 6 7 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_and3_dec

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver
* pin Z
* pin A
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver 1 2 3 4
* net 1 Z
* net 2 A
* net 3 vdd
* net 4 gnd
* cell instance $1 r0 *1 0,0
X$1 2 1 3 4 freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_1
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pdriver

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_0
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_0 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,1.56 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.56 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2_0

* cell dummy_cell_1rw
* pin wl
* pin vdd
* pin gnd
.SUBCKT dummy_cell_1rw 2 6 7
* net 2 wl
* net 6 vdd
* net 7 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 1 6 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.00945P PS=0.39U PD=0.39U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 6 5 1 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.00945P PS=0.39U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 1 7 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.021525P PS=0.62U
+ PD=0.62U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 7 5 1 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.021525P PS=0.62U
+ PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 3 2 5 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 1 2 4 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS dummy_cell_1rw

* cell replica_cell_1rw
* pin bl
* pin wl
* pin br
* pin vdd
* pin gnd
.SUBCKT replica_cell_1rw 1 2 4 5 6
* net 1 bl
* net 2 wl
* net 4 br
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 3 5 5 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0099P PS=0.39U PD=0.4U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 5 5 3 5 PMOS_VTG L=0.05U W=0.09U AS=0.0099P AD=0.00945P PS=0.4U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 3 6 6 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.02255P PS=0.62U PD=0.63U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 6 5 3 6 NMOS_VTG L=0.05U W=0.205U AS=0.02255P AD=0.021525P PS=0.63U PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 4 2 5 6 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 3 2 1 6 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS replica_cell_1rw

* cell cell_1rw
* pin bl
* pin wl
* pin br
* pin vdd
* pin gnd
.SUBCKT cell_1rw 1 2 4 6 7
* net 1 bl
* net 2 wl
* net 3 Q
* net 4 br
* net 5 Q_bar
* net 6 vdd
* net 7 gnd
* device instance $1 r0 *1 0.61,1.2075 PMOS_VTG
M$1 5 3 6 6 PMOS_VTG L=0.05U W=0.09U AS=0.00945P AD=0.0099P PS=0.39U PD=0.4U
* device instance $2 r0 *1 0.095,1.2075 PMOS_VTG
M$2 6 5 3 6 PMOS_VTG L=0.05U W=0.09U AS=0.0099P AD=0.00945P PS=0.4U PD=0.39U
* device instance $3 r0 *1 0.61,0.67 NMOS_VTG
M$3 5 3 7 7 NMOS_VTG L=0.05U W=0.205U AS=0.021525P AD=0.02255P PS=0.62U PD=0.63U
* device instance $4 r0 *1 0.095,0.67 NMOS_VTG
M$4 7 5 3 7 NMOS_VTG L=0.05U W=0.205U AS=0.02255P AD=0.021525P PS=0.63U PD=0.62U
* device instance $5 r0 *1 0.53,0.315 NMOS_VTG
M$5 4 2 5 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
* device instance $6 r0 *1 0.175,0.315 NMOS_VTG
M$6 3 2 1 7 NMOS_VTG L=0.05U W=0.135U AS=0.014175P AD=0.014175P PS=0.48U
+ PD=0.48U
.ENDS cell_1rw

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,2.21 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_2

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2
* pin A
* pin B
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2 1 2 3 4 5
* net 1 A
* net 2 B
* net 3 Z
* net 4 vdd
* net 5 gnd
* device instance $1 r0 *1 0.2325,1.105 PMOS_VTG
M$1 4 1 3 4 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.105 PMOS_VTG
M$2 3 2 4 4 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $3 r0 *1 0.2325,0.215 NMOS_VTG
M$3 5 1 6 5 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $4 r0 *1 0.4475,0.215 NMOS_VTG
M$4 6 2 3 5 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand2

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.17 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.09U AS=0.011475P AD=0.011475P PS=0.435U
+ PD=0.435U
* device instance $2 r0 *1 0.2325,1.105 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.034425P PS=0.795U
+ PD=0.795U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3
* pin A
* pin B
* pin C
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3 1 2 3 4 5 6
* net 1 A
* net 2 B
* net 3 C
* net 4 Z
* net 5 vdd
* net 6 gnd
* device instance $1 r0 *1 0.2325,1.105 PMOS_VTG
M$1 5 1 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.034425P AD=0.022275P PS=0.795U
+ PD=0.435U
* device instance $2 r0 *1 0.4475,1.105 PMOS_VTG
M$2 4 2 5 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.022275P PS=0.435U
+ PD=0.435U
* device instance $3 r0 *1 0.6625,1.105 PMOS_VTG
M$3 5 3 4 5 PMOS_VTG L=0.05U W=0.27U AS=0.022275P AD=0.034425P PS=0.435U
+ PD=0.795U
* device instance $4 r0 *1 0.2325,0.215 NMOS_VTG
M$4 6 1 8 6 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.01485P PS=0.615U PD=0.345U
* device instance $5 r0 *1 0.4475,0.215 NMOS_VTG
M$5 8 2 7 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.01485P PS=0.345U PD=0.345U
* device instance $6 r0 *1 0.6625,0.215 NMOS_VTG
M$6 7 3 4 6 NMOS_VTG L=0.05U W=0.18U AS=0.01485P AD=0.02295P PS=0.345U PD=0.615U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pnand3

* cell freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_1
* pin A
* pin Z
* pin vdd
* pin gnd
.SUBCKT freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_1 1 2 3 4
* net 1 A
* net 2 Z
* net 3 vdd
* net 4 gnd
* device instance $1 r0 *1 0.2325,0.215 NMOS_VTG
M$1 4 1 2 4 NMOS_VTG L=0.05U W=0.18U AS=0.02295P AD=0.02295P PS=0.615U PD=0.615U
* device instance $2 r0 *1 0.2325,1.425 PMOS_VTG
M$2 3 1 2 3 PMOS_VTG L=0.05U W=0.54U AS=0.06885P AD=0.06885P PS=1.335U PD=1.335U
.ENDS freepdk45_sram_4kbytes_1rw_32x1024_8_pinv_1
