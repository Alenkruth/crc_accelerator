VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO freepdk45_sram_4kbytes_1rw_32x1024_8
   CLASS BLOCK ;
   SIZE 239.82 BY 218.26 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.6 0.0 47.74 0.42 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.4 0.0 50.54 0.42 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.48 0.0 53.62 0.42 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.28 0.0 56.42 0.42 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.8 0.0 58.94 0.42 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.88 0.0 62.02 0.42 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.96 0.0 65.1 0.42 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.48 0.0 67.62 0.42 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.56 0.0 70.7 0.42 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.08 0.0 73.22 0.42 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.16 0.0 76.3 0.42 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.96 0.0 79.1 0.42 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.04 0.0 82.18 0.42 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.84 0.0 84.98 0.42 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.64 0.0 87.78 0.42 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.44 0.0 90.58 0.42 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.52 0.0 93.66 0.42 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.32 0.0 96.46 0.42 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.12 0.0 99.26 0.42 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.92 0.0 102.06 0.42 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.72 0.0 104.86 0.42 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.8 0.0 107.94 0.42 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.32 0.0 110.46 0.42 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.4 0.0 113.54 0.42 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.2 0.0 116.34 0.42 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.28 0.0 119.42 0.42 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  122.08 0.0 122.22 0.42 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  124.6 0.0 124.74 0.42 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  127.68 0.0 127.82 0.42 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  130.48 0.0 130.62 0.42 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  133.28 0.0 133.42 0.42 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  136.08 0.0 136.22 0.42 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  139.16 0.0 139.3 0.42 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  27.72 0.0 27.86 0.42 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  30.52 0.0 30.66 0.42 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  33.04 0.0 33.18 0.42 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 71.4 0.42 71.54 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 73.92 0.42 74.06 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 76.16 0.42 76.3 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 79.24 0.42 79.38 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 80.92 0.42 81.06 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 83.72 0.42 83.86 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 86.24 0.42 86.38 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 88.76 0.42 88.9 ;
      END
   END addr0[10]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 15.68 0.42 15.82 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 18.2 0.42 18.34 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 15.96 0.42 16.1 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  36.12 0.0 36.26 0.42 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.92 0.0 39.06 0.42 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.72 0.0 41.86 0.42 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.8 0.0 44.94 0.42 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  141.96 0.0 142.1 0.42 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  54.32 0.0 54.46 0.42 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  59.08 0.0 59.22 0.42 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.68 0.0 64.82 0.42 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.28 0.0 70.42 0.42 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.72 0.0 76.86 0.42 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  82.32 0.0 82.46 0.42 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  86.8 0.0 86.94 0.42 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.8 0.0 93.94 0.42 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  98.0 0.0 98.14 0.42 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  103.88 0.0 104.02 0.42 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  109.48 0.0 109.62 0.42 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  115.36 0.0 115.5 0.42 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  120.96 0.0 121.1 0.42 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  126.56 0.0 126.7 0.42 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  132.44 0.0 132.58 0.42 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  138.04 0.0 138.18 0.42 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  143.36 0.0 143.5 0.42 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  149.24 0.0 149.38 0.42 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  154.84 0.0 154.98 0.42 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  160.44 0.0 160.58 0.42 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  166.04 0.0 166.18 0.42 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  171.92 0.0 172.06 0.42 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  177.52 0.0 177.66 0.42 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  183.12 0.0 183.26 0.42 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  188.44 0.0 188.58 0.42 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  194.32 0.0 194.46 0.42 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  199.92 0.0 200.06 0.42 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  205.52 0.0 205.66 0.42 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  211.4 0.0 211.54 0.42 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.4 22.96 239.82 23.1 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.4 24.08 239.82 24.22 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.4 23.24 239.82 23.38 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  239.4 23.52 239.82 23.66 ;
      END
   END dout0[32]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  1.4 216.16 238.42 216.86 ;
         LAYER metal4 ;
         RECT  237.72 1.4 238.42 216.86 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 216.86 ;
         LAYER metal3 ;
         RECT  1.4 1.4 238.42 2.1 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 0.0 239.82 0.7 ;
         LAYER metal4 ;
         RECT  239.12 0.0 239.82 218.26 ;
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 218.26 ;
         LAYER metal3 ;
         RECT  0.0 217.56 239.82 218.26 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 239.68 218.12 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 239.68 218.12 ;
   LAYER  metal3 ;
      RECT  0.56 71.26 239.68 71.68 ;
      RECT  0.14 71.68 0.56 73.78 ;
      RECT  0.14 74.2 0.56 76.02 ;
      RECT  0.14 76.44 0.56 79.1 ;
      RECT  0.14 79.52 0.56 80.78 ;
      RECT  0.14 81.2 0.56 83.58 ;
      RECT  0.14 84.0 0.56 86.1 ;
      RECT  0.14 86.52 0.56 88.62 ;
      RECT  0.14 18.48 0.56 71.26 ;
      RECT  0.14 16.24 0.56 18.06 ;
      RECT  0.56 22.82 239.26 23.24 ;
      RECT  0.56 23.24 239.26 71.26 ;
      RECT  239.26 24.36 239.68 71.26 ;
      RECT  239.26 23.8 239.68 23.94 ;
      RECT  0.56 71.68 1.26 216.02 ;
      RECT  0.56 216.02 1.26 217.0 ;
      RECT  1.26 71.68 238.56 216.02 ;
      RECT  238.56 71.68 239.68 216.02 ;
      RECT  238.56 216.02 239.68 217.0 ;
      RECT  0.56 1.26 1.26 2.24 ;
      RECT  0.56 2.24 1.26 22.82 ;
      RECT  1.26 2.24 238.56 22.82 ;
      RECT  238.56 1.26 239.26 2.24 ;
      RECT  238.56 2.24 239.26 22.82 ;
      RECT  0.14 0.84 0.56 15.54 ;
      RECT  239.26 0.84 239.68 22.82 ;
      RECT  0.56 0.84 1.26 1.26 ;
      RECT  1.26 0.84 238.56 1.26 ;
      RECT  238.56 0.84 239.26 1.26 ;
      RECT  0.14 89.04 0.56 217.42 ;
      RECT  0.56 217.0 1.26 217.42 ;
      RECT  1.26 217.0 238.56 217.42 ;
      RECT  238.56 217.0 239.68 217.42 ;
   LAYER  metal4 ;
      RECT  47.32 0.7 48.02 218.12 ;
      RECT  48.02 0.14 50.12 0.7 ;
      RECT  50.82 0.14 53.2 0.7 ;
      RECT  56.7 0.14 58.52 0.7 ;
      RECT  65.38 0.14 67.2 0.7 ;
      RECT  70.98 0.14 72.8 0.7 ;
      RECT  73.5 0.14 75.88 0.7 ;
      RECT  79.38 0.14 81.76 0.7 ;
      RECT  88.06 0.14 90.16 0.7 ;
      RECT  90.86 0.14 93.24 0.7 ;
      RECT  99.54 0.14 101.64 0.7 ;
      RECT  105.14 0.14 107.52 0.7 ;
      RECT  110.74 0.14 113.12 0.7 ;
      RECT  116.62 0.14 119.0 0.7 ;
      RECT  122.5 0.14 124.32 0.7 ;
      RECT  128.1 0.14 130.2 0.7 ;
      RECT  133.7 0.14 135.8 0.7 ;
      RECT  28.14 0.14 30.24 0.7 ;
      RECT  30.94 0.14 32.76 0.7 ;
      RECT  33.46 0.14 35.84 0.7 ;
      RECT  36.54 0.14 38.64 0.7 ;
      RECT  39.34 0.14 41.44 0.7 ;
      RECT  42.14 0.14 44.52 0.7 ;
      RECT  45.22 0.14 47.32 0.7 ;
      RECT  139.58 0.14 141.68 0.7 ;
      RECT  53.9 0.14 54.04 0.7 ;
      RECT  54.74 0.14 56.0 0.7 ;
      RECT  59.5 0.14 61.6 0.7 ;
      RECT  62.3 0.14 64.4 0.7 ;
      RECT  67.9 0.14 70.0 0.7 ;
      RECT  77.14 0.14 78.68 0.7 ;
      RECT  82.74 0.14 84.56 0.7 ;
      RECT  85.26 0.14 86.52 0.7 ;
      RECT  87.22 0.14 87.36 0.7 ;
      RECT  94.22 0.14 96.04 0.7 ;
      RECT  96.74 0.14 97.72 0.7 ;
      RECT  98.42 0.14 98.84 0.7 ;
      RECT  102.34 0.14 103.6 0.7 ;
      RECT  104.3 0.14 104.44 0.7 ;
      RECT  108.22 0.14 109.2 0.7 ;
      RECT  109.9 0.14 110.04 0.7 ;
      RECT  113.82 0.14 115.08 0.7 ;
      RECT  115.78 0.14 115.92 0.7 ;
      RECT  119.7 0.14 120.68 0.7 ;
      RECT  121.38 0.14 121.8 0.7 ;
      RECT  125.02 0.14 126.28 0.7 ;
      RECT  126.98 0.14 127.4 0.7 ;
      RECT  130.9 0.14 132.16 0.7 ;
      RECT  132.86 0.14 133.0 0.7 ;
      RECT  136.5 0.14 137.76 0.7 ;
      RECT  138.46 0.14 138.88 0.7 ;
      RECT  142.38 0.14 143.08 0.7 ;
      RECT  143.78 0.14 148.96 0.7 ;
      RECT  149.66 0.14 154.56 0.7 ;
      RECT  155.26 0.14 160.16 0.7 ;
      RECT  160.86 0.14 165.76 0.7 ;
      RECT  166.46 0.14 171.64 0.7 ;
      RECT  172.34 0.14 177.24 0.7 ;
      RECT  177.94 0.14 182.84 0.7 ;
      RECT  183.54 0.14 188.16 0.7 ;
      RECT  188.86 0.14 194.04 0.7 ;
      RECT  194.74 0.14 199.64 0.7 ;
      RECT  200.34 0.14 205.24 0.7 ;
      RECT  205.94 0.14 211.12 0.7 ;
      RECT  48.02 0.7 237.44 1.12 ;
      RECT  48.02 1.12 237.44 217.14 ;
      RECT  48.02 217.14 237.44 218.12 ;
      RECT  237.44 0.7 238.7 1.12 ;
      RECT  237.44 217.14 238.7 218.12 ;
      RECT  1.12 0.7 2.38 1.12 ;
      RECT  1.12 217.14 2.38 218.12 ;
      RECT  2.38 0.7 47.32 1.12 ;
      RECT  2.38 1.12 47.32 217.14 ;
      RECT  2.38 217.14 47.32 218.12 ;
      RECT  211.82 0.14 238.84 0.7 ;
      RECT  238.7 0.7 238.84 1.12 ;
      RECT  238.7 1.12 238.84 217.14 ;
      RECT  238.7 217.14 238.84 218.12 ;
      RECT  0.98 0.14 27.44 0.7 ;
      RECT  0.98 0.7 1.12 1.12 ;
      RECT  0.98 1.12 1.12 217.14 ;
      RECT  0.98 217.14 1.12 218.12 ;
   END
END    freepdk45_sram_4kbytes_1rw_32x1024_8
END    LIBRARY
